module fake_jpeg_13425_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_51),
.B(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_54),
.B(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_56),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_13),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_12),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_88),
.Y(n_118)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_12),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_64),
.B(n_73),
.Y(n_113)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_12),
.B(n_11),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_69),
.B(n_76),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_23),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_17),
.B(n_0),
.CON(n_74),
.SN(n_74)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_86),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_11),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_11),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_23),
.B(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_92),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_17),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_32),
.B(n_10),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_98),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_33),
.B(n_10),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_48),
.B1(n_46),
.B2(n_36),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_116),
.B1(n_120),
.B2(n_140),
.Y(n_159)
);

CKINVDCx12_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_105),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_48),
.B1(n_46),
.B2(n_36),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_49),
.A2(n_48),
.B1(n_46),
.B2(n_36),
.Y(n_120)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_74),
.A2(n_48),
.B1(n_40),
.B2(n_39),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_63),
.B(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_66),
.B(n_37),
.Y(n_145)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_149),
.Y(n_193)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_84),
.B(n_37),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_30),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_90),
.A2(n_35),
.B1(n_31),
.B2(n_34),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_93),
.B1(n_91),
.B2(n_82),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_94),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_156),
.A2(n_97),
.B1(n_96),
.B2(n_95),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_160),
.A2(n_202),
.B1(n_75),
.B2(n_70),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_88),
.B1(n_30),
.B2(n_28),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_71),
.C(n_87),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_205),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_100),
.B(n_51),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_53),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_177),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_40),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_37),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_127),
.B(n_39),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_179),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_113),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_21),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_185),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_129),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_186),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_114),
.B(n_21),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_112),
.B(n_39),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_106),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_25),
.B1(n_27),
.B2(n_24),
.Y(n_208)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_195),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_103),
.B(n_39),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_40),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_201),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_198),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_147),
.B(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_207),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_204),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_101),
.A2(n_56),
.B(n_30),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_144),
.B(n_27),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_27),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_208),
.A2(n_21),
.B(n_24),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_158),
.A2(n_120),
.B1(n_116),
.B2(n_144),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_220),
.B1(n_221),
.B2(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_159),
.A2(n_141),
.B1(n_102),
.B2(n_155),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_225),
.B(n_173),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_165),
.A2(n_155),
.B1(n_157),
.B2(n_150),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_167),
.A2(n_157),
.B1(n_150),
.B2(n_111),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_148),
.B1(n_139),
.B2(n_108),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_185),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_203),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_160),
.A2(n_111),
.B1(n_133),
.B2(n_136),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_194),
.B1(n_108),
.B2(n_168),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_238),
.B(n_25),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_180),
.B(n_148),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_242),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_146),
.B1(n_109),
.B2(n_136),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_243),
.B1(n_207),
.B2(n_188),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_139),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_162),
.A2(n_146),
.B1(n_109),
.B2(n_133),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_25),
.B(n_24),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_179),
.B(n_181),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_171),
.C(n_190),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_209),
.B(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_247),
.B(n_251),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_176),
.B1(n_184),
.B2(n_193),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_249),
.A2(n_250),
.B(n_260),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_191),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_256),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_261),
.B1(n_240),
.B2(n_210),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_209),
.B(n_187),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_264),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_182),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_259),
.Y(n_294)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_182),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_238),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_217),
.B1(n_211),
.B2(n_218),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_263),
.B1(n_217),
.B2(n_234),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_50),
.B1(n_81),
.B2(n_79),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_266),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_200),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_268),
.Y(n_295)
);

BUFx12_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_269),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_279),
.B(n_208),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_272),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_200),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_199),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_161),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_215),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_128),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_246),
.Y(n_301)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_224),
.A2(n_193),
.B1(n_161),
.B2(n_173),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_280),
.A2(n_291),
.B1(n_298),
.B2(n_307),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_285),
.A2(n_296),
.B1(n_299),
.B2(n_312),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_253),
.Y(n_286)
);

INVx13_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_287),
.A2(n_250),
.B(n_249),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_289),
.B(n_271),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_211),
.B1(n_230),
.B2(n_225),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_230),
.A3(n_222),
.B1(n_213),
.B2(n_244),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_300),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_248),
.A2(n_228),
.B1(n_208),
.B2(n_225),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_261),
.A2(n_243),
.B1(n_221),
.B2(n_225),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_248),
.A2(n_260),
.B1(n_252),
.B2(n_250),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_266),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_302),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_245),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_301),
.C(n_297),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_256),
.Y(n_303)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_225),
.B1(n_215),
.B2(n_237),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_248),
.A2(n_244),
.B1(n_227),
.B2(n_223),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_265),
.A2(n_237),
.B1(n_241),
.B2(n_233),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_313),
.A2(n_260),
.B1(n_263),
.B2(n_262),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_269),
.Y(n_314)
);

INVx13_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_259),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_315),
.B(n_326),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_321),
.C(n_329),
.Y(n_351)
);

OAI221xp5_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_257),
.B1(n_273),
.B2(n_251),
.C(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_320),
.B(n_330),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_322),
.A2(n_287),
.B(n_307),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_304),
.Y(n_323)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_323),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_296),
.A2(n_249),
.B(n_263),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_324),
.A2(n_334),
.B(n_281),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_260),
.C(n_277),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_294),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_294),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_338),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_333),
.A2(n_283),
.B1(n_282),
.B2(n_237),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_279),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_311),
.A2(n_270),
.B(n_279),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_335),
.A2(n_166),
.B(n_189),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_262),
.B1(n_277),
.B2(n_258),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_336),
.A2(n_346),
.B1(n_60),
.B2(n_67),
.Y(n_379)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_305),
.B(n_226),
.C(n_229),
.Y(n_338)
);

INVx3_ASAP7_75t_SL g339 ( 
.A(n_312),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_305),
.B(n_293),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_343),
.C(n_345),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_229),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_344),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_241),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_284),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_311),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_285),
.A2(n_258),
.B1(n_237),
.B2(n_223),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_288),
.B(n_216),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_343),
.C(n_328),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_306),
.Y(n_348)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_349),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_308),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_356),
.Y(n_387)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_354),
.A2(n_360),
.B(n_375),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_SL g355 ( 
.A(n_335),
.B(n_345),
.Y(n_355)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_280),
.Y(n_356)
);

AOI22x1_ASAP7_75t_L g357 ( 
.A1(n_316),
.A2(n_298),
.B1(n_304),
.B2(n_309),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_364),
.B1(n_370),
.B2(n_382),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_340),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_380),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_332),
.A2(n_281),
.B1(n_283),
.B2(n_314),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_366),
.A2(n_367),
.B1(n_372),
.B2(n_327),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_282),
.B1(n_290),
.B2(n_216),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_290),
.Y(n_369)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_199),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_324),
.A2(n_226),
.B1(n_268),
.B2(n_278),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_317),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_175),
.Y(n_374)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_193),
.C(n_187),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_322),
.C(n_346),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_323),
.B(n_175),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_197),
.B1(n_169),
.B2(n_31),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_269),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_339),
.A2(n_47),
.B1(n_43),
.B2(n_45),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_317),
.B(n_278),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_198),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_385),
.B(n_390),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_333),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_386),
.B(n_400),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_391),
.A2(n_395),
.B1(n_357),
.B2(n_198),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_352),
.B(n_334),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_399),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_350),
.A2(n_365),
.B1(n_368),
.B2(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_325),
.B1(n_324),
.B2(n_327),
.Y(n_394)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_371),
.A2(n_325),
.B1(n_338),
.B2(n_337),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_396),
.Y(n_428)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_349),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_169),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_377),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_401),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_367),
.A2(n_268),
.B1(n_34),
.B2(n_35),
.Y(n_402)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_269),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_406),
.Y(n_431)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_404),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_358),
.Y(n_405)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_269),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_383),
.A2(n_164),
.B1(n_35),
.B2(n_34),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_409),
.A2(n_377),
.B1(n_381),
.B2(n_370),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_164),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_411),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_357),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_353),
.B(n_0),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_413),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_363),
.C(n_359),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_414),
.B(n_420),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_396),
.Y(n_418)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_405),
.Y(n_419)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_380),
.C(n_364),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_422),
.A2(n_391),
.B1(n_408),
.B2(n_407),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_376),
.C(n_366),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_438),
.C(n_412),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_360),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_427),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_354),
.B(n_375),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_426),
.A2(n_390),
.B(n_389),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_372),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_433),
.A2(n_40),
.B(n_22),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_68),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_198),
.C(n_35),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_421),
.A2(n_398),
.B(n_384),
.Y(n_439)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_440),
.A2(n_457),
.B(n_22),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_446),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_385),
.C(n_410),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_445),
.C(n_452),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_417),
.A2(n_397),
.B(n_410),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_443),
.A2(n_427),
.B(n_435),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_399),
.C(n_392),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_395),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_447),
.A2(n_458),
.B1(n_416),
.B2(n_434),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_404),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_449),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_409),
.Y(n_451)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_34),
.C(n_102),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_102),
.C(n_68),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_456),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_420),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_22),
.C(n_20),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_447),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_473),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_464),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_448),
.A2(n_424),
.B(n_433),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_463),
.A2(n_477),
.B(n_458),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_432),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_432),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_476),
.Y(n_478)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_428),
.B1(n_436),
.B2(n_416),
.Y(n_468)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_445),
.A2(n_426),
.B1(n_422),
.B2(n_438),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_437),
.B1(n_40),
.B2(n_4),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_469),
.A2(n_453),
.B(n_444),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_485),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_472),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_482),
.B(n_484),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_444),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_468),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_442),
.C(n_455),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_486),
.B(n_489),
.Y(n_498)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_487),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_473),
.A2(n_463),
.B(n_475),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_456),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_22),
.C(n_5),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_452),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_491),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_493),
.A2(n_454),
.B1(n_477),
.B2(n_465),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_497),
.Y(n_512)
);

NOR3xp33_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_474),
.C(n_464),
.Y(n_497)
);

AOI321xp33_ASAP7_75t_L g499 ( 
.A1(n_480),
.A2(n_462),
.A3(n_22),
.B1(n_4),
.B2(n_5),
.C(n_0),
.Y(n_499)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_499),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_486),
.A2(n_0),
.B(n_3),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_500),
.A2(n_502),
.B(n_485),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_479),
.A2(n_0),
.B(n_3),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_504),
.B(n_505),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_481),
.C(n_483),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_508),
.Y(n_515)
);

AOI322xp5_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_498),
.A3(n_494),
.B1(n_501),
.B2(n_492),
.C1(n_496),
.C2(n_505),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_511),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_481),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_501),
.B(n_491),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_478),
.C(n_5),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g514 ( 
.A(n_512),
.B(n_478),
.C(n_487),
.Y(n_514)
);

NOR3xp33_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_516),
.C(n_517),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_510),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_518),
.B(n_506),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_521),
.B(n_6),
.Y(n_522)
);

AOI322xp5_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_482),
.C2(n_503),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_522),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_519),
.B(n_6),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_6),
.Y(n_525)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_525),
.Y(n_526)
);


endmodule