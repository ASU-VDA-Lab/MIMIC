module fake_ibex_1096_n_863 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_863);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_863;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_841;
wire n_679;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_801;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_179;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_285;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_231;
wire n_298;
wire n_159;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_18),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_0),
.Y(n_154)
);

BUFx8_ASAP7_75t_SL g155 ( 
.A(n_86),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_26),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_38),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_90),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_31),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_78),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_54),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_21),
.B(n_70),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_55),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_53),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_82),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_10),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_30),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_36),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_121),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_58),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_18),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_21),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_84),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_29),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_67),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_19),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_87),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_107),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_56),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_88),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_43),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_63),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_1),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_51),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_2),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_66),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_4),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_131),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_136),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_100),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_L g213 ( 
.A(n_117),
.B(n_77),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_42),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_26),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_75),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_72),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_44),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g224 ( 
.A(n_125),
.B(n_22),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_105),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_146),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_143),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_19),
.Y(n_228)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_139),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_5),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_76),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_49),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_31),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_32),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_115),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_17),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_35),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_92),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_17),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_79),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_47),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_81),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_122),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_102),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_60),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_101),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_89),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_46),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_95),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_57),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_133),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_94),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_23),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_190),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_176),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_176),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_152),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_3),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g271 ( 
.A1(n_215),
.A2(n_74),
.B(n_149),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_160),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_73),
.B(n_148),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_181),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_157),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_158),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_194),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_157),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_155),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_174),
.B(n_6),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_199),
.Y(n_284)
);

BUFx8_ASAP7_75t_SL g285 ( 
.A(n_190),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_155),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_175),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_210),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_162),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_197),
.B(n_8),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_197),
.B(n_9),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_200),
.B(n_9),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_165),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_153),
.B(n_10),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_154),
.B(n_163),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_166),
.A2(n_80),
.B(n_147),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_230),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_203),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_156),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_203),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_177),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_168),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_14),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_170),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_172),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_173),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g309 ( 
.A(n_167),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_175),
.A2(n_15),
.B1(n_16),
.B2(n_20),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_210),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_180),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_203),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_193),
.B(n_20),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_183),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_257),
.B(n_24),
.Y(n_316)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_182),
.Y(n_319)
);

CKINVDCx8_ASAP7_75t_R g320 ( 
.A(n_229),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_210),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_184),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_186),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_223),
.B(n_25),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_243),
.B(n_25),
.Y(n_325)
);

OAI22x1_ASAP7_75t_SL g326 ( 
.A1(n_183),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_202),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_187),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_216),
.Y(n_330)
);

CKINVDCx6p67_ASAP7_75t_R g331 ( 
.A(n_164),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_228),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_236),
.B(n_28),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_275),
.A2(n_260),
.B1(n_232),
.B2(n_235),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_280),
.B(n_164),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_280),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_286),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_329),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_261),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_269),
.B(n_191),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_269),
.B(n_195),
.Y(n_347)
);

NAND2xp33_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_161),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_223),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_290),
.A2(n_260),
.B1(n_232),
.B2(n_241),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_277),
.B(n_289),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_286),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_241),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_331),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_277),
.B(n_205),
.Y(n_358)
);

AND3x2_ASAP7_75t_L g359 ( 
.A(n_287),
.B(n_250),
.C(n_244),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_290),
.A2(n_178),
.B1(n_185),
.B2(n_208),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_261),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_161),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_267),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_273),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_279),
.B(n_224),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_289),
.B(n_212),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_304),
.B(n_214),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_278),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_329),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_291),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_291),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_278),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_329),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_316),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_278),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_279),
.B(n_169),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_278),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_284),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_273),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_282),
.B(n_169),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_284),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_327),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_282),
.B(n_171),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_284),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_288),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_300),
.B(n_171),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_276),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_293),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_276),
.A2(n_196),
.B1(n_198),
.B2(n_246),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_300),
.B(n_318),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_308),
.B(n_219),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_308),
.B(n_221),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_300),
.B(n_222),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_SL g399 ( 
.A(n_324),
.B(n_196),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_272),
.B(n_207),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_296),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_318),
.B(n_207),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_318),
.B(n_231),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_324),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_299),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_296),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_296),
.Y(n_409)
);

BUFx6f_ASAP7_75t_SL g410 ( 
.A(n_312),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_299),
.Y(n_411)
);

OR2x6_ASAP7_75t_L g412 ( 
.A(n_265),
.B(n_198),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_406),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_270),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_387),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_372),
.A2(n_309),
.B1(n_292),
.B2(n_281),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_317),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_317),
.Y(n_422)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_410),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_373),
.A2(n_363),
.B1(n_348),
.B2(n_349),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_360),
.B(n_400),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_340),
.Y(n_426)
);

NOR2x1p5_ASAP7_75t_L g427 ( 
.A(n_337),
.B(n_270),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_340),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_356),
.B(n_317),
.Y(n_429)
);

BUFx8_ASAP7_75t_L g430 ( 
.A(n_410),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_378),
.B(n_317),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_376),
.B(n_320),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_350),
.B(n_320),
.Y(n_433)
);

NOR3xp33_ASAP7_75t_L g434 ( 
.A(n_334),
.B(n_325),
.C(n_298),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_319),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_301),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_410),
.B(n_233),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_328),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_338),
.B(n_303),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_336),
.A2(n_343),
.B1(n_344),
.B2(n_341),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_409),
.B(n_330),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_395),
.B(n_332),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_335),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_393),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_352),
.B(n_233),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_345),
.B(n_294),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_338),
.B(n_294),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_398),
.B(n_306),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_361),
.B(n_315),
.C(n_310),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_362),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_394),
.B(n_348),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_351),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_363),
.A2(n_242),
.B1(n_246),
.B2(n_307),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_377),
.Y(n_457)
);

BUFx5_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

NOR3xp33_ASAP7_75t_L g460 ( 
.A(n_399),
.B(n_307),
.C(n_323),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_353),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_326),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_354),
.B(n_266),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_355),
.B(n_366),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_366),
.B(n_283),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_366),
.B(n_266),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_392),
.B(n_159),
.Y(n_468)
);

NOR2x1p5_ASAP7_75t_L g469 ( 
.A(n_357),
.B(n_285),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_346),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_365),
.B(n_271),
.C(n_322),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_347),
.A2(n_271),
.B(n_297),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_347),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_357),
.B(n_268),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_339),
.B(n_179),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_381),
.A2(n_271),
.B(n_297),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_358),
.B(n_262),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_371),
.B(n_189),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_399),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_358),
.B(n_263),
.Y(n_480)
);

OAI221xp5_ASAP7_75t_L g481 ( 
.A1(n_368),
.A2(n_264),
.B1(n_274),
.B2(n_254),
.C(n_253),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_375),
.B(n_192),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_359),
.Y(n_483)
);

OAI221xp5_ASAP7_75t_L g484 ( 
.A1(n_369),
.A2(n_274),
.B1(n_234),
.B2(n_237),
.C(n_245),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_369),
.B(n_204),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_420),
.B(n_415),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_443),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_441),
.A2(n_242),
.B1(n_396),
.B2(n_397),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_472),
.A2(n_297),
.B(n_383),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_423),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_476),
.A2(n_389),
.B(n_401),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_440),
.B(n_412),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_423),
.B(n_211),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_471),
.A2(n_401),
.B(n_405),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_412),
.Y(n_500)
);

AO22x2_ASAP7_75t_L g501 ( 
.A1(n_454),
.A2(n_285),
.B1(n_412),
.B2(n_258),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_463),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_435),
.A2(n_439),
.B(n_442),
.C(n_477),
.Y(n_503)
);

NOR3xp33_ASAP7_75t_L g504 ( 
.A(n_452),
.B(n_201),
.C(n_227),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_426),
.B(n_217),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_450),
.B(n_448),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_428),
.B(n_218),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_455),
.A2(n_370),
.B(n_374),
.Y(n_508)
);

A2O1A1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_439),
.A2(n_248),
.B(n_239),
.C(n_255),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_425),
.B(n_220),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_414),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_225),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_455),
.A2(n_383),
.B(n_379),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_421),
.A2(n_422),
.B(n_451),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_456),
.A2(n_249),
.B1(n_256),
.B2(n_247),
.Y(n_516)
);

INVx11_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

OAI21xp33_ASAP7_75t_L g518 ( 
.A1(n_438),
.A2(n_226),
.B(n_251),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_433),
.B(n_32),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_33),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_424),
.A2(n_213),
.B1(n_321),
.B2(n_388),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_321),
.Y(n_523)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_442),
.A2(n_299),
.B(n_311),
.C(n_321),
.Y(n_524)
);

AO21x1_ASAP7_75t_L g525 ( 
.A1(n_460),
.A2(n_411),
.B(n_407),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_432),
.Y(n_526)
);

AO21x1_ASAP7_75t_L g527 ( 
.A1(n_460),
.A2(n_411),
.B(n_407),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_436),
.A2(n_321),
.B1(n_311),
.B2(n_390),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_465),
.B(n_33),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_416),
.A2(n_431),
.B(n_429),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_470),
.B(n_34),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_445),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_474),
.B(n_35),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_427),
.B(n_36),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_457),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_473),
.A2(n_98),
.B(n_40),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_447),
.B(n_37),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_446),
.B(n_48),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_479),
.B(n_52),
.Y(n_540)
);

OAI321xp33_ASAP7_75t_L g541 ( 
.A1(n_467),
.A2(n_484),
.A3(n_481),
.B1(n_466),
.B2(n_464),
.C(n_449),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_453),
.A2(n_449),
.B(n_464),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_434),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_434),
.B(n_64),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_467),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_545)
);

CKINVDCx10_ASAP7_75t_R g546 ( 
.A(n_463),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_477),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_R g548 ( 
.A(n_461),
.B(n_145),
.Y(n_548)
);

O2A1O1Ixp33_ASAP7_75t_L g549 ( 
.A1(n_485),
.A2(n_142),
.B(n_83),
.C(n_85),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_458),
.B(n_140),
.Y(n_550)
);

O2A1O1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_468),
.A2(n_91),
.B(n_93),
.C(n_96),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_458),
.B(n_480),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_458),
.B(n_482),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_503),
.A2(n_514),
.B(n_542),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_489),
.A2(n_486),
.B1(n_496),
.B2(n_520),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_547),
.A2(n_475),
.B(n_478),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_515),
.B(n_458),
.Y(n_557)
);

A2O1A1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_534),
.A2(n_469),
.B(n_463),
.C(n_108),
.Y(n_558)
);

AO31x2_ASAP7_75t_L g559 ( 
.A1(n_525),
.A2(n_527),
.A3(n_522),
.B(n_531),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_538),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_489),
.B(n_118),
.Y(n_561)
);

AND3x4_ASAP7_75t_L g562 ( 
.A(n_546),
.B(n_119),
.C(n_120),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_492),
.B(n_128),
.Y(n_563)
);

OAI21xp33_ASAP7_75t_L g564 ( 
.A1(n_509),
.A2(n_130),
.B(n_132),
.Y(n_564)
);

CKINVDCx8_ASAP7_75t_R g565 ( 
.A(n_491),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_530),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_519),
.Y(n_567)
);

AO31x2_ASAP7_75t_L g568 ( 
.A1(n_524),
.A2(n_134),
.A3(n_135),
.B(n_138),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_487),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_526),
.B(n_500),
.Y(n_570)
);

AO32x2_ASAP7_75t_L g571 ( 
.A1(n_516),
.A2(n_545),
.A3(n_548),
.B1(n_504),
.B2(n_541),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_506),
.B(n_535),
.Y(n_572)
);

AO21x1_ASAP7_75t_L g573 ( 
.A1(n_537),
.A2(n_549),
.B(n_543),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_532),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g575 ( 
.A1(n_508),
.A2(n_513),
.B(n_550),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_SL g576 ( 
.A1(n_537),
.A2(n_540),
.B(n_541),
.C(n_551),
.Y(n_576)
);

OA22x2_ASAP7_75t_L g577 ( 
.A1(n_518),
.A2(n_519),
.B1(n_501),
.B2(n_544),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_510),
.B(n_512),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_501),
.B(n_502),
.Y(n_579)
);

CKINVDCx8_ASAP7_75t_R g580 ( 
.A(n_517),
.Y(n_580)
);

NAND3x1_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_494),
.C(n_492),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_494),
.B(n_499),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_499),
.B(n_529),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_497),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_488),
.B(n_490),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_505),
.B(n_507),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_553),
.B(n_539),
.Y(n_587)
);

OAI21xp33_ASAP7_75t_SL g588 ( 
.A1(n_552),
.A2(n_548),
.B(n_523),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_533),
.B(n_536),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_533),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_536),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_486),
.B(n_406),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_528),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_486),
.B(n_406),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_492),
.B(n_494),
.Y(n_595)
);

AOI221x1_ASAP7_75t_L g596 ( 
.A1(n_504),
.A2(n_522),
.B1(n_493),
.B2(n_476),
.C(n_531),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_486),
.B(n_406),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_489),
.A2(n_456),
.B1(n_503),
.B2(n_424),
.Y(n_598)
);

NOR2x1_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_553),
.Y(n_599)
);

OAI21xp33_ASAP7_75t_L g600 ( 
.A1(n_503),
.A2(n_413),
.B(n_486),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_486),
.B(n_406),
.Y(n_601)
);

NAND2x1p5_ASAP7_75t_L g602 ( 
.A(n_492),
.B(n_494),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_499),
.Y(n_603)
);

NAND2x1_ASAP7_75t_L g604 ( 
.A(n_492),
.B(n_494),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_489),
.A2(n_190),
.B1(n_446),
.B2(n_196),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_499),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_489),
.A2(n_486),
.B1(n_496),
.B2(n_434),
.Y(n_607)
);

BUFx8_ASAP7_75t_L g608 ( 
.A(n_491),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_491),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_498),
.A2(n_495),
.B(n_476),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_486),
.B(n_452),
.C(n_496),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_491),
.B(n_415),
.Y(n_612)
);

INVx3_ASAP7_75t_SL g613 ( 
.A(n_519),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_486),
.B(n_406),
.Y(n_614)
);

AO31x2_ASAP7_75t_L g615 ( 
.A1(n_525),
.A2(n_527),
.A3(n_522),
.B(n_476),
.Y(n_615)
);

NOR2x1_ASAP7_75t_SL g616 ( 
.A(n_489),
.B(n_526),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_503),
.A2(n_472),
.B(n_514),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_511),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_503),
.A2(n_472),
.B(n_514),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_489),
.A2(n_448),
.B1(n_438),
.B2(n_331),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_486),
.B(n_406),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_511),
.Y(n_622)
);

AO31x2_ASAP7_75t_L g623 ( 
.A1(n_525),
.A2(n_527),
.A3(n_522),
.B(n_476),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_503),
.A2(n_472),
.B(n_514),
.Y(n_624)
);

AO21x2_ASAP7_75t_L g625 ( 
.A1(n_493),
.A2(n_476),
.B(n_525),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_526),
.B(n_496),
.Y(n_626)
);

AOI221x1_ASAP7_75t_L g627 ( 
.A1(n_504),
.A2(n_522),
.B1(n_493),
.B2(n_476),
.C(n_531),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_491),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_517),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_486),
.B(n_406),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_486),
.B(n_406),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_526),
.B(n_496),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_511),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_511),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_489),
.A2(n_456),
.B1(n_503),
.B2(n_424),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_491),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_486),
.B(n_406),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_491),
.B(n_415),
.Y(n_639)
);

NOR2x1_ASAP7_75t_SL g640 ( 
.A(n_557),
.B(n_609),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_608),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_611),
.A2(n_635),
.B1(n_598),
.B2(n_600),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_555),
.A2(n_605),
.B1(n_607),
.B2(n_620),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_607),
.B(n_592),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_608),
.Y(n_645)
);

OA21x2_ASAP7_75t_L g646 ( 
.A1(n_596),
.A2(n_627),
.B(n_575),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_565),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_618),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_622),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_633),
.Y(n_650)
);

CKINVDCx8_ASAP7_75t_R g651 ( 
.A(n_636),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_594),
.B(n_597),
.Y(n_652)
);

OA21x2_ASAP7_75t_L g653 ( 
.A1(n_554),
.A2(n_617),
.B(n_619),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_593),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_600),
.A2(n_577),
.B1(n_555),
.B2(n_638),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_601),
.B(n_614),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_634),
.Y(n_657)
);

AND2x2_ASAP7_75t_SL g658 ( 
.A(n_579),
.B(n_561),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_628),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_580),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_621),
.B(n_630),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_560),
.B(n_566),
.Y(n_662)
);

BUFx2_ASAP7_75t_R g663 ( 
.A(n_637),
.Y(n_663)
);

AO21x2_ASAP7_75t_L g664 ( 
.A1(n_619),
.A2(n_624),
.B(n_625),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_631),
.A2(n_578),
.B(n_558),
.C(n_572),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_574),
.A2(n_632),
.B1(n_626),
.B2(n_599),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_605),
.B(n_639),
.Y(n_667)
);

O2A1O1Ixp5_ASAP7_75t_L g668 ( 
.A1(n_576),
.A2(n_587),
.B(n_563),
.C(n_589),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_612),
.B(n_569),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_615),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_570),
.B(n_613),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_586),
.B(n_616),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_623),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_588),
.A2(n_556),
.B(n_583),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_636),
.B(n_606),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_591),
.A2(n_562),
.B1(n_581),
.B2(n_636),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_564),
.A2(n_584),
.B1(n_606),
.B2(n_603),
.Y(n_677)
);

AO21x2_ASAP7_75t_L g678 ( 
.A1(n_585),
.A2(n_571),
.B(n_588),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_603),
.A2(n_604),
.B(n_582),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_629),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_595),
.A2(n_602),
.B(n_623),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_568),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_590),
.A2(n_571),
.B(n_559),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_559),
.Y(n_685)
);

OAI21x1_ASAP7_75t_SL g686 ( 
.A1(n_571),
.A2(n_568),
.B(n_623),
.Y(n_686)
);

OA21x2_ASAP7_75t_L g687 ( 
.A1(n_596),
.A2(n_627),
.B(n_610),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_591),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_555),
.A2(n_607),
.B1(n_448),
.B2(n_489),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_580),
.Y(n_690)
);

OAI222xp33_ASAP7_75t_L g691 ( 
.A1(n_605),
.A2(n_607),
.B1(n_577),
.B2(n_555),
.C1(n_635),
.C2(n_598),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_636),
.B(n_492),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_611),
.A2(n_635),
.B1(n_598),
.B2(n_600),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_636),
.B(n_492),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_555),
.A2(n_605),
.B1(n_489),
.B2(n_456),
.Y(n_695)
);

OA21x2_ASAP7_75t_L g696 ( 
.A1(n_596),
.A2(n_627),
.B(n_610),
.Y(n_696)
);

AO31x2_ASAP7_75t_L g697 ( 
.A1(n_596),
.A2(n_627),
.A3(n_573),
.B(n_527),
.Y(n_697)
);

NAND2x1p5_ASAP7_75t_L g698 ( 
.A(n_636),
.B(n_492),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_595),
.Y(n_699)
);

NAND2x1p5_ASAP7_75t_L g700 ( 
.A(n_636),
.B(n_492),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_607),
.B(n_611),
.Y(n_701)
);

BUFx2_ASAP7_75t_SL g702 ( 
.A(n_580),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_629),
.B(n_423),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_593),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_701),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_667),
.B(n_671),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_648),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_704),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_682),
.B(n_654),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_649),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_650),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_704),
.B(n_662),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_652),
.B(n_656),
.Y(n_713)
);

AO21x2_ASAP7_75t_L g714 ( 
.A1(n_686),
.A2(n_684),
.B(n_683),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_665),
.A2(n_644),
.B(n_693),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_661),
.B(n_695),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_704),
.Y(n_717)
);

BUFx16f_ASAP7_75t_R g718 ( 
.A(n_675),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_657),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_643),
.A2(n_658),
.B1(n_640),
.B2(n_676),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_704),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_660),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_670),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_659),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_670),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_689),
.A2(n_658),
.B1(n_666),
.B2(n_662),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_689),
.B(n_655),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_688),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_663),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_673),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_642),
.A2(n_672),
.B1(n_647),
.B2(n_685),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_688),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_651),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_668),
.A2(n_691),
.B(n_674),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_675),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_653),
.B(n_664),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_653),
.B(n_664),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_692),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_669),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_647),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_641),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_680),
.B(n_672),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_699),
.B(n_675),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_703),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_687),
.Y(n_745)
);

HB1xp67_ASAP7_75t_SL g746 ( 
.A(n_702),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_692),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_685),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_694),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_736),
.B(n_646),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_736),
.B(n_646),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_748),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_737),
.B(n_646),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_737),
.B(n_696),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_716),
.B(n_691),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_725),
.Y(n_757)
);

BUFx4f_ASAP7_75t_L g758 ( 
.A(n_712),
.Y(n_758)
);

INVxp33_ASAP7_75t_L g759 ( 
.A(n_712),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_705),
.B(n_697),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_726),
.A2(n_677),
.B1(n_678),
.B2(n_645),
.Y(n_761)
);

AND2x4_ASAP7_75t_SL g762 ( 
.A(n_735),
.B(n_749),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_722),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_727),
.B(n_730),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_712),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_715),
.B(n_739),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_755),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_750),
.B(n_714),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_750),
.B(n_709),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_755),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_750),
.B(n_714),
.Y(n_771)
);

NOR2x1_ASAP7_75t_L g772 ( 
.A(n_765),
.B(n_721),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_766),
.B(n_745),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_756),
.B(n_707),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_760),
.B(n_707),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_751),
.B(n_753),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_756),
.B(n_710),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_762),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_766),
.B(n_710),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_757),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_765),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_766),
.B(n_711),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_751),
.B(n_714),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_751),
.B(n_714),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_774),
.B(n_753),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_776),
.B(n_753),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_767),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_779),
.B(n_764),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_780),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_768),
.B(n_754),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_777),
.B(n_729),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_782),
.B(n_773),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_773),
.B(n_764),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_768),
.B(n_764),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_770),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_769),
.B(n_752),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_778),
.B(n_741),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_771),
.B(n_754),
.Y(n_798)
);

AOI211xp5_ASAP7_75t_L g799 ( 
.A1(n_791),
.A2(n_778),
.B(n_759),
.C(n_734),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_785),
.B(n_728),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_792),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_786),
.B(n_771),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_792),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_790),
.B(n_783),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_787),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_787),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_796),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_L g808 ( 
.A1(n_797),
.A2(n_706),
.B(n_740),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_796),
.B(n_769),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_790),
.B(n_783),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_796),
.A2(n_720),
.B1(n_761),
.B2(n_769),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_798),
.B(n_784),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_801),
.Y(n_813)
);

OAI32xp33_ASAP7_75t_L g814 ( 
.A1(n_803),
.A2(n_759),
.A3(n_794),
.B1(n_793),
.B2(n_786),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_799),
.A2(n_772),
.B1(n_758),
.B2(n_789),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_805),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_806),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_811),
.A2(n_772),
.B1(n_758),
.B2(n_794),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_804),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_802),
.B(n_798),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_802),
.B(n_800),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_L g822 ( 
.A1(n_807),
.A2(n_765),
.B1(n_781),
.B2(n_793),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_SL g823 ( 
.A1(n_800),
.A2(n_762),
.B1(n_765),
.B2(n_732),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_821),
.B(n_724),
.Y(n_824)
);

OAI322xp33_ASAP7_75t_L g825 ( 
.A1(n_818),
.A2(n_812),
.A3(n_810),
.B1(n_788),
.B2(n_724),
.C1(n_775),
.C2(n_795),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_816),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_823),
.B(n_809),
.Y(n_827)
);

XNOR2xp5_ASAP7_75t_L g828 ( 
.A(n_823),
.B(n_763),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_828),
.A2(n_814),
.B(n_815),
.Y(n_829)
);

AOI32xp33_ASAP7_75t_L g830 ( 
.A1(n_827),
.A2(n_822),
.A3(n_807),
.B1(n_813),
.B2(n_809),
.Y(n_830)
);

AOI21xp33_ASAP7_75t_SL g831 ( 
.A1(n_824),
.A2(n_808),
.B(n_660),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_829),
.B(n_819),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_831),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_833),
.B(n_826),
.Y(n_834)
);

NOR2x1_ASAP7_75t_L g835 ( 
.A(n_833),
.B(n_733),
.Y(n_835)
);

NAND4xp75_ASAP7_75t_L g836 ( 
.A(n_835),
.B(n_832),
.C(n_746),
.D(n_830),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_834),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_L g838 ( 
.A(n_837),
.B(n_832),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_836),
.B(n_690),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_838),
.A2(n_690),
.B(n_681),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_839),
.Y(n_841)
);

OAI221xp5_ASAP7_75t_L g842 ( 
.A1(n_838),
.A2(n_733),
.B1(n_681),
.B2(n_703),
.C(n_744),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_841),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_840),
.A2(n_825),
.B1(n_817),
.B2(n_733),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_842),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_841),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_841),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_843),
.B(n_711),
.Y(n_848)
);

AOI22x1_ASAP7_75t_L g849 ( 
.A1(n_846),
.A2(n_700),
.B1(n_698),
.B2(n_694),
.Y(n_849)
);

OAI32xp33_ASAP7_75t_L g850 ( 
.A1(n_846),
.A2(n_700),
.A3(n_698),
.B1(n_721),
.B2(n_713),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_847),
.A2(n_820),
.B1(n_703),
.B2(n_731),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_845),
.Y(n_852)
);

AO22x1_ASAP7_75t_L g853 ( 
.A1(n_844),
.A2(n_699),
.B1(n_721),
.B2(n_708),
.Y(n_853)
);

AO22x2_ASAP7_75t_SL g854 ( 
.A1(n_843),
.A2(n_717),
.B1(n_719),
.B2(n_718),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_848),
.A2(n_849),
.B1(n_851),
.B2(n_852),
.Y(n_855)
);

XNOR2xp5_ASAP7_75t_L g856 ( 
.A(n_853),
.B(n_742),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_854),
.A2(n_809),
.B1(n_721),
.B2(n_747),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_850),
.A2(n_708),
.B(n_747),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_SL g859 ( 
.A1(n_856),
.A2(n_717),
.B(n_743),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_855),
.A2(n_858),
.B(n_857),
.Y(n_860)
);

OA21x2_ASAP7_75t_L g861 ( 
.A1(n_860),
.A2(n_719),
.B(n_679),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_861),
.B(n_859),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_862),
.A2(n_738),
.B1(n_717),
.B2(n_749),
.Y(n_863)
);


endmodule