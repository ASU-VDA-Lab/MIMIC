module fake_jpeg_22802_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_SL g19 ( 
.A(n_18),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_9),
.B1(n_14),
.B2(n_11),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_34),
.B1(n_19),
.B2(n_13),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_17),
.B1(n_12),
.B2(n_9),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_19),
.B1(n_10),
.B2(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_17),
.B1(n_12),
.B2(n_18),
.Y(n_34)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_45),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_24),
.B1(n_25),
.B2(n_23),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_19),
.B1(n_41),
.B2(n_27),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_24),
.C(n_26),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_21),
.Y(n_54)
);

OAI22x1_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_30),
.B1(n_13),
.B2(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

OR2x4_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_25),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_27),
.B(n_15),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_42),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_53),
.B1(n_30),
.B2(n_37),
.Y(n_64)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_54),
.B(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_38),
.B(n_40),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_64),
.B(n_65),
.Y(n_67)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_49),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_70),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_53),
.B1(n_52),
.B2(n_46),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_75),
.B1(n_42),
.B2(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_47),
.B1(n_55),
.B2(n_49),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_46),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_62),
.C(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_83),
.C(n_76),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_50),
.B(n_66),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_84),
.B(n_42),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_64),
.C(n_63),
.Y(n_83)
);

BUFx12f_ASAP7_75t_SL g85 ( 
.A(n_81),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_78),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_28),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_36),
.C(n_35),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_84),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_58),
.B1(n_61),
.B2(n_28),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_94),
.B(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_58),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_97),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_95),
.C(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_100),
.B(n_101),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.C(n_1),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_103),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_106)
);

AOI321xp33_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_93),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);


endmodule