module fake_netlist_1_11138_n_28 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
NOR2xp33_ASAP7_75t_R g12 ( .A(n_9), .B(n_3), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_0), .B(n_3), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_13), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_16), .B(n_1), .C(n_2), .Y(n_19) );
INVxp67_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
AOI221xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_19), .B1(n_16), .B2(n_17), .C(n_15), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_14), .B(n_12), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_19), .B1(n_14), .B2(n_12), .Y(n_23) );
NOR4xp25_ASAP7_75t_L g24 ( .A(n_23), .B(n_1), .C(n_2), .D(n_4), .Y(n_24) );
NAND5xp2_ASAP7_75t_L g25 ( .A(n_23), .B(n_4), .C(n_6), .D(n_7), .E(n_8), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_6), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI222xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_26), .B1(n_25), .B2(n_24), .C1(n_11), .C2(n_10), .Y(n_28) );
endmodule