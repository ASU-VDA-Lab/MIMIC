module fake_jpeg_13877_n_521 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_521);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_521;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_62),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_63),
.Y(n_189)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_65),
.Y(n_200)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_68),
.Y(n_164)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_72),
.Y(n_175)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_73),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_74),
.B(n_84),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g186 ( 
.A(n_78),
.Y(n_186)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_79),
.Y(n_199)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_16),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_86),
.B(n_91),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_90),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_0),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_92),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_25),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_93),
.A2(n_113),
.B1(n_41),
.B2(n_34),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_18),
.B(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_115),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_105),
.Y(n_145)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

NAND2x1_ASAP7_75t_SL g158 ( 
.A(n_107),
.B(n_110),
.Y(n_158)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_46),
.B(n_5),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_27),
.C(n_57),
.Y(n_134)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_46),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_38),
.B(n_5),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_119),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_120),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_118),
.B(n_48),
.Y(n_190)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_38),
.B(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_122),
.Y(n_162)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

NAND2x1p5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_55),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_133),
.B(n_164),
.C(n_182),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_134),
.B(n_169),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_53),
.B1(n_43),
.B2(n_57),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_136),
.A2(n_154),
.B1(n_160),
.B2(n_48),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_95),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_143),
.A2(n_144),
.B1(n_155),
.B2(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_43),
.B1(n_27),
.B2(n_42),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_56),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_148),
.B(n_150),
.C(n_180),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_80),
.B(n_40),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_58),
.A2(n_42),
.B1(n_34),
.B2(n_47),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_69),
.A2(n_55),
.B1(n_50),
.B2(n_28),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_157),
.A2(n_181),
.B(n_192),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_99),
.A2(n_47),
.B1(n_45),
.B2(n_41),
.Y(n_160)
);

CKINVDCx12_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_161),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_45),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_163),
.B(n_173),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_59),
.A2(n_40),
.B1(n_28),
.B2(n_29),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_101),
.B(n_6),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_60),
.B(n_100),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_62),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_174),
.A2(n_178),
.B1(n_185),
.B2(n_123),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_63),
.A2(n_33),
.B1(n_36),
.B2(n_48),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_106),
.B(n_6),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_72),
.A2(n_111),
.B1(n_81),
.B2(n_88),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_65),
.B(n_7),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_196),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_104),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_120),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_67),
.A2(n_33),
.B1(n_36),
.B2(n_26),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_190),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_117),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_75),
.B(n_10),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_77),
.B(n_10),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_141),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_203),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_140),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_204),
.B(n_216),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_143),
.A2(n_85),
.B1(n_89),
.B2(n_87),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_206),
.A2(n_213),
.B1(n_235),
.B2(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_208),
.Y(n_313)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_94),
.B1(n_92),
.B2(n_90),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_212),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_154),
.A2(n_110),
.B1(n_105),
.B2(n_78),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_194),
.A2(n_48),
.B1(n_26),
.B2(n_36),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_125),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_124),
.B1(n_142),
.B2(n_133),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_217),
.A2(n_220),
.B1(n_239),
.B2(n_243),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_246),
.Y(n_289)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_26),
.B1(n_36),
.B2(n_48),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_221),
.Y(n_277)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_137),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_225),
.B(n_248),
.Y(n_278)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_226),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_227),
.B(n_240),
.Y(n_286)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_229),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_12),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_232),
.B(n_249),
.C(n_253),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_149),
.A2(n_26),
.B1(n_13),
.B2(n_14),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_234),
.A2(n_237),
.B1(n_255),
.B2(n_270),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_131),
.A2(n_26),
.B1(n_13),
.B2(n_14),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_126),
.Y(n_236)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_149),
.A2(n_12),
.B1(n_14),
.B2(n_158),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_181),
.A2(n_157),
.B1(n_169),
.B2(n_153),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_138),
.B(n_186),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_126),
.Y(n_242)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_201),
.B1(n_179),
.B2(n_151),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_245),
.B(n_259),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_167),
.B(n_135),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_258),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_186),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_130),
.B(n_178),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_193),
.A2(n_201),
.B1(n_179),
.B2(n_151),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_141),
.A2(n_129),
.B1(n_168),
.B2(n_200),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_260),
.B1(n_248),
.B2(n_209),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_252),
.B(n_223),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_156),
.B(n_197),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_257),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_129),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_166),
.B(n_171),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_186),
.B(n_164),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_168),
.A2(n_189),
.B1(n_200),
.B2(n_176),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_156),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_262),
.Y(n_315)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_189),
.A2(n_132),
.B1(n_176),
.B2(n_139),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_263),
.A2(n_266),
.B1(n_268),
.B2(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_264),
.B(n_267),
.Y(n_316)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_265),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_139),
.A2(n_171),
.B1(n_202),
.B2(n_158),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_123),
.B(n_191),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_232),
.C(n_270),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_147),
.A2(n_187),
.B(n_145),
.C(n_137),
.Y(n_269)
);

AO22x2_ASAP7_75t_L g314 ( 
.A1(n_269),
.A2(n_261),
.B1(n_265),
.B2(n_242),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_228),
.A2(n_187),
.B1(n_191),
.B2(n_145),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_280),
.B1(n_297),
.B2(n_302),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_228),
.A2(n_191),
.B1(n_233),
.B2(n_246),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_205),
.B(n_245),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_300),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g296 ( 
.A1(n_231),
.A2(n_211),
.A3(n_249),
.B1(n_205),
.B2(n_217),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_317),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_233),
.A2(n_211),
.B1(n_252),
.B2(n_212),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_232),
.B(n_247),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_239),
.A2(n_249),
.B1(n_258),
.B2(n_223),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_291),
.C(n_307),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_238),
.A2(n_223),
.B1(n_219),
.B2(n_226),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_302),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_SL g346 ( 
.A1(n_309),
.A2(n_299),
.B(n_273),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_266),
.A2(n_263),
.B1(n_262),
.B2(n_254),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_311),
.A2(n_318),
.B1(n_321),
.B2(n_275),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_253),
.B(n_268),
.CI(n_269),
.CON(n_312),
.SN(n_312)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_312),
.B(n_321),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_312),
.Y(n_344)
);

OAI32xp33_ASAP7_75t_L g317 ( 
.A1(n_207),
.A2(n_214),
.A3(n_229),
.B1(n_222),
.B2(n_236),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_221),
.A2(n_255),
.B1(n_264),
.B2(n_257),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_225),
.A2(n_244),
.B1(n_267),
.B2(n_253),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_224),
.B(n_230),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_323),
.A2(n_326),
.B(n_339),
.Y(n_365)
);

BUFx12_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

INVx13_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_299),
.A2(n_256),
.B(n_275),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_308),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_327),
.B(n_338),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_331),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_281),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g377 ( 
.A1(n_332),
.A2(n_344),
.B(n_355),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_316),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_358),
.Y(n_366)
);

BUFx24_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

INVx13_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_335),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_293),
.C(n_310),
.Y(n_373)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_284),
.Y(n_338)
);

A2O1A1O1Ixp25_ASAP7_75t_L g339 ( 
.A1(n_305),
.A2(n_300),
.B(n_271),
.C(n_304),
.D(n_296),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_285),
.B(n_278),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_340),
.B(n_342),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_271),
.B(n_305),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_343),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_280),
.Y(n_343)
);

BUFx24_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_345),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_348),
.B1(n_351),
.B2(n_359),
.Y(n_381)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_279),
.A2(n_289),
.B1(n_306),
.B2(n_303),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_298),
.B(n_319),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_349),
.B(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_279),
.B(n_289),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_289),
.A2(n_287),
.B1(n_288),
.B2(n_314),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_282),
.B(n_283),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_357),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_354),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_283),
.A2(n_319),
.B(n_298),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_360),
.Y(n_384)
);

A2O1A1O1Ixp25_ASAP7_75t_L g357 ( 
.A1(n_315),
.A2(n_314),
.B(n_301),
.C(n_320),
.D(n_294),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_318),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_314),
.A2(n_274),
.B1(n_295),
.B2(n_277),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_314),
.A2(n_294),
.B(n_320),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_329),
.A2(n_274),
.B1(n_295),
.B2(n_293),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_367),
.A2(n_374),
.B1(n_392),
.B2(n_351),
.Y(n_406)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_322),
.C(n_323),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_329),
.A2(n_272),
.B1(n_310),
.B2(n_350),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_272),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_379),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_338),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

OA22x2_ASAP7_75t_L g383 ( 
.A1(n_345),
.A2(n_344),
.B1(n_343),
.B2(n_358),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_390),
.Y(n_398)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_334),
.Y(n_387)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

CKINVDCx12_ASAP7_75t_R g388 ( 
.A(n_334),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_388),
.Y(n_418)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_344),
.A2(n_332),
.B1(n_325),
.B2(n_360),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_394),
.C(n_399),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_336),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_328),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_341),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_330),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_401),
.C(n_403),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_330),
.C(n_339),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_339),
.C(n_348),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_333),
.Y(n_404)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_404),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_363),
.B(n_327),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_407),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_406),
.A2(n_361),
.B1(n_372),
.B2(n_383),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_340),
.C(n_345),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_381),
.A2(n_325),
.B1(n_355),
.B2(n_346),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_412),
.B1(n_417),
.B2(n_392),
.Y(n_421)
);

XOR2x1_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_357),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_410),
.B(n_375),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_381),
.A2(n_352),
.B1(n_326),
.B2(n_357),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_342),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_361),
.C(n_383),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_384),
.A2(n_334),
.B(n_359),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_415),
.A2(n_419),
.B(n_398),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_366),
.B(n_331),
.Y(n_416)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_416),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_378),
.A2(n_382),
.B1(n_389),
.B2(n_369),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_421),
.A2(n_423),
.B1(n_436),
.B2(n_406),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_416),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_422),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_409),
.A2(n_374),
.B1(n_369),
.B2(n_378),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_404),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_432),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_408),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_412),
.B(n_383),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_433),
.B(n_437),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_386),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_L g450 ( 
.A1(n_434),
.A2(n_438),
.B(n_443),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_377),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_414),
.Y(n_445)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_439),
.B(n_435),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_372),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_396),
.C(n_419),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_393),
.B(n_387),
.C(n_385),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_410),
.C(n_415),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_442),
.A2(n_398),
.B(n_411),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_452),
.C(n_453),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_448),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_455),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_449),
.A2(n_451),
.B1(n_433),
.B2(n_443),
.Y(n_469)
);

XNOR2x1_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_403),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_429),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_429),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_454),
.A2(n_434),
.B(n_437),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_401),
.C(n_394),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_399),
.C(n_417),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_456),
.A2(n_458),
.B1(n_460),
.B2(n_430),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_387),
.C(n_385),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_367),
.C(n_413),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_388),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_461),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_449),
.A2(n_436),
.B1(n_425),
.B2(n_422),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_463),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_459),
.A2(n_423),
.B1(n_425),
.B2(n_427),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_472),
.B1(n_460),
.B2(n_413),
.Y(n_484)
);

AO221x1_ASAP7_75t_L g468 ( 
.A1(n_457),
.A2(n_440),
.B1(n_432),
.B2(n_426),
.C(n_420),
.Y(n_468)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_468),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_470),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_473),
.B(n_444),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_457),
.A2(n_428),
.B1(n_438),
.B2(n_420),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_454),
.A2(n_428),
.B(n_433),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_450),
.A2(n_461),
.B1(n_433),
.B2(n_462),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_474),
.Y(n_487)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_477),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_453),
.C(n_452),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_479),
.B(n_480),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_455),
.C(n_458),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_467),
.B(n_456),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_482),
.A2(n_467),
.B(n_480),
.Y(n_493)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_451),
.C(n_448),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_445),
.C(n_471),
.Y(n_498)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_488),
.A2(n_474),
.B(n_463),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_465),
.C(n_469),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_491),
.A2(n_496),
.B(n_483),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_493),
.A2(n_497),
.B(n_499),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_487),
.A2(n_477),
.B1(n_464),
.B2(n_476),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_498),
.C(n_489),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_478),
.A2(n_466),
.B1(n_468),
.B2(n_464),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_371),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_473),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_395),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_501),
.B(n_502),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_486),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_504),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_485),
.C(n_478),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_497),
.A2(n_371),
.B(n_376),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_506),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_337),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_371),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_507),
.A2(n_499),
.B(n_496),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_510),
.A2(n_391),
.B(n_324),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_513),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_364),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_509),
.A2(n_364),
.B(n_370),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_515),
.B(n_514),
.Y(n_518)
);

O2A1O1Ixp33_ASAP7_75t_SL g517 ( 
.A1(n_516),
.A2(n_512),
.B(n_391),
.C(n_324),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_517),
.A2(n_518),
.B1(n_391),
.B2(n_324),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_510),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_508),
.Y(n_521)
);


endmodule