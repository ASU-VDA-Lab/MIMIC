module fake_jpeg_720_n_222 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_222);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_12),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_1),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_87),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_73),
.B(n_67),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_75),
.CI(n_74),
.CON(n_105),
.SN(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_75),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_55),
.B1(n_69),
.B2(n_74),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_108),
.B1(n_114),
.B2(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_64),
.B1(n_52),
.B2(n_63),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_101),
.B1(n_107),
.B2(n_94),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_63),
.B1(n_54),
.B2(n_59),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_114),
.B(n_94),
.C(n_53),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_111),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_52),
.B1(n_54),
.B2(n_71),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_73),
.B1(n_69),
.B2(n_55),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_59),
.B1(n_65),
.B2(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_93),
.Y(n_117)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_115),
.Y(n_125)
);

OR2x4_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_74),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_62),
.C(n_60),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_118),
.B1(n_120),
.B2(n_136),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_126),
.C(n_133),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_65),
.B1(n_72),
.B2(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_27),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_97),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_53),
.B1(n_2),
.B2(n_4),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_131),
.B1(n_51),
.B2(n_30),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_113),
.B1(n_102),
.B2(n_109),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_53),
.B(n_5),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_8),
.B(n_9),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_25),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_13),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_7),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_7),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_143),
.Y(n_172)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_158),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_148),
.B1(n_17),
.B2(n_19),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_147),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_155),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_10),
.B(n_11),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_154),
.B(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_14),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_157),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_164),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_135),
.B1(n_136),
.B2(n_134),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_35),
.C(n_47),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_177),
.C(n_178),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_33),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_154),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_31),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_44),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_49),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_32),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_146),
.B(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_145),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_191),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_148),
.B(n_37),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_188),
.Y(n_195)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_190),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_40),
.B(n_41),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_43),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_193),
.C(n_178),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_203),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_160),
.B1(n_165),
.B2(n_174),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_169),
.B1(n_188),
.B2(n_177),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_181),
.C(n_167),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_166),
.C(n_45),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_208),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_181),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_186),
.B(n_189),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_209),
.B(n_210),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_204),
.A2(n_196),
.B1(n_195),
.B2(n_201),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_199),
.B1(n_198),
.B2(n_194),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_206),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_216),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_199),
.CI(n_211),
.CON(n_218),
.SN(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_211),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_219),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_221),
.A2(n_217),
.B(n_214),
.Y(n_222)
);


endmodule