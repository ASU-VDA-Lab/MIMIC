module real_aes_10453_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g1160 ( .A(n_0), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_1), .A2(n_65), .B1(n_558), .B2(n_560), .Y(n_1384) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1), .Y(n_1414) );
AO22x2_ASAP7_75t_L g865 ( .A1(n_2), .A2(n_866), .B1(n_909), .B2(n_910), .Y(n_865) );
INVxp67_ASAP7_75t_L g909 ( .A(n_2), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_3), .A2(n_194), .B1(n_688), .B2(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g735 ( .A(n_3), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g1037 ( .A(n_4), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_5), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_5), .B(n_176), .Y(n_369) );
AND2x2_ASAP7_75t_L g379 ( .A(n_5), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g407 ( .A(n_5), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_6), .A2(n_132), .B1(n_331), .B2(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g433 ( .A(n_6), .Y(n_433) );
INVx1_ASAP7_75t_L g828 ( .A(n_7), .Y(n_828) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_7), .A2(n_118), .B1(n_576), .B2(n_854), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_8), .Y(n_701) );
INVx1_ASAP7_75t_L g1259 ( .A(n_9), .Y(n_1259) );
XNOR2x2_ASAP7_75t_L g766 ( .A(n_10), .B(n_767), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g999 ( .A(n_11), .Y(n_999) );
AOI21xp33_ASAP7_75t_L g783 ( .A1(n_12), .A2(n_527), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g810 ( .A(n_12), .Y(n_810) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_13), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_13), .A2(n_213), .B1(n_842), .B2(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g511 ( .A(n_14), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_14), .A2(n_173), .B1(n_562), .B2(n_563), .Y(n_561) );
XNOR2xp5_ASAP7_75t_L g568 ( .A(n_15), .B(n_569), .Y(n_568) );
AO221x2_ASAP7_75t_L g1186 ( .A1(n_15), .A2(n_49), .B1(n_1158), .B2(n_1177), .C(n_1187), .Y(n_1186) );
AO22x2_ASAP7_75t_L g1084 ( .A1(n_16), .A2(n_1085), .B1(n_1086), .B2(n_1137), .Y(n_1084) );
INVxp67_ASAP7_75t_SL g1085 ( .A(n_16), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_17), .A2(n_42), .B1(n_642), .B2(n_645), .Y(n_704) );
INVx1_ASAP7_75t_L g757 ( .A(n_17), .Y(n_757) );
INVx1_ASAP7_75t_L g1205 ( .A(n_18), .Y(n_1205) );
OR2x2_ASAP7_75t_L g275 ( .A(n_19), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g314 ( .A(n_19), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_20), .A2(n_139), .B1(n_794), .B2(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g806 ( .A(n_20), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_21), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_22), .A2(n_71), .B1(n_596), .B2(n_836), .Y(n_835) );
INVxp33_ASAP7_75t_L g861 ( .A(n_22), .Y(n_861) );
INVx1_ASAP7_75t_L g1188 ( .A(n_23), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_24), .A2(n_189), .B1(n_562), .B2(n_563), .Y(n_1386) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_24), .A2(n_189), .B1(n_441), .B2(n_795), .Y(n_1420) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_25), .Y(n_303) );
INVx1_ASAP7_75t_L g277 ( .A(n_26), .Y(n_277) );
BUFx2_ASAP7_75t_L g329 ( .A(n_26), .Y(n_329) );
BUFx2_ASAP7_75t_L g351 ( .A(n_26), .Y(n_351) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_26), .B(n_369), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_27), .A2(n_169), .B1(n_532), .B2(n_598), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_27), .A2(n_169), .B1(n_665), .B2(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g582 ( .A(n_28), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_28), .A2(n_168), .B1(n_596), .B2(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g1257 ( .A(n_29), .Y(n_1257) );
INVx1_ASAP7_75t_L g825 ( .A(n_30), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_30), .A2(n_58), .B1(n_337), .B2(n_846), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g874 ( .A1(n_31), .A2(n_201), .B1(n_576), .B2(n_875), .C(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g883 ( .A(n_31), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_32), .A2(n_54), .B1(n_250), .B2(n_519), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_32), .A2(n_146), .B1(n_672), .B2(n_673), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_33), .A2(n_39), .B1(n_375), .B2(n_416), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_33), .A2(n_39), .B1(n_343), .B2(n_588), .C(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_34), .A2(n_61), .B1(n_1121), .B2(n_1124), .Y(n_1123) );
INVxp67_ASAP7_75t_SL g1129 ( .A(n_34), .Y(n_1129) );
INVx1_ASAP7_75t_L g952 ( .A(n_35), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_35), .A2(n_52), .B1(n_979), .B2(n_981), .Y(n_978) );
CKINVDCx16_ASAP7_75t_R g1202 ( .A(n_36), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_37), .A2(n_195), .B1(n_586), .B2(n_588), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_37), .A2(n_195), .B1(n_603), .B2(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g1253 ( .A(n_38), .Y(n_1253) );
XNOR2xp5_ASAP7_75t_L g1375 ( .A(n_38), .B(n_1376), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_38), .A2(n_1429), .B1(n_1433), .B2(n_1437), .Y(n_1428) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_40), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_41), .A2(n_229), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_41), .A2(n_229), .B1(n_551), .B2(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g696 ( .A(n_42), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_43), .A2(n_73), .B1(n_596), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_43), .A2(n_73), .B1(n_842), .B2(n_843), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_44), .Y(n_717) );
INVx1_ASAP7_75t_L g462 ( .A(n_45), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_45), .A2(n_124), .B1(n_537), .B2(n_540), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_46), .A2(n_196), .B1(n_479), .B2(n_576), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_46), .A2(n_196), .B1(n_505), .B2(n_620), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_47), .Y(n_773) );
INVx1_ASAP7_75t_L g287 ( .A(n_48), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_48), .A2(n_50), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_397) );
INVx1_ASAP7_75t_L g278 ( .A(n_50), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_51), .A2(n_85), .B1(n_603), .B2(n_838), .Y(n_837) );
INVxp67_ASAP7_75t_SL g852 ( .A(n_51), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g955 ( .A1(n_52), .A2(n_63), .B1(n_603), .B2(n_838), .C(n_956), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_53), .A2(n_122), .B1(n_562), .B2(n_563), .Y(n_932) );
INVx1_ASAP7_75t_L g969 ( .A(n_53), .Y(n_969) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_54), .A2(n_192), .B1(n_642), .B2(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g475 ( .A(n_55), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_55), .A2(n_103), .B1(n_542), .B2(n_545), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g1109 ( .A1(n_56), .A2(n_101), .B1(n_530), .B2(n_1110), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_56), .A2(n_101), .B1(n_1121), .B2(n_1122), .Y(n_1120) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_57), .Y(n_779) );
INVxp33_ASAP7_75t_L g822 ( .A(n_58), .Y(n_822) );
INVx1_ASAP7_75t_L g1216 ( .A(n_59), .Y(n_1216) );
CKINVDCx16_ASAP7_75t_R g1221 ( .A(n_60), .Y(n_1221) );
INVxp33_ASAP7_75t_L g1136 ( .A(n_61), .Y(n_1136) );
INVx1_ASAP7_75t_L g991 ( .A(n_62), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g1054 ( .A1(n_62), .A2(n_113), .B1(n_1055), .B2(n_1056), .C(n_1058), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_63), .A2(n_174), .B1(n_280), .B2(n_977), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g1393 ( .A(n_64), .Y(n_1393) );
INVx1_ASAP7_75t_L g1411 ( .A(n_65), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_66), .A2(n_208), .B1(n_289), .B2(n_670), .Y(n_1385) );
OAI211xp5_ASAP7_75t_SL g1397 ( .A1(n_66), .A2(n_375), .B(n_1398), .C(n_1407), .Y(n_1397) );
INVx1_ASAP7_75t_L g881 ( .A(n_67), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_67), .A2(n_184), .B1(n_298), .B2(n_902), .Y(n_908) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_68), .Y(n_1095) );
AOI22xp33_ASAP7_75t_SL g1113 ( .A1(n_68), .A2(n_97), .B1(n_528), .B2(n_1110), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_69), .A2(n_191), .B1(n_596), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_69), .A2(n_191), .B1(n_842), .B2(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g1166 ( .A(n_70), .Y(n_1166) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_71), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_72), .A2(n_107), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_72), .A2(n_107), .B1(n_598), .B2(n_607), .Y(n_661) );
XNOR2x2_ASAP7_75t_L g453 ( .A(n_74), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g636 ( .A(n_75), .Y(n_636) );
OAI222xp33_ASAP7_75t_L g649 ( .A1(n_75), .A2(n_146), .B1(n_159), .B2(n_650), .C1(n_651), .C2(n_652), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_76), .A2(n_102), .B1(n_562), .B2(n_563), .Y(n_1126) );
INVxp33_ASAP7_75t_SL g1133 ( .A(n_76), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_77), .A2(n_138), .B1(n_347), .B2(n_349), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_77), .A2(n_138), .B1(n_441), .B2(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g1390 ( .A(n_78), .Y(n_1390) );
AOI221xp5_ASAP7_75t_L g1404 ( .A1(n_78), .A2(n_153), .B1(n_497), .B2(n_956), .C(n_1405), .Y(n_1404) );
CKINVDCx16_ASAP7_75t_R g1223 ( .A(n_79), .Y(n_1223) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_80), .A2(n_121), .B1(n_1171), .B2(n_1174), .Y(n_1183) );
INVx1_ASAP7_75t_L g1021 ( .A(n_81), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_81), .A2(n_230), .B1(n_1072), .B2(n_1074), .Y(n_1071) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_82), .Y(n_728) );
INVx1_ASAP7_75t_L g276 ( .A(n_83), .Y(n_276) );
INVx1_ASAP7_75t_L g327 ( .A(n_83), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_84), .A2(n_135), .B1(n_588), .B2(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g626 ( .A(n_84), .Y(n_626) );
INVxp33_ASAP7_75t_L g858 ( .A(n_85), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_86), .A2(n_88), .B1(n_318), .B2(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g958 ( .A(n_86), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_87), .A2(n_114), .B1(n_332), .B2(n_347), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_87), .A2(n_114), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g960 ( .A(n_88), .Y(n_960) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_89), .Y(n_725) );
INVx1_ASAP7_75t_L g1204 ( .A(n_90), .Y(n_1204) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_91), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_92), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_93), .A2(n_152), .B1(n_553), .B2(n_665), .Y(n_1383) );
INVx1_ASAP7_75t_L g1416 ( .A(n_93), .Y(n_1416) );
INVx1_ASAP7_75t_L g572 ( .A(n_94), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_94), .A2(n_164), .B1(n_530), .B2(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g937 ( .A(n_95), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g961 ( .A1(n_95), .A2(n_416), .B1(n_438), .B2(n_962), .C(n_965), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_96), .B(n_640), .Y(n_703) );
INVx1_ASAP7_75t_L g755 ( .A(n_96), .Y(n_755) );
INVxp33_ASAP7_75t_SL g1089 ( .A(n_97), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_98), .A2(n_225), .B1(n_603), .B2(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_98), .A2(n_225), .B1(n_574), .B2(n_586), .Y(n_844) );
AO221x2_ASAP7_75t_L g1151 ( .A1(n_99), .A2(n_156), .B1(n_1152), .B2(n_1158), .C(n_1159), .Y(n_1151) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_100), .Y(n_316) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_102), .Y(n_1134) );
INVx1_ASAP7_75t_L g457 ( .A(n_103), .Y(n_457) );
INVx1_ASAP7_75t_L g241 ( .A(n_104), .Y(n_241) );
OA22x2_ASAP7_75t_L g682 ( .A1(n_105), .A2(n_683), .B1(n_764), .B2(n_765), .Y(n_682) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_105), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_106), .Y(n_579) );
INVx1_ASAP7_75t_L g877 ( .A(n_108), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_108), .A2(n_120), .B1(n_495), .B2(n_603), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_109), .Y(n_1043) );
XNOR2xp5_ASAP7_75t_L g261 ( .A(n_110), .B(n_262), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_110), .A2(n_151), .B1(n_1158), .B2(n_1177), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_111), .Y(n_1031) );
INVx1_ASAP7_75t_L g498 ( .A(n_112), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_112), .A2(n_178), .B1(n_558), .B2(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g1002 ( .A(n_113), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_115), .Y(n_790) );
OAI221xp5_ASAP7_75t_L g807 ( .A1(n_115), .A2(n_305), .B1(n_318), .B2(n_355), .C(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g1035 ( .A(n_116), .Y(n_1035) );
INVx1_ASAP7_75t_L g1189 ( .A(n_117), .Y(n_1189) );
INVxp67_ASAP7_75t_SL g826 ( .A(n_118), .Y(n_826) );
INVx1_ASAP7_75t_L g890 ( .A(n_119), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g906 ( .A1(n_119), .A2(n_123), .B1(n_588), .B2(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g869 ( .A(n_120), .Y(n_869) );
INVx1_ASAP7_75t_L g973 ( .A(n_122), .Y(n_973) );
INVx1_ASAP7_75t_L g885 ( .A(n_123), .Y(n_885) );
INVx1_ASAP7_75t_L g471 ( .A(n_124), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_125), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_126), .A2(n_202), .B1(n_349), .B2(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g622 ( .A(n_126), .Y(n_622) );
INVx1_ASAP7_75t_L g655 ( .A(n_127), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_127), .A2(n_131), .B1(n_562), .B2(n_563), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_128), .A2(n_158), .B1(n_400), .B2(n_495), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_128), .A2(n_158), .B1(n_586), .B2(n_588), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_129), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_130), .A2(n_154), .B1(n_526), .B2(n_528), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_130), .A2(n_154), .B1(n_556), .B2(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g656 ( .A(n_131), .Y(n_656) );
INVx1_ASAP7_75t_L g435 ( .A(n_132), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_133), .A2(n_143), .B1(n_1171), .B2(n_1174), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_134), .A2(n_187), .B1(n_337), .B2(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g424 ( .A(n_134), .Y(n_424) );
INVx1_ASAP7_75t_L g618 ( .A(n_135), .Y(n_618) );
INVxp33_ASAP7_75t_SL g1090 ( .A(n_136), .Y(n_1090) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_136), .A2(n_175), .B1(n_1105), .B2(n_1112), .Y(n_1111) );
AOI22x1_ASAP7_75t_SL g628 ( .A1(n_137), .A2(n_629), .B1(n_676), .B2(n_677), .Y(n_628) );
INVx1_ASAP7_75t_L g676 ( .A(n_137), .Y(n_676) );
INVx1_ASAP7_75t_L g805 ( .A(n_139), .Y(n_805) );
INVx1_ASAP7_75t_L g1395 ( .A(n_140), .Y(n_1395) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_141), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g995 ( .A(n_142), .Y(n_995) );
INVx1_ASAP7_75t_L g633 ( .A(n_144), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_144), .A2(n_192), .B1(n_495), .B2(n_526), .Y(n_662) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_145), .Y(n_243) );
AND3x2_ASAP7_75t_L g1156 ( .A(n_145), .B(n_241), .C(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_145), .B(n_241), .Y(n_1163) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_147), .A2(n_182), .B1(n_1152), .B2(n_1195), .Y(n_1194) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_148), .Y(n_697) );
INVx2_ASAP7_75t_L g254 ( .A(n_149), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_150), .Y(n_872) );
INVx1_ASAP7_75t_L g1418 ( .A(n_152), .Y(n_1418) );
INVx1_ASAP7_75t_L g1392 ( .A(n_153), .Y(n_1392) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_155), .A2(n_162), .B1(n_1158), .B2(n_1177), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_157), .A2(n_179), .B1(n_1105), .B2(n_1107), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_157), .A2(n_179), .B1(n_1116), .B2(n_1118), .Y(n_1115) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_159), .Y(n_635) );
INVx1_ASAP7_75t_L g477 ( .A(n_160), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_160), .A2(n_188), .B1(n_503), .B2(n_505), .Y(n_502) );
INVx1_ASAP7_75t_L g1157 ( .A(n_161), .Y(n_1157) );
INVx1_ASAP7_75t_L g359 ( .A(n_163), .Y(n_359) );
INVx1_ASAP7_75t_L g578 ( .A(n_164), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g814 ( .A(n_165), .Y(n_814) );
INVx1_ASAP7_75t_L g1255 ( .A(n_166), .Y(n_1255) );
XOR2xp5_ASAP7_75t_L g1434 ( .A(n_167), .B(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g581 ( .A(n_168), .Y(n_581) );
INVx1_ASAP7_75t_L g945 ( .A(n_170), .Y(n_945) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_171), .A2(n_211), .B1(n_495), .B2(n_544), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_171), .A2(n_211), .B1(n_560), .B2(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g1024 ( .A(n_172), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g1067 ( .A1(n_172), .A2(n_226), .B1(n_1055), .B2(n_1068), .C(n_1070), .Y(n_1067) );
INVx1_ASAP7_75t_L g514 ( .A(n_173), .Y(n_514) );
INVx1_ASAP7_75t_L g954 ( .A(n_174), .Y(n_954) );
INVxp33_ASAP7_75t_L g1093 ( .A(n_175), .Y(n_1093) );
INVx1_ASAP7_75t_L g256 ( .A(n_176), .Y(n_256) );
INVx2_ASAP7_75t_L g380 ( .A(n_176), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_177), .A2(n_200), .B1(n_551), .B2(n_943), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_177), .A2(n_200), .B1(n_441), .B2(n_446), .Y(n_974) );
INVx1_ASAP7_75t_L g517 ( .A(n_178), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_180), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_181), .A2(n_206), .B1(n_1171), .B2(n_1174), .Y(n_1170) );
INVx1_ASAP7_75t_L g775 ( .A(n_183), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g799 ( .A1(n_183), .A2(n_203), .B1(n_588), .B2(n_800), .C(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g880 ( .A(n_184), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_185), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g986 ( .A(n_186), .B(n_987), .Y(n_986) );
XNOR2x1_ASAP7_75t_L g1140 ( .A(n_186), .B(n_987), .Y(n_1140) );
INVx1_ASAP7_75t_L g428 ( .A(n_187), .Y(n_428) );
INVx1_ASAP7_75t_L g483 ( .A(n_188), .Y(n_483) );
INVx1_ASAP7_75t_L g941 ( .A(n_190), .Y(n_941) );
OAI211xp5_ASAP7_75t_SL g947 ( .A1(n_190), .A2(n_375), .B(n_948), .C(n_957), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_193), .Y(n_782) );
INVx1_ASAP7_75t_L g736 ( .A(n_194), .Y(n_736) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_197), .A2(n_637), .B(n_706), .C(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g762 ( .A(n_197), .Y(n_762) );
INVx1_ASAP7_75t_L g789 ( .A(n_198), .Y(n_789) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_198), .Y(n_808) );
INVx1_ASAP7_75t_L g823 ( .A(n_199), .Y(n_823) );
INVx1_ASAP7_75t_L g884 ( .A(n_201), .Y(n_884) );
INVx1_ASAP7_75t_L g624 ( .A(n_202), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g777 ( .A1(n_203), .A2(n_370), .B(n_741), .Y(n_777) );
INVx1_ASAP7_75t_L g1217 ( .A(n_204), .Y(n_1217) );
INVx1_ASAP7_75t_L g1155 ( .A(n_205), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_205), .B(n_1165), .Y(n_1168) );
INVx1_ASAP7_75t_L g1096 ( .A(n_207), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_207), .A2(n_222), .B1(n_620), .B2(n_652), .Y(n_1131) );
OAI221xp5_ASAP7_75t_L g1408 ( .A1(n_208), .A2(n_416), .B1(n_438), .B2(n_1409), .C(n_1415), .Y(n_1408) );
INVx1_ASAP7_75t_L g1092 ( .A(n_209), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_210), .Y(n_267) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_212), .A2(n_419), .B(n_693), .C(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g733 ( .A(n_212), .Y(n_733) );
INVx1_ASAP7_75t_L g819 ( .A(n_213), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_214), .Y(n_931) );
INVx2_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_216), .Y(n_1033) );
OAI221xp5_ASAP7_75t_L g1004 ( .A1(n_217), .A2(n_220), .B1(n_1005), .B2(n_1012), .C(n_1014), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_217), .A2(n_220), .B1(n_1049), .B2(n_1052), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_218), .A2(n_219), .B1(n_338), .B2(n_343), .Y(n_342) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_218), .A2(n_375), .B(n_385), .C(n_408), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_219), .A2(n_416), .B1(n_418), .B2(n_432), .C(n_438), .Y(n_415) );
INVx1_ASAP7_75t_L g873 ( .A(n_221), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_221), .A2(n_223), .B1(n_596), .B2(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g1097 ( .A(n_222), .Y(n_1097) );
INVx1_ASAP7_75t_L g870 ( .A(n_223), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_224), .Y(n_721) );
INVx1_ASAP7_75t_L g1026 ( .A(n_226), .Y(n_1026) );
INVx1_ASAP7_75t_L g273 ( .A(n_227), .Y(n_273) );
BUFx3_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
BUFx3_ASAP7_75t_L g272 ( .A(n_228), .Y(n_272) );
INVx1_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
INVx1_ASAP7_75t_L g1028 ( .A(n_230), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_231), .Y(n_1389) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_232), .Y(n_711) );
XNOR2xp5_ASAP7_75t_L g916 ( .A(n_233), .B(n_917), .Y(n_916) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_257), .B(n_1144), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_244), .Y(n_238) );
AND2x4_ASAP7_75t_L g1427 ( .A(n_239), .B(n_245), .Y(n_1427) );
NOR2xp33_ASAP7_75t_SL g239 ( .A(n_240), .B(n_242), .Y(n_239) );
INVx1_ASAP7_75t_SL g1432 ( .A(n_240), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_240), .B(n_242), .Y(n_1442) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_242), .B(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x6_ASAP7_75t_L g520 ( .A(n_247), .B(n_351), .Y(n_520) );
OR2x2_ASAP7_75t_L g684 ( .A(n_247), .B(n_351), .Y(n_684) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g431 ( .A(n_248), .B(n_256), .Y(n_431) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g741 ( .A(n_249), .B(n_510), .Y(n_741) );
INVx8_ASAP7_75t_L g516 ( .A(n_250), .Y(n_516) );
OR2x6_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_251), .Y(n_427) );
OR2x6_ASAP7_75t_L g519 ( .A(n_251), .B(n_509), .Y(n_519) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_251), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1041 ( .A(n_251), .B(n_1011), .Y(n_1041) );
INVx1_ASAP7_75t_L g1413 ( .A(n_251), .Y(n_1413) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g372 ( .A(n_253), .B(n_254), .Y(n_372) );
INVx1_ASAP7_75t_L g383 ( .A(n_253), .Y(n_383) );
INVx2_ASAP7_75t_L g390 ( .A(n_253), .Y(n_390) );
AND2x4_ASAP7_75t_L g396 ( .A(n_253), .B(n_384), .Y(n_396) );
INVx1_ASAP7_75t_L g423 ( .A(n_253), .Y(n_423) );
INVx2_ASAP7_75t_L g384 ( .A(n_254), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_254), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g411 ( .A(n_254), .Y(n_411) );
INVx1_ASAP7_75t_L g422 ( .A(n_254), .Y(n_422) );
INVx1_ASAP7_75t_L g445 ( .A(n_254), .Y(n_445) );
AND2x4_ASAP7_75t_L g504 ( .A(n_255), .B(n_411), .Y(n_504) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g505 ( .A(n_256), .B(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g652 ( .A(n_256), .B(n_506), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_913), .B1(n_1142), .B2(n_1143), .Y(n_257) );
INVx1_ASAP7_75t_L g1142 ( .A(n_258), .Y(n_1142) );
AO22x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_678), .B1(n_679), .B2(n_912), .Y(n_258) );
INVx1_ASAP7_75t_L g912 ( .A(n_259), .Y(n_912) );
XOR2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_451), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND3xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_358), .C(n_373), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_301), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_286), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B1(n_278), .B2(n_279), .Y(n_266) );
OAI221xp5_ASAP7_75t_L g385 ( .A1(n_267), .A2(n_296), .B1(n_386), .B2(n_391), .C(n_397), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_268), .A2(n_279), .B1(n_780), .B2(n_782), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_268), .A2(n_279), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
CKINVDCx6p67_ASAP7_75t_R g268 ( .A(n_269), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
OR2x2_ASAP7_75t_L g977 ( .A(n_270), .B(n_274), .Y(n_977) );
INVx2_ASAP7_75t_L g1074 ( .A(n_270), .Y(n_1074) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g335 ( .A(n_271), .Y(n_335) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_271), .Y(n_473) );
INVx1_ASAP7_75t_L g564 ( .A(n_271), .Y(n_564) );
BUFx6f_ASAP7_75t_L g903 ( .A(n_271), .Y(n_903) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g294 ( .A(n_272), .Y(n_294) );
AND2x2_ASAP7_75t_L g341 ( .A(n_272), .B(n_293), .Y(n_341) );
INVx1_ASAP7_75t_L g283 ( .A(n_273), .Y(n_283) );
OR2x6_ASAP7_75t_L g280 ( .A(n_274), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
OR2x2_ASAP7_75t_L g979 ( .A(n_274), .B(n_980), .Y(n_979) );
OR2x2_ASAP7_75t_L g981 ( .A(n_274), .B(n_982), .Y(n_981) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx2_ASAP7_75t_L g1047 ( .A(n_275), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_275), .B(n_644), .Y(n_1079) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_275), .B(n_335), .Y(n_1081) );
INVx1_ASAP7_75t_L g312 ( .A(n_276), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_277), .Y(n_315) );
AND2x4_ASAP7_75t_L g994 ( .A(n_277), .B(n_379), .Y(n_994) );
CKINVDCx6p67_ASAP7_75t_R g279 ( .A(n_280), .Y(n_279) );
BUFx3_ASAP7_75t_L g732 ( .A(n_281), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_281), .A2(n_927), .B1(n_930), .B2(n_931), .C(n_932), .Y(n_926) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g730 ( .A(n_282), .Y(n_730) );
BUFx4f_ASAP7_75t_L g940 ( .A(n_282), .Y(n_940) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
OR2x2_ASAP7_75t_L g644 ( .A(n_283), .B(n_284), .Y(n_644) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g300 ( .A(n_285), .B(n_293), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B1(n_296), .B2(n_297), .Y(n_286) );
AOI222xp33_ASAP7_75t_L g809 ( .A1(n_288), .A2(n_297), .B1(n_361), .B2(n_779), .C1(n_786), .C2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_288), .A2(n_297), .B1(n_1392), .B2(n_1393), .Y(n_1391) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_295), .Y(n_288) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_289), .Y(n_1121) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g560 ( .A(n_290), .Y(n_560) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g337 ( .A(n_291), .Y(n_337) );
INVx6_ASAP7_75t_L g345 ( .A(n_291), .Y(n_345) );
AND2x2_ASAP7_75t_L g362 ( .A(n_291), .B(n_311), .Y(n_362) );
AND2x4_ASAP7_75t_L g468 ( .A(n_291), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
AND2x2_ASAP7_75t_L g297 ( .A(n_295), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g615 ( .A(n_299), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_299), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g331 ( .A(n_300), .Y(n_331) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
AND2x6_ASAP7_75t_L g463 ( .A(n_300), .B(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_300), .Y(n_552) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_300), .Y(n_667) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_300), .Y(n_709) );
BUFx2_ASAP7_75t_L g842 ( .A(n_300), .Y(n_842) );
BUFx3_ASAP7_75t_L g1117 ( .A(n_300), .Y(n_1117) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_322), .C(n_353), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_316), .B2(n_317), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_303), .A2(n_316), .B1(n_409), .B2(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g924 ( .A(n_304), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_304), .A2(n_317), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g1051 ( .A(n_307), .Y(n_1051) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g482 ( .A(n_308), .Y(n_482) );
INVx2_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
OR2x6_ASAP7_75t_L g318 ( .A(n_310), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_311), .B(n_315), .Y(n_310) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_311), .B(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1053 ( .A(n_311), .Y(n_1053) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x4_ASAP7_75t_L g352 ( .A(n_313), .B(n_327), .Y(n_352) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g326 ( .A(n_314), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g460 ( .A(n_314), .Y(n_460) );
INVx1_ASAP7_75t_L g465 ( .A(n_314), .Y(n_465) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_314), .Y(n_470) );
OR2x6_ASAP7_75t_L g547 ( .A(n_315), .B(n_405), .Y(n_547) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_319), .B(n_1053), .Y(n_1052) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x6_ASAP7_75t_L g484 ( .A(n_321), .B(n_465), .Y(n_484) );
AOI33xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_330), .A3(n_336), .B1(n_342), .B2(n_346), .B3(n_350), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_323), .A2(n_566), .B1(n_799), .B2(n_803), .C(n_807), .Y(n_798) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_324), .Y(n_549) );
OAI22xp5_ASAP7_75t_SL g925 ( .A1(n_324), .A2(n_926), .B1(n_933), .B2(n_935), .Y(n_925) );
OR2x6_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
OR2x2_ASAP7_75t_L g715 ( .A(n_325), .B(n_328), .Y(n_715) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g593 ( .A(n_326), .Y(n_593) );
INVx2_ASAP7_75t_SL g1070 ( .A(n_326), .Y(n_1070) );
INVx1_ASAP7_75t_L g491 ( .A(n_327), .Y(n_491) );
INVx2_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
BUFx2_ASAP7_75t_L g450 ( .A(n_328), .Y(n_450) );
AND2x4_ASAP7_75t_L g524 ( .A(n_328), .B(n_431), .Y(n_524) );
OR2x2_ASAP7_75t_L g592 ( .A(n_328), .B(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g658 ( .A(n_328), .B(n_431), .Y(n_658) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g492 ( .A(n_329), .Y(n_492) );
OR2x6_ASAP7_75t_L g740 ( .A(n_329), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g349 ( .A(n_333), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_333), .A2(n_720), .B1(n_805), .B2(n_806), .Y(n_804) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g723 ( .A(n_335), .Y(n_723) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g558 ( .A(n_339), .Y(n_558) );
INVx2_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_340), .Y(n_356) );
BUFx4f_ASAP7_75t_L g476 ( .A(n_340), .Y(n_476) );
BUFx3_ASAP7_75t_L g670 ( .A(n_340), .Y(n_670) );
INVx1_ASAP7_75t_L g847 ( .A(n_340), .Y(n_847) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_340), .B(n_1047), .Y(n_1066) );
INVx1_ASAP7_75t_L g1069 ( .A(n_340), .Y(n_1069) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_341), .Y(n_488) );
INVx4_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g613 ( .A(n_344), .Y(n_613) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g461 ( .A(n_345), .Y(n_461) );
INVx2_ASAP7_75t_L g557 ( .A(n_345), .Y(n_557) );
INVx2_ASAP7_75t_L g587 ( .A(n_345), .Y(n_587) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_345), .Y(n_801) );
INVx1_ASAP7_75t_L g907 ( .A(n_345), .Y(n_907) );
BUFx4f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g562 ( .A(n_348), .Y(n_562) );
INVx1_ASAP7_75t_L g982 ( .A(n_348), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_350), .B(n_612), .C(n_614), .Y(n_611) );
AOI33xp33_ASAP7_75t_L g839 ( .A1(n_350), .A2(n_840), .A3(n_841), .B1(n_844), .B2(n_845), .B3(n_848), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g905 ( .A(n_350), .B(n_906), .C(n_908), .Y(n_905) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x4_ASAP7_75t_L g361 ( .A(n_351), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g566 ( .A(n_351), .B(n_352), .Y(n_566) );
INVx2_ASAP7_75t_L g1062 ( .A(n_352), .Y(n_1062) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND3xp33_ASAP7_75t_SL g1378 ( .A(n_355), .B(n_1379), .C(n_1382), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g1125 ( .A(n_356), .Y(n_1125) );
AND2x2_ASAP7_75t_L g920 ( .A(n_357), .B(n_921), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_360), .B(n_945), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_360), .B(n_1395), .Y(n_1394) );
OR2x6_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx2_ASAP7_75t_L g1042 ( .A(n_361), .Y(n_1042) );
NOR2xp67_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx2_ASAP7_75t_L g797 ( .A(n_364), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_370), .Y(n_365) );
AND2x2_ASAP7_75t_L g409 ( .A(n_366), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g959 ( .A(n_366), .B(n_410), .Y(n_959) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x6_ASAP7_75t_L g413 ( .A(n_367), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g438 ( .A(n_367), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g792 ( .A(n_367), .Y(n_792) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g603 ( .A(n_370), .Y(n_603) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g527 ( .A(n_371), .Y(n_527) );
INVx2_ASAP7_75t_SL g1001 ( .A(n_371), .Y(n_1001) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
OAI31xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_415), .A3(n_440), .B(n_448), .Y(n_373) );
INVx8_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
AND2x4_ASAP7_75t_L g447 ( .A(n_377), .B(n_394), .Y(n_447) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g417 ( .A(n_379), .B(n_402), .Y(n_417) );
AND2x2_ASAP7_75t_L g442 ( .A(n_379), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g406 ( .A(n_380), .Y(n_406) );
INVx1_ASAP7_75t_L g510 ( .A(n_380), .Y(n_510) );
INVx1_ASAP7_75t_L g399 ( .A(n_381), .Y(n_399) );
BUFx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_382), .Y(n_497) );
AND2x4_ASAP7_75t_L g499 ( .A(n_382), .B(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_382), .Y(n_530) );
BUFx2_ASAP7_75t_L g888 ( .A(n_382), .Y(n_888) );
BUFx3_ASAP7_75t_L g997 ( .A(n_382), .Y(n_997) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g434 ( .A(n_388), .Y(n_434) );
INVx1_ASAP7_75t_L g968 ( .A(n_388), .Y(n_968) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g690 ( .A(n_389), .Y(n_690) );
INVx1_ASAP7_75t_L g751 ( .A(n_389), .Y(n_751) );
INVx1_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
AND2x4_ASAP7_75t_L g443 ( .A(n_390), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g608 ( .A(n_393), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_393), .A2(n_717), .B1(n_721), .B2(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g1403 ( .A(n_395), .Y(n_1403) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g437 ( .A(n_396), .Y(n_437) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_396), .Y(n_535) );
INVx3_ASAP7_75t_L g601 ( .A(n_396), .Y(n_601) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g1130 ( .A(n_399), .Y(n_1130) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g695 ( .A(n_401), .Y(n_695) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_402), .Y(n_544) );
INVx2_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g956 ( .A(n_404), .Y(n_956) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g784 ( .A(n_405), .Y(n_784) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g501 ( .A(n_406), .Y(n_501) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_411), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g1009 ( .A(n_411), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_412), .A2(n_958), .B1(n_959), .B2(n_960), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_412), .A2(n_959), .B1(n_1380), .B2(n_1381), .Y(n_1407) );
CKINVDCx11_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g791 ( .A(n_414), .Y(n_791) );
CKINVDCx6p67_ASAP7_75t_R g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_424), .B1(n_425), .B2(n_428), .C(n_429), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g962 ( .A1(n_419), .A2(n_930), .B1(n_931), .B2(n_963), .C(n_964), .Y(n_962) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g439 ( .A(n_421), .Y(n_439) );
INVx2_ASAP7_75t_L g651 ( .A(n_421), .Y(n_651) );
INVx3_ASAP7_75t_L g776 ( .A(n_421), .Y(n_776) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_422), .B(n_423), .Y(n_761) );
INVx1_ASAP7_75t_L g506 ( .A(n_423), .Y(n_506) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_427), .A2(n_725), .B1(n_728), .B2(n_743), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_427), .A2(n_757), .B1(n_758), .B2(n_762), .Y(n_756) );
BUFx2_ASAP7_75t_L g963 ( .A(n_427), .Y(n_963) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_SL g964 ( .A(n_431), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_435), .B2(n_436), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_434), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_434), .A2(n_599), .B1(n_779), .B2(n_780), .Y(n_778) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g513 ( .A(n_437), .Y(n_513) );
INVx1_ASAP7_75t_L g744 ( .A(n_439), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_439), .B(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g794 ( .A(n_442), .Y(n_794) );
AND2x4_ASAP7_75t_L g508 ( .A(n_443), .B(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g532 ( .A(n_443), .Y(n_532) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_443), .Y(n_539) );
INVx1_ASAP7_75t_L g597 ( .A(n_443), .Y(n_597) );
BUFx2_ASAP7_75t_L g607 ( .A(n_443), .Y(n_607) );
BUFx6f_ASAP7_75t_L g1106 ( .A(n_443), .Y(n_1106) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g795 ( .A(n_447), .Y(n_795) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
CKINVDCx8_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
OAI31xp33_ASAP7_75t_L g946 ( .A1(n_450), .A2(n_947), .A3(n_961), .B(n_974), .Y(n_946) );
XNOR2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_567), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI211x1_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_489), .B(n_493), .C(n_521), .Y(n_454) );
NAND4xp25_ASAP7_75t_SL g455 ( .A(n_456), .B(n_466), .C(n_474), .D(n_485), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_462), .B2(n_463), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_458), .A2(n_468), .B1(n_578), .B2(n_579), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_458), .A2(n_472), .B1(n_869), .B2(n_870), .Y(n_868) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
AND2x6_ASAP7_75t_L g472 ( .A(n_459), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g859 ( .A(n_459), .B(n_461), .Y(n_859) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g855 ( .A(n_460), .B(n_856), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_463), .A2(n_472), .B1(n_581), .B2(n_582), .Y(n_580) );
CKINVDCx6p67_ASAP7_75t_R g639 ( .A(n_463), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_463), .A2(n_472), .B1(n_861), .B2(n_862), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_463), .A2(n_468), .B1(n_872), .B2(n_873), .C(n_874), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_463), .A2(n_859), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
INVx1_ASAP7_75t_L g487 ( .A(n_464), .Y(n_487) );
INVx1_ASAP7_75t_L g643 ( .A(n_464), .Y(n_643) );
AND2x2_ASAP7_75t_L g707 ( .A(n_464), .B(n_574), .Y(n_707) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_471), .B2(n_472), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_467), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_515) );
INVx4_ASAP7_75t_L g645 ( .A(n_468), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_468), .A2(n_823), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_468), .A2(n_472), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
AND2x4_ASAP7_75t_L g480 ( .A(n_469), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_SL g712 ( .A(n_469), .B(n_481), .Y(n_712) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx4_ASAP7_75t_L g640 ( .A(n_472), .Y(n_640) );
INVx2_ASAP7_75t_L g554 ( .A(n_473), .Y(n_554) );
INVx1_ASAP7_75t_L g737 ( .A(n_473), .Y(n_737) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_473), .Y(n_843) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_473), .Y(n_849) );
INVx1_ASAP7_75t_L g1119 ( .A(n_473), .Y(n_1119) );
AOI222xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_477), .B2(n_478), .C1(n_483), .C2(n_484), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_480), .A2(n_484), .B1(n_635), .B2(n_636), .Y(n_634) );
AOI222xp33_ASAP7_75t_L g1094 ( .A1(n_480), .A2(n_484), .B1(n_670), .B2(n_1095), .C1(n_1096), .C2(n_1097), .Y(n_1094) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g856 ( .A(n_482), .Y(n_856) );
INVx3_ASAP7_75t_L g576 ( .A(n_484), .Y(n_576) );
AOI322xp5_ASAP7_75t_L g708 ( .A1(n_484), .A2(n_697), .A3(n_701), .B1(n_709), .B2(n_710), .C1(n_711), .C2(n_712), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g1087 ( .A(n_485), .B(n_1088), .C(n_1091), .D(n_1094), .Y(n_1087) );
INVx5_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_486), .A2(n_572), .B(n_573), .C(n_575), .Y(n_571) );
CKINVDCx8_ASAP7_75t_R g637 ( .A(n_486), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g851 ( .A1(n_486), .A2(n_707), .B(n_852), .C(n_853), .Y(n_851) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g876 ( .A1(n_487), .A2(n_674), .B(n_877), .Y(n_876) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_488), .Y(n_574) );
INVx2_ASAP7_75t_L g589 ( .A(n_488), .Y(n_589) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_488), .Y(n_674) );
INVx1_ASAP7_75t_L g922 ( .A(n_488), .Y(n_922) );
AOI221x1_ASAP7_75t_L g866 ( .A1(n_489), .A2(n_816), .B1(n_867), .B2(n_878), .C(n_891), .Y(n_866) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AO211x2_ASAP7_75t_L g569 ( .A1(n_490), .A2(n_570), .B(n_583), .C(n_616), .Y(n_569) );
INVx1_ASAP7_75t_L g1099 ( .A(n_490), .Y(n_1099) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_L g646 ( .A(n_491), .B(n_492), .Y(n_646) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_492), .Y(n_1083) );
INVx2_ASAP7_75t_L g1422 ( .A(n_492), .Y(n_1422) );
AOI31xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_507), .A3(n_515), .B(n_520), .Y(n_493) );
AOI211xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B(n_499), .C(n_502), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_497), .Y(n_610) );
BUFx2_ASAP7_75t_L g838 ( .A(n_497), .Y(n_838) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_499), .A2(n_528), .B(n_618), .C(n_619), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_499), .B(n_649), .C(n_653), .Y(n_648) );
CKINVDCx11_ASAP7_75t_R g693 ( .A(n_499), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g1128 ( .A1(n_499), .A2(n_1129), .B(n_1130), .C(n_1131), .Y(n_1128) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_L g700 ( .A(n_501), .Y(n_700) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g620 ( .A(n_504), .Y(n_620) );
INVx2_ASAP7_75t_L g650 ( .A(n_504), .Y(n_650) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_504), .A2(n_689), .A3(n_695), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_701), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g882 ( .A1(n_504), .A2(n_698), .B1(n_883), .B2(n_884), .C1(n_885), .C2(n_886), .Y(n_882) );
INVx1_ASAP7_75t_L g699 ( .A(n_506), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .B1(n_512), .B2(n_514), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_508), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_508), .A2(n_623), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_508), .A2(n_512), .B1(n_819), .B2(n_820), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_508), .A2(n_512), .B1(n_880), .B2(n_881), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g1132 ( .A1(n_508), .A2(n_512), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
AND2x4_ASAP7_75t_L g512 ( .A(n_509), .B(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g623 ( .A(n_509), .B(n_513), .Y(n_623) );
INVx1_ASAP7_75t_L g689 ( .A(n_509), .Y(n_689) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_516), .A2(n_579), .B1(n_626), .B2(n_627), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_516), .A2(n_686), .B(n_687), .C(n_692), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_516), .A2(n_518), .B1(n_822), .B2(n_823), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_516), .A2(n_518), .B1(n_872), .B2(n_890), .Y(n_889) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_516), .A2(n_627), .B1(n_1092), .B2(n_1136), .Y(n_1135) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g627 ( .A(n_519), .Y(n_627) );
AOI31xp33_ASAP7_75t_L g616 ( .A1(n_520), .A2(n_617), .A3(n_621), .B(n_625), .Y(n_616) );
AO21x1_ASAP7_75t_SL g647 ( .A1(n_520), .A2(n_648), .B(n_654), .Y(n_647) );
CKINVDCx16_ASAP7_75t_R g816 ( .A(n_520), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_548), .Y(n_521) );
AOI33xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_525), .A3(n_531), .B1(n_536), .B2(n_541), .B3(n_546), .Y(n_522) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_524), .B(n_606), .C(n_609), .Y(n_605) );
INVx2_ASAP7_75t_L g1103 ( .A(n_524), .Y(n_1103) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g545 ( .A(n_529), .Y(n_545) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_530), .Y(n_832) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g540 ( .A(n_535), .Y(n_540) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_535), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_535), .Y(n_1032) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_539), .B(n_994), .Y(n_1003) );
INVx1_ASAP7_75t_L g1419 ( .A(n_540), .Y(n_1419) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_544), .A2(n_786), .B(n_787), .C(n_792), .Y(n_785) );
AOI222xp33_ASAP7_75t_L g824 ( .A1(n_545), .A2(n_698), .B1(n_825), .B2(n_826), .C1(n_827), .C2(n_828), .Y(n_824) );
AOI33xp33_ASAP7_75t_L g657 ( .A1(n_546), .A2(n_658), .A3(n_659), .B1(n_660), .B2(n_661), .B3(n_662), .Y(n_657) );
INVx2_ASAP7_75t_L g763 ( .A(n_546), .Y(n_763) );
AOI33xp33_ASAP7_75t_L g830 ( .A1(n_546), .A2(n_658), .A3(n_831), .B1(n_833), .B2(n_835), .B3(n_837), .Y(n_830) );
INVx6_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx5_ASAP7_75t_L g604 ( .A(n_547), .Y(n_604) );
AOI33xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .A3(n_555), .B1(n_559), .B2(n_561), .B3(n_565), .Y(n_548) );
AOI33xp33_ASAP7_75t_L g663 ( .A1(n_549), .A2(n_566), .A3(n_664), .B1(n_669), .B2(n_671), .B3(n_675), .Y(n_663) );
AOI33xp33_ASAP7_75t_L g1114 ( .A1(n_549), .A2(n_566), .A3(n_1115), .B1(n_1120), .B2(n_1123), .B3(n_1126), .Y(n_1114) );
AOI33xp33_ASAP7_75t_L g1382 ( .A1(n_549), .A2(n_565), .A3(n_1383), .B1(n_1384), .B2(n_1385), .B3(n_1386), .Y(n_1382) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g943 ( .A(n_554), .Y(n_943) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_557), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_558), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g668 ( .A(n_564), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_564), .A2(n_666), .B1(n_771), .B2(n_773), .Y(n_802) );
BUFx4f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx4_ASAP7_75t_L g738 ( .A(n_566), .Y(n_738) );
BUFx4f_ASAP7_75t_L g934 ( .A(n_566), .Y(n_934) );
XNOR2x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_628), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_577), .C(n_580), .Y(n_570) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_574), .Y(n_1122) );
NAND4xp25_ASAP7_75t_L g583 ( .A(n_584), .B(n_594), .C(n_605), .D(n_611), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .C(n_591), .Y(n_584) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g1073 ( .A(n_587), .Y(n_1073) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_591), .B(n_901), .C(n_904), .Y(n_900) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_602), .C(n_604), .Y(n_594) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g834 ( .A(n_599), .Y(n_834) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g772 ( .A(n_600), .Y(n_772) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g754 ( .A(n_601), .Y(n_754) );
INVx3_ASAP7_75t_L g972 ( .A(n_601), .Y(n_972) );
NAND3xp33_ASAP7_75t_L g896 ( .A(n_604), .B(n_897), .C(n_899), .Y(n_896) );
AOI33xp33_ASAP7_75t_L g1101 ( .A1(n_604), .A2(n_1102), .A3(n_1104), .B1(n_1109), .B2(n_1111), .B3(n_1113), .Y(n_1101) );
INVx1_ASAP7_75t_L g953 ( .A(n_608), .Y(n_953) );
INVx1_ASAP7_75t_L g827 ( .A(n_620), .Y(n_827) );
INVx5_ASAP7_75t_SL g691 ( .A(n_623), .Y(n_691) );
AND4x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_647), .C(n_657), .D(n_663), .Y(n_629) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_630), .B(n_647), .C(n_657), .D(n_663), .Y(n_677) );
OAI31xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_638), .A3(n_641), .B(n_646), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .C(n_637), .Y(n_631) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g710 ( .A(n_643), .Y(n_710) );
INVx2_ASAP7_75t_L g727 ( .A(n_644), .Y(n_727) );
INVx1_ASAP7_75t_L g929 ( .A(n_644), .Y(n_929) );
BUFx2_ASAP7_75t_L g1060 ( .A(n_644), .Y(n_1060) );
OAI31xp33_ASAP7_75t_SL g702 ( .A1(n_646), .A2(n_703), .A3(n_704), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_SL g863 ( .A(n_646), .Y(n_863) );
OAI21xp33_ASAP7_75t_L g781 ( .A1(n_651), .A2(n_782), .B(n_783), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_658), .B(n_893), .C(n_895), .Y(n_892) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g1046 ( .A(n_667), .B(n_1047), .Y(n_1046) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_667), .Y(n_1055) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_674), .B(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
XNOR2x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_812), .Y(n_680) );
XNOR2x1_ASAP7_75t_L g681 ( .A(n_682), .B(n_766), .Y(n_681) );
INVx1_ASAP7_75t_L g764 ( .A(n_683), .Y(n_764) );
OAI211xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B(n_702), .C(n_713), .Y(n_683) );
AOI31xp33_ASAP7_75t_L g1127 ( .A1(n_684), .A2(n_1128), .A3(n_1132), .B(n_1135), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_686), .A2(n_726), .B1(n_732), .B2(n_733), .Y(n_731) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx2_ASAP7_75t_L g747 ( .A(n_690), .Y(n_747) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_690), .Y(n_1027) );
NAND4xp25_ASAP7_75t_SL g817 ( .A(n_693), .B(n_818), .C(n_821), .D(n_824), .Y(n_817) );
NAND4xp25_ASAP7_75t_SL g878 ( .A(n_693), .B(n_879), .C(n_882), .D(n_889), .Y(n_878) );
AND2x4_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g720 ( .A(n_709), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_711), .A2(n_749), .B1(n_752), .B2(n_755), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_739), .Y(n_713) );
OAI33xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .A3(n_724), .B1(n_731), .B2(n_734), .B3(n_738), .Y(n_714) );
INVx1_ASAP7_75t_SL g840 ( .A(n_715), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_721), .B2(n_722), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI22xp33_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_726), .B1(n_728), .B2(n_729), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g936 ( .A(n_727), .Y(n_936) );
INVx1_ASAP7_75t_L g980 ( .A(n_727), .Y(n_980) );
BUFx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI33xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_742), .A3(n_745), .B1(n_748), .B2(n_756), .B3(n_763), .Y(n_739) );
OAI33xp33_ASAP7_75t_L g1016 ( .A1(n_740), .A2(n_763), .A3(n_1017), .B1(n_1025), .B2(n_1030), .B3(n_1034), .Y(n_1016) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g1417 ( .A(n_750), .Y(n_1417) );
BUFx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g951 ( .A(n_751), .Y(n_951) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g898 ( .A(n_754), .Y(n_898) );
INVx2_ASAP7_75t_L g1108 ( .A(n_754), .Y(n_1108) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND4xp25_ASAP7_75t_L g767 ( .A(n_768), .B(n_798), .C(n_809), .D(n_811), .Y(n_767) );
OAI31xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_793), .A3(n_796), .B(n_797), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_774), .B1(n_778), .B2(n_781), .C(n_785), .Y(n_769) );
INVx2_ASAP7_75t_L g836 ( .A(n_772), .Y(n_836) );
INVx2_ASAP7_75t_SL g894 ( .A(n_772), .Y(n_894) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g1023 ( .A(n_776), .Y(n_1023) );
BUFx2_ASAP7_75t_L g1410 ( .A(n_776), .Y(n_1410) );
NAND2x1p5_ASAP7_75t_L g1013 ( .A(n_791), .B(n_1010), .Y(n_1013) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OA22x2_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_864), .B1(n_865), .B2(n_911), .Y(n_812) );
INVx1_ASAP7_75t_L g911 ( .A(n_813), .Y(n_911) );
XNOR2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_814), .A2(n_1200), .B1(n_1201), .B2(n_1202), .Y(n_1199) );
AOI211xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B(n_829), .C(n_850), .Y(n_815) );
NAND2xp5_ASAP7_75t_SL g829 ( .A(n_830), .B(n_839), .Y(n_829) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
AOI31xp33_ASAP7_75t_SL g850 ( .A1(n_851), .A2(n_857), .A3(n_860), .B(n_863), .Y(n_850) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g875 ( .A(n_855), .Y(n_875) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g910 ( .A(n_866), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_871), .Y(n_867) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND4xp25_ASAP7_75t_L g891 ( .A(n_892), .B(n_896), .C(n_900), .D(n_905), .Y(n_891) );
BUFx6f_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g1057 ( .A(n_903), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g1143 ( .A(n_913), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_983), .B1(n_984), .B2(n_1141), .Y(n_913) );
INVx1_ASAP7_75t_L g1141 ( .A(n_914), .Y(n_1141) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
AND4x1_ASAP7_75t_L g917 ( .A(n_918), .B(n_944), .C(n_946), .D(n_975), .Y(n_917) );
NOR3xp33_ASAP7_75t_SL g918 ( .A(n_919), .B(n_923), .C(n_925), .Y(n_918) );
BUFx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
BUFx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g933 ( .A(n_934), .Y(n_933) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_941), .C(n_942), .Y(n_935) );
BUFx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g1059 ( .A(n_940), .Y(n_1059) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_952), .B1(n_953), .B2(n_954), .C(n_955), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
BUFx2_ASAP7_75t_L g1399 ( .A(n_951), .Y(n_1399) );
OAI221xp5_ASAP7_75t_L g1409 ( .A1(n_964), .A2(n_1410), .B1(n_1411), .B2(n_1412), .C(n_1414), .Y(n_1409) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_969), .B1(n_970), .B2(n_973), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_971), .Y(n_970) );
BUFx3_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
AND2x4_ASAP7_75t_L g993 ( .A(n_972), .B(n_994), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g975 ( .A(n_976), .B(n_978), .Y(n_975) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVxp67_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
AOI22x1_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_1084), .B1(n_1138), .B2(n_1139), .Y(n_985) );
AND2x2_ASAP7_75t_L g987 ( .A(n_988), .B(n_1038), .Y(n_987) );
NOR3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_1004), .C(n_1016), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_998), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .B1(n_995), .B2(n_996), .Y(n_990) );
BUFx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AND2x6_ASAP7_75t_L g996 ( .A(n_994), .B(n_997), .Y(n_996) );
AND2x4_ASAP7_75t_L g1000 ( .A(n_994), .B(n_1001), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g1058 ( .A1(n_995), .A2(n_999), .B1(n_1059), .B2(n_1060), .C(n_1061), .Y(n_1058) );
NAND2x1p5_ASAP7_75t_L g1015 ( .A(n_997), .B(n_1010), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1000), .B1(n_1002), .B2(n_1003), .Y(n_998) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_1001), .Y(n_1110) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1001), .Y(n_1406) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
NAND2x1_ASAP7_75t_SL g1007 ( .A(n_1008), .B(n_1010), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx3_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
BUFx4f_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
OAI22xp33_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1021), .B1(n_1022), .B2(n_1024), .Y(n_1017) );
OAI22xp33_ASAP7_75t_L g1034 ( .A1(n_1018), .A2(n_1035), .B1(n_1036), .B2(n_1037), .Y(n_1034) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1023), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1027), .B1(n_1028), .B2(n_1029), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_1027), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1030) );
AOI211xp5_ASAP7_75t_L g1045 ( .A1(n_1031), .A2(n_1046), .B(n_1048), .C(n_1054), .Y(n_1045) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1032), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_1033), .A2(n_1035), .B1(n_1078), .B2(n_1080), .Y(n_1077) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_1037), .A2(n_1064), .B1(n_1067), .B2(n_1071), .C(n_1075), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1043), .B(n_1044), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
AND2x4_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
AOI31xp33_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1063), .A3(n_1077), .B(n_1082), .Y(n_1044) );
INVx2_ASAP7_75t_SL g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_SL g1076 ( .A(n_1053), .Y(n_1076) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx6_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx4_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1084), .Y(n_1138) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1086), .Y(n_1137) );
AOI211x1_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1098), .B(n_1100), .C(n_1127), .Y(n_1086) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1114), .Y(n_1100) );
INVx2_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
BUFx3_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx3_ASAP7_75t_SL g1139 ( .A(n_1140), .Y(n_1139) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1370), .B1(n_1372), .B2(n_1423), .C(n_1428), .Y(n_1144) );
NOR2x1_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1307), .Y(n_1145) );
NAND3xp33_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1244), .C(n_1268), .Y(n_1146) );
AOI211xp5_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1178), .B(n_1206), .C(n_1236), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1148), .B(n_1227), .Y(n_1310) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_1149), .A2(n_1169), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1169), .Y(n_1149) );
INVx2_ASAP7_75t_SL g1232 ( .A(n_1150), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1150), .B(n_1192), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1150), .B(n_1169), .Y(n_1316) );
INVx2_ASAP7_75t_SL g1150 ( .A(n_1151), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1211 ( .A(n_1151), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1151), .B(n_1169), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1151), .B(n_1169), .Y(n_1289) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1152), .Y(n_1222) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1152), .Y(n_1254) );
BUFx3_ASAP7_75t_L g1371 ( .A(n_1152), .Y(n_1371) );
AND2x4_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1156), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1153), .B(n_1156), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g1441 ( .A(n_1153), .Y(n_1441) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_1154), .B(n_1156), .Y(n_1158) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1155), .B(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1157), .Y(n_1165) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1158), .Y(n_1196) );
INVx1_ASAP7_75t_SL g1201 ( .A(n_1158), .Y(n_1201) );
OAI22xp33_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B1(n_1166), .B2(n_1167), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_1161), .A2(n_1167), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
OAI22xp33_ASAP7_75t_L g1215 ( .A1(n_1161), .A2(n_1216), .B1(n_1217), .B2(n_1218), .Y(n_1215) );
BUFx3_ASAP7_75t_L g1258 ( .A(n_1161), .Y(n_1258) );
BUFx6f_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1162), .A2(n_1167), .B1(n_1188), .B2(n_1189), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1164), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_1163), .B(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1163), .Y(n_1173) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1164), .Y(n_1172) );
HB1xp67_ASAP7_75t_L g1440 ( .A(n_1165), .Y(n_1440) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1167), .Y(n_1219) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1168), .Y(n_1175) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1169), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1169), .B(n_1213), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1169), .B(n_1213), .Y(n_1265) );
OAI21xp33_ASAP7_75t_L g1269 ( .A1(n_1169), .A2(n_1270), .B(n_1272), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1169), .B(n_1214), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1176), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1173), .Y(n_1171) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1173), .B(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1177), .Y(n_1200) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1190), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1180), .B(n_1291), .Y(n_1290) );
NOR2xp33_ASAP7_75t_L g1301 ( .A(n_1180), .B(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1181), .B(n_1197), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1181), .B(n_1198), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1185), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1182), .B(n_1186), .Y(n_1209) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1182), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1182), .B(n_1198), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1182), .B(n_1186), .Y(n_1329) );
NOR2xp33_ASAP7_75t_SL g1359 ( .A(n_1182), .B(n_1360), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1184), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1185), .B(n_1197), .Y(n_1229) );
NOR3xp33_ASAP7_75t_L g1249 ( .A(n_1185), .B(n_1227), .C(n_1250), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1185), .B(n_1197), .Y(n_1280) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1186), .B(n_1197), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1186), .B(n_1242), .Y(n_1241) );
OAI322xp33_ASAP7_75t_L g1313 ( .A1(n_1186), .A2(n_1314), .A3(n_1317), .B1(n_1318), .B2(n_1320), .C1(n_1322), .C2(n_1324), .Y(n_1313) );
NOR2xp33_ASAP7_75t_L g1323 ( .A(n_1186), .B(n_1197), .Y(n_1323) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1197), .Y(n_1191) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1192), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1192), .B(n_1197), .Y(n_1243) );
INVx4_ASAP7_75t_L g1248 ( .A(n_1192), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_1192), .B(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1192), .B(n_1316), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1192), .B(n_1319), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1192), .B(n_1214), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1192), .B(n_1232), .Y(n_1360) );
AND2x6_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1194), .Y(n_1192) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_1196), .A2(n_1253), .B1(n_1254), .B2(n_1255), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1197), .B(n_1209), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1197), .B(n_1247), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1197), .B(n_1241), .Y(n_1303) );
CKINVDCx6p67_ASAP7_75t_R g1197 ( .A(n_1198), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1198), .B(n_1247), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1198), .B(n_1241), .Y(n_1283) );
AOI32xp33_ASAP7_75t_L g1285 ( .A1(n_1198), .A2(n_1264), .A3(n_1286), .B1(n_1290), .B2(n_1292), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1198), .B(n_1209), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1198), .B(n_1329), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1198), .B(n_1358), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1198), .B(n_1364), .Y(n_1363) );
OR2x6_ASAP7_75t_SL g1198 ( .A(n_1199), .B(n_1203), .Y(n_1198) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_1201), .A2(n_1221), .B1(n_1222), .B2(n_1223), .Y(n_1220) );
OAI221xp5_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1210), .B1(n_1225), .B2(n_1230), .C(n_1233), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1209), .B(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1209), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1212), .Y(n_1210) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1211), .Y(n_1342) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1211), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1212), .B(n_1234), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1224), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1213), .B(n_1232), .Y(n_1231) );
INVx3_ASAP7_75t_L g1277 ( .A(n_1213), .Y(n_1277) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1213), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1213), .B(n_1261), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1213), .B(n_1251), .Y(n_1317) );
INVx3_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1214), .B(n_1289), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1220), .Y(n_1214) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_1218), .Y(n_1260) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
NOR2x1_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1229), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1227), .B(n_1283), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1334 ( .A(n_1227), .B(n_1335), .Y(n_1334) );
NOR2x1_ASAP7_75t_R g1350 ( .A(n_1227), .B(n_1291), .Y(n_1350) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1228), .B(n_1235), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1228), .B(n_1279), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1228), .B(n_1295), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1368 ( .A(n_1228), .B(n_1283), .Y(n_1368) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1229), .Y(n_1297) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
AOI322xp5_ASAP7_75t_L g1296 ( .A1(n_1231), .A2(n_1277), .A3(n_1297), .B1(n_1298), .B2(n_1300), .C1(n_1301), .C2(n_1303), .Y(n_1296) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1232), .Y(n_1238) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1232), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1232), .B(n_1300), .Y(n_1321) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1232), .Y(n_1337) );
NOR2xp33_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1240), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1239), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1243), .Y(n_1240) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1241), .Y(n_1291) );
AOI211xp5_ASAP7_75t_L g1345 ( .A1(n_1242), .A2(n_1346), .B(n_1347), .C(n_1350), .Y(n_1345) );
O2A1O1Ixp33_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1249), .B(n_1261), .C(n_1262), .Y(n_1244) );
INVxp67_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1248), .B(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1248), .Y(n_1274) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_1248), .B(n_1329), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1248), .B(n_1288), .Y(n_1366) );
OAI31xp33_ASAP7_75t_L g1268 ( .A1(n_1250), .A2(n_1269), .A3(n_1281), .B(n_1284), .Y(n_1268) );
OAI221xp5_ASAP7_75t_L g1355 ( .A1(n_1250), .A2(n_1289), .B1(n_1356), .B2(n_1361), .C(n_1365), .Y(n_1355) );
CKINVDCx5p33_ASAP7_75t_R g1250 ( .A(n_1251), .Y(n_1250) );
AOI22xp5_ASAP7_75t_L g1330 ( .A1(n_1251), .A2(n_1331), .B1(n_1340), .B2(n_1341), .Y(n_1330) );
OR2x6_ASAP7_75t_SL g1251 ( .A(n_1252), .B(n_1256), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1258), .B1(n_1259), .B2(n_1260), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1261), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1266), .Y(n_1263) );
AOI322xp5_ASAP7_75t_L g1356 ( .A1(n_1264), .A2(n_1277), .A3(n_1280), .B1(n_1315), .B2(n_1316), .C1(n_1357), .C2(n_1359), .Y(n_1356) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1266), .B(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1267), .Y(n_1293) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
OAI21xp5_ASAP7_75t_SL g1272 ( .A1(n_1273), .A2(n_1275), .B(n_1280), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1274), .B(n_1295), .Y(n_1294) );
NOR2xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1278), .Y(n_1275) );
INVx1_ASAP7_75t_SL g1276 ( .A(n_1277), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1277), .B(n_1282), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1277), .B(n_1303), .Y(n_1339) );
AOI21xp5_ASAP7_75t_L g1338 ( .A1(n_1278), .A2(n_1291), .B(n_1332), .Y(n_1338) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1278), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1280), .B(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1283), .Y(n_1312) );
NAND3xp33_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1296), .C(n_1304), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1288), .B(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1294), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1293), .B(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1295), .Y(n_1332) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
A2O1A1Ixp33_ASAP7_75t_L g1352 ( .A1(n_1299), .A2(n_1312), .B(n_1328), .C(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1300), .Y(n_1335) );
AOI211xp5_ASAP7_75t_SL g1351 ( .A1(n_1300), .A2(n_1352), .B(n_1355), .C(n_1367), .Y(n_1351) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1302), .Y(n_1354) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1303), .B(n_1323), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1303), .B(n_1337), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1303), .B(n_1354), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1306), .Y(n_1304) );
AOI211xp5_ASAP7_75t_L g1333 ( .A1(n_1305), .A2(n_1334), .B(n_1336), .C(n_1338), .Y(n_1333) );
NAND3xp33_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1330), .C(n_1351), .Y(n_1307) );
AOI211xp5_ASAP7_75t_SL g1308 ( .A1(n_1309), .A2(n_1311), .B(n_1313), .C(n_1326), .Y(n_1308) );
INVxp67_ASAP7_75t_SL g1309 ( .A(n_1310), .Y(n_1309) );
OAI211xp5_ASAP7_75t_L g1341 ( .A1(n_1312), .A2(n_1342), .B(n_1343), .C(n_1345), .Y(n_1341) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1317), .Y(n_1340) );
OAI211xp5_ASAP7_75t_L g1331 ( .A1(n_1320), .A2(n_1332), .B(n_1333), .C(n_1339), .Y(n_1331) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
NOR2xp33_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1328), .Y(n_1326) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1329), .Y(n_1358) );
AOI21xp5_ASAP7_75t_L g1367 ( .A1(n_1361), .A2(n_1368), .B(n_1369), .Y(n_1367) );
INVxp67_ASAP7_75t_SL g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
HB1xp67_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
HB1xp67_ASAP7_75t_L g1436 ( .A(n_1376), .Y(n_1436) );
AND3x1_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1394), .C(n_1396), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1377 ( .A(n_1378), .B(n_1387), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .Y(n_1387) );
OAI221xp5_ASAP7_75t_L g1398 ( .A1(n_1389), .A2(n_1393), .B1(n_1399), .B2(n_1400), .C(n_1404), .Y(n_1398) );
OAI31xp33_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1408), .A3(n_1420), .B(n_1421), .Y(n_1396) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
OAI22xp5_ASAP7_75t_L g1415 ( .A1(n_1416), .A2(n_1417), .B1(n_1418), .B2(n_1419), .Y(n_1415) );
BUFx8_ASAP7_75t_SL g1421 ( .A(n_1422), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g1423 ( .A(n_1424), .Y(n_1423) );
BUFx2_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
CKINVDCx5p33_ASAP7_75t_R g1430 ( .A(n_1431), .Y(n_1430) );
A2O1A1Ixp33_ASAP7_75t_L g1438 ( .A1(n_1432), .A2(n_1439), .B(n_1441), .C(n_1442), .Y(n_1438) );
INVxp33_ASAP7_75t_SL g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
HB1xp67_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
endmodule