module real_aes_17445_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g113 ( .A(n_0), .B(n_114), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_1), .A2(n_4), .B1(n_265), .B2(n_266), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_2), .A2(n_43), .B1(n_166), .B2(n_214), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_3), .A2(n_25), .B1(n_214), .B2(n_248), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_5), .A2(n_17), .B1(n_515), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_6), .A2(n_60), .B1(n_151), .B2(n_152), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_7), .A2(n_18), .B1(n_166), .B2(n_167), .Y(n_165) );
INVx1_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_9), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_10), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_11), .A2(n_19), .B1(n_516), .B2(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_12), .A2(n_127), .B1(n_791), .B2(n_792), .Y(n_126) );
INVx1_ASAP7_75t_L g791 ( .A(n_12), .Y(n_791) );
OR2x2_ASAP7_75t_L g106 ( .A(n_13), .B(n_38), .Y(n_106) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_14), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_15), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_16), .A2(n_100), .B1(n_115), .B2(n_823), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_20), .A2(n_96), .B1(n_266), .B2(n_515), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_21), .A2(n_39), .B1(n_144), .B2(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_22), .B(n_142), .Y(n_576) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_23), .A2(n_58), .B(n_157), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_24), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_26), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_27), .B(n_139), .Y(n_206) );
INVx4_ASAP7_75t_R g190 ( .A(n_28), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_29), .A2(n_47), .B1(n_170), .B2(n_263), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_30), .A2(n_54), .B1(n_170), .B2(n_515), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_31), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_32), .B(n_540), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_33), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_34), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g270 ( .A(n_35), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_36), .A2(n_138), .B(n_166), .C(n_246), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_37), .A2(n_55), .B1(n_166), .B2(n_170), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_40), .A2(n_84), .B1(n_166), .B2(n_507), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_41), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_806) );
INVx1_ASAP7_75t_L g809 ( .A(n_41), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_42), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_44), .A2(n_46), .B1(n_166), .B2(n_167), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_45), .A2(n_59), .B1(n_515), .B2(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g210 ( .A(n_48), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_49), .B(n_166), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_50), .Y(n_224) );
INVx2_ASAP7_75t_L g121 ( .A(n_51), .Y(n_121) );
INVx1_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
BUFx3_ASAP7_75t_L g124 ( .A(n_52), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_53), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_56), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_57), .A2(n_85), .B1(n_166), .B2(n_170), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_61), .A2(n_73), .B1(n_263), .B2(n_532), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_62), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_63), .A2(n_76), .B1(n_166), .B2(n_167), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_64), .A2(n_95), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g157 ( .A(n_65), .Y(n_157) );
AND2x4_ASAP7_75t_L g160 ( .A(n_66), .B(n_161), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_67), .A2(n_87), .B1(n_170), .B2(n_263), .Y(n_262) );
AO22x1_ASAP7_75t_L g140 ( .A1(n_68), .A2(n_74), .B1(n_141), .B2(n_144), .Y(n_140) );
INVx1_ASAP7_75t_L g161 ( .A(n_69), .Y(n_161) );
AND2x2_ASAP7_75t_L g249 ( .A(n_70), .B(n_202), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_71), .B(n_151), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_72), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_75), .B(n_214), .Y(n_225) );
INVx2_ASAP7_75t_L g139 ( .A(n_77), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_78), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_79), .B(n_202), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_80), .A2(n_94), .B1(n_151), .B2(n_170), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_81), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_82), .B(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_83), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_86), .B(n_202), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_88), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_89), .B(n_202), .Y(n_221) );
INVx1_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_90), .B(n_800), .Y(n_799) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_91), .B(n_142), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_92), .A2(n_151), .B(n_172), .C(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g195 ( .A(n_93), .B(n_196), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g229 ( .A(n_97), .B(n_191), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_98), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g823 ( .A(n_102), .Y(n_823) );
INVx6_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g125 ( .A(n_106), .Y(n_125) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_106), .B(n_124), .Y(n_822) );
NOR2x1p5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND3x2_ASAP7_75t_L g814 ( .A(n_108), .B(n_111), .C(n_125), .Y(n_814) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g800 ( .A(n_109), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g487 ( .A(n_112), .Y(n_487) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_801), .Y(n_115) );
OAI21xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_126), .B(n_793), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x6_ASAP7_75t_SL g119 ( .A(n_120), .B(n_122), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g804 ( .A(n_121), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_121), .B(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_SL g798 ( .A(n_125), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g792 ( .A(n_127), .Y(n_792) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_485), .B1(n_488), .B2(n_790), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_395), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_324), .C(n_366), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_298), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_197), .B1(n_273), .B2(n_284), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_178), .Y(n_134) );
AOI21xp33_ASAP7_75t_L g317 ( .A1(n_135), .A2(n_318), .B(n_320), .Y(n_317) );
AOI21xp33_ASAP7_75t_L g390 ( .A1(n_135), .A2(n_391), .B(n_392), .Y(n_390) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_162), .Y(n_135) );
INVx2_ASAP7_75t_L g310 ( .A(n_136), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_136), .B(n_163), .Y(n_340) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_146), .C(n_158), .Y(n_137) );
INVx6_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_138), .A2(n_229), .B(n_230), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_138), .B(n_140), .Y(n_282) );
O2A1O1Ixp5_ASAP7_75t_L g574 ( .A1(n_138), .A2(n_167), .B(n_575), .C(n_576), .Y(n_574) );
BUFx8_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx1_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
INVx1_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
INVxp67_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g515 ( .A(n_142), .Y(n_515) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g145 ( .A(n_143), .Y(n_145) );
INVx1_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx1_ASAP7_75t_L g153 ( .A(n_143), .Y(n_153) );
INVx3_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_143), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_143), .Y(n_214) );
INVx1_ASAP7_75t_L g242 ( .A(n_143), .Y(n_242) );
INVx2_ASAP7_75t_L g248 ( .A(n_143), .Y(n_248) );
OAI21xp33_ASAP7_75t_SL g205 ( .A1(n_144), .A2(n_206), .B(n_207), .Y(n_205) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g281 ( .A(n_146), .Y(n_281) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B(n_154), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_147), .A2(n_212), .B(n_213), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_147), .A2(n_168), .B1(n_253), .B2(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g498 ( .A(n_148), .Y(n_498) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g227 ( .A(n_149), .Y(n_227) );
INVx1_ASAP7_75t_L g560 ( .A(n_152), .Y(n_560) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_153), .B(n_187), .Y(n_186) );
OAI21xp33_ASAP7_75t_L g158 ( .A1(n_154), .A2(n_155), .B(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx2_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
INVx2_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g283 ( .A(n_158), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_159), .A2(n_238), .B(n_245), .Y(n_237) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx10_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
BUFx10_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
INVx1_ASAP7_75t_L g268 ( .A(n_160), .Y(n_268) );
AND2x2_ASAP7_75t_L g380 ( .A(n_162), .B(n_219), .Y(n_380) );
INVx1_ASAP7_75t_L g413 ( .A(n_162), .Y(n_413) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g275 ( .A(n_163), .B(n_220), .Y(n_275) );
AND2x2_ASAP7_75t_L g306 ( .A(n_163), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g315 ( .A(n_163), .Y(n_315) );
OR2x2_ASAP7_75t_L g334 ( .A(n_163), .B(n_180), .Y(n_334) );
AND2x2_ASAP7_75t_L g349 ( .A(n_163), .B(n_180), .Y(n_349) );
AO31x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_173), .A3(n_174), .B(n_175), .Y(n_163) );
OAI22x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B1(n_169), .B2(n_171), .Y(n_164) );
INVx4_ASAP7_75t_L g167 ( .A(n_166), .Y(n_167) );
INVx1_ASAP7_75t_L g516 ( .A(n_166), .Y(n_516) );
INVx1_ASAP7_75t_L g532 ( .A(n_166), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_167), .A2(n_224), .B(n_225), .C(n_226), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_168), .A2(n_171), .B1(n_262), .B2(n_264), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_168), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_168), .A2(n_171), .B1(n_506), .B2(n_508), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_168), .A2(n_514), .B1(n_517), .B2(n_518), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_168), .A2(n_498), .B1(n_530), .B2(n_531), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_168), .A2(n_498), .B1(n_539), .B2(n_541), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_168), .A2(n_498), .B1(n_549), .B2(n_550), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_168), .A2(n_518), .B1(n_559), .B2(n_561), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_168), .A2(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_170), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g265 ( .A(n_170), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_171), .B(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_SL g518 ( .A(n_172), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_173), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_173), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g194 ( .A(n_174), .Y(n_194) );
AO31x2_ASAP7_75t_L g495 ( .A1(n_174), .A2(n_255), .A3(n_496), .B(n_500), .Y(n_495) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_174), .A2(n_504), .A3(n_538), .B(n_543), .Y(n_537) );
AO31x2_ASAP7_75t_L g557 ( .A1(n_174), .A2(n_236), .A3(n_558), .B(n_562), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVx2_ASAP7_75t_L g196 ( .A(n_177), .Y(n_196) );
BUFx2_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_177), .B(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_177), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_179), .B(n_348), .Y(n_391) );
OR2x2_ASAP7_75t_L g479 ( .A(n_179), .B(n_340), .Y(n_479) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g307 ( .A(n_180), .Y(n_307) );
AND2x2_ASAP7_75t_L g316 ( .A(n_180), .B(n_279), .Y(n_316) );
AND2x2_ASAP7_75t_L g319 ( .A(n_180), .B(n_220), .Y(n_319) );
AND2x2_ASAP7_75t_L g338 ( .A(n_180), .B(n_219), .Y(n_338) );
AND2x4_ASAP7_75t_L g357 ( .A(n_180), .B(n_280), .Y(n_357) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B(n_195), .Y(n_180) );
AO31x2_ASAP7_75t_L g528 ( .A1(n_181), .A2(n_519), .A3(n_529), .B(n_533), .Y(n_528) );
AO31x2_ASAP7_75t_L g547 ( .A1(n_181), .A2(n_267), .A3(n_548), .B(n_551), .Y(n_547) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_183), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_SL g562 ( .A(n_183), .B(n_563), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B(n_194), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_189) );
INVx2_ASAP7_75t_L g263 ( .A(n_191), .Y(n_263) );
INVx1_ASAP7_75t_L g540 ( .A(n_191), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_192), .Y(n_542) );
INVx1_ASAP7_75t_L g519 ( .A(n_194), .Y(n_519) );
OAI21xp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_217), .B(n_258), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_198), .B(n_352), .Y(n_455) );
CKINVDCx14_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_200), .B(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g288 ( .A(n_200), .Y(n_288) );
OR2x2_ASAP7_75t_L g296 ( .A(n_200), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_200), .B(n_289), .Y(n_321) );
AND2x2_ASAP7_75t_L g346 ( .A(n_200), .B(n_260), .Y(n_346) );
AND2x2_ASAP7_75t_L g364 ( .A(n_200), .B(n_294), .Y(n_364) );
INVx1_ASAP7_75t_L g403 ( .A(n_200), .Y(n_403) );
AND2x2_ASAP7_75t_L g405 ( .A(n_200), .B(n_406), .Y(n_405) );
NAND2x1p5_ASAP7_75t_SL g424 ( .A(n_200), .B(n_345), .Y(n_424) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_204), .Y(n_200) );
NOR2x1_ASAP7_75t_L g231 ( .A(n_202), .B(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g255 ( .A(n_202), .Y(n_255) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g215 ( .A(n_203), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_203), .B(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g504 ( .A(n_203), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_203), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_203), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g572 ( .A(n_203), .Y(n_572) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_211), .B(n_215), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
BUFx4f_ASAP7_75t_L g244 ( .A(n_209), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_214), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g232 ( .A(n_216), .Y(n_232) );
AO31x2_ASAP7_75t_L g251 ( .A1(n_216), .A2(n_252), .A3(n_255), .B(n_256), .Y(n_251) );
OAI32xp33_ASAP7_75t_L g308 ( .A1(n_217), .A2(n_300), .A3(n_309), .B1(n_311), .B2(n_313), .Y(n_308) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_233), .Y(n_217) );
INVx1_ASAP7_75t_L g348 ( .A(n_218), .Y(n_348) );
AND2x2_ASAP7_75t_L g356 ( .A(n_218), .B(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g355 ( .A(n_219), .B(n_279), .Y(n_355) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx3_ASAP7_75t_L g305 ( .A(n_220), .Y(n_305) );
AND2x2_ASAP7_75t_L g314 ( .A(n_220), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g420 ( .A(n_220), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_228), .B(n_231), .Y(n_222) );
INVx2_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g290 ( .A(n_233), .Y(n_290) );
OR2x2_ASAP7_75t_L g300 ( .A(n_233), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g422 ( .A(n_233), .Y(n_422) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_250), .Y(n_233) );
AND2x2_ASAP7_75t_L g323 ( .A(n_234), .B(n_251), .Y(n_323) );
INVx2_ASAP7_75t_L g345 ( .A(n_234), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_234), .B(n_260), .Y(n_365) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g272 ( .A(n_235), .Y(n_272) );
AOI21x1_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_249), .Y(n_235) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_236), .A2(n_261), .A3(n_267), .B(n_269), .Y(n_260) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_236), .A2(n_513), .A3(n_519), .B(n_520), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_241), .B(n_244), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_SL g507 ( .A(n_248), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_250), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g354 ( .A(n_250), .Y(n_354) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
OR2x2_ASAP7_75t_L g360 ( .A(n_251), .B(n_260), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_251), .B(n_260), .Y(n_393) );
INVx2_ASAP7_75t_L g341 ( .A(n_258), .Y(n_341) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_271), .Y(n_258) );
OR2x2_ASAP7_75t_L g328 ( .A(n_259), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g406 ( .A(n_259), .Y(n_406) );
INVx1_ASAP7_75t_L g289 ( .A(n_260), .Y(n_289) );
INVx1_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
INVx1_ASAP7_75t_L g312 ( .A(n_260), .Y(n_312) );
AO31x2_ASAP7_75t_L g503 ( .A1(n_267), .A2(n_504), .A3(n_505), .B(n_509), .Y(n_503) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g580 ( .A(n_268), .Y(n_580) );
OR2x2_ASAP7_75t_L g416 ( .A(n_271), .B(n_393), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_272), .B(n_288), .Y(n_329) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_272), .Y(n_331) );
OR2x2_ASAP7_75t_L g430 ( .A(n_272), .B(n_354), .Y(n_430) );
INVxp67_ASAP7_75t_L g454 ( .A(n_272), .Y(n_454) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NAND2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_275), .B(n_316), .Y(n_383) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g332 ( .A(n_277), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g445 ( .A(n_278), .Y(n_445) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g474 ( .A(n_279), .B(n_307), .Y(n_474) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g400 ( .A(n_280), .B(n_307), .Y(n_400) );
AOI21x1_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_291), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_287), .B(n_323), .Y(n_437) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g301 ( .A(n_288), .Y(n_301) );
AND2x2_ASAP7_75t_L g351 ( .A(n_288), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_288), .B(n_345), .Y(n_394) );
OR2x2_ASAP7_75t_L g466 ( .A(n_288), .B(n_353), .Y(n_466) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g386 ( .A(n_292), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx2_ASAP7_75t_L g377 ( .A(n_293), .Y(n_377) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g367 ( .A(n_296), .B(n_368), .Y(n_367) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_296), .Y(n_378) );
OR2x2_ASAP7_75t_L g429 ( .A(n_296), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g484 ( .A(n_296), .Y(n_484) );
AOI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B(n_308), .C(n_317), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g373 ( .A(n_301), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_301), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g446 ( .A(n_301), .B(n_323), .Y(n_446) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_304), .B(n_349), .Y(n_371) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_304), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g456 ( .A(n_304), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g399 ( .A(n_305), .Y(n_399) );
AND2x2_ASAP7_75t_L g427 ( .A(n_306), .B(n_355), .Y(n_427) );
INVx2_ASAP7_75t_L g450 ( .A(n_306), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_306), .B(n_348), .Y(n_482) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_309), .B(n_314), .Y(n_436) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g389 ( .A(n_310), .B(n_315), .Y(n_389) );
OR2x2_ASAP7_75t_L g441 ( .A(n_310), .B(n_334), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_311), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_311), .B(n_323), .Y(n_477) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g425 ( .A(n_312), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g408 ( .A(n_314), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_314), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g458 ( .A(n_315), .Y(n_458) );
BUFx2_ASAP7_75t_L g326 ( .A(n_316), .Y(n_326) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g444 ( .A(n_319), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g368 ( .A(n_323), .Y(n_368) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_323), .Y(n_385) );
NAND3xp33_ASAP7_75t_SL g324 ( .A(n_325), .B(n_335), .C(n_350), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_327), .B1(n_330), .B2(n_332), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_332), .A2(n_358), .B1(n_439), .B2(n_442), .C1(n_444), .C2(n_446), .Y(n_438) );
AND2x2_ASAP7_75t_L g470 ( .A(n_333), .B(n_419), .Y(n_470) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g418 ( .A(n_334), .B(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_341), .B1(n_342), .B2(n_347), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx2_ASAP7_75t_SL g414 ( .A(n_338), .Y(n_414) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
AND2x2_ASAP7_75t_L g401 ( .A(n_343), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g359 ( .A(n_344), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g353 ( .A(n_345), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g468 ( .A(n_346), .Y(n_468) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_349), .B(n_445), .Y(n_464) );
INVx1_ASAP7_75t_L g481 ( .A(n_349), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B1(n_356), .B2(n_358), .C1(n_361), .C2(n_362), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_357), .Y(n_361) );
AND2x2_ASAP7_75t_L g379 ( .A(n_357), .B(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g410 ( .A(n_357), .Y(n_410) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g374 ( .A(n_360), .Y(n_374) );
OR2x2_ASAP7_75t_L g443 ( .A(n_360), .B(n_424), .Y(n_443) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_372), .C(n_381), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B(n_379), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_373), .A2(n_411), .B1(n_460), .B2(n_463), .C(n_465), .Y(n_459) );
AND2x4_ASAP7_75t_L g402 ( .A(n_374), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
AOI211x1_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_386), .C(n_390), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g451 ( .A(n_389), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_392), .B(n_440), .C(n_441), .Y(n_439) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g475 ( .A(n_393), .Y(n_475) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_396), .B(n_447), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g396 ( .A(n_397), .B(n_404), .C(n_426), .D(n_438), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
AND2x2_ASAP7_75t_L g457 ( .A(n_400), .B(n_458), .Y(n_457) );
AOI221x1_ASAP7_75t_L g426 ( .A1(n_402), .A2(n_427), .B1(n_428), .B2(n_431), .C(n_434), .Y(n_426) );
AND2x2_ASAP7_75t_L g452 ( .A(n_402), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g462 ( .A(n_403), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_411), .B2(n_415), .C(n_417), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_409), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_414), .A2(n_418), .B1(n_421), .B2(n_423), .Y(n_417) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_418), .A2(n_435), .B(n_437), .Y(n_434) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g440 ( .A(n_420), .Y(n_440) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g461 ( .A(n_430), .Y(n_461) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_443), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_459), .C(n_471), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_452), .B1(n_455), .B2(n_456), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g467 ( .A(n_454), .B(n_468), .Y(n_467) );
NAND2x1_ASAP7_75t_L g483 ( .A(n_454), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_469), .Y(n_465) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B1(n_476), .B2(n_478), .C(n_480), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
INVx4_ASAP7_75t_L g790 ( .A(n_485), .Y(n_790) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g821 ( .A(n_487), .B(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g808 ( .A(n_488), .Y(n_808) );
NOR2x1p5_ASAP7_75t_L g488 ( .A(n_489), .B(n_700), .Y(n_488) );
NAND4xp75_ASAP7_75t_L g489 ( .A(n_490), .B(n_645), .C(n_665), .D(n_681), .Y(n_489) );
NOR2x1p5_ASAP7_75t_SL g490 ( .A(n_491), .B(n_615), .Y(n_490) );
NAND4xp75_ASAP7_75t_L g491 ( .A(n_492), .B(n_553), .C(n_592), .D(n_601), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_522), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_502), .Y(n_493) );
AND2x4_ASAP7_75t_L g725 ( .A(n_494), .B(n_652), .Y(n_725) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_495), .Y(n_568) );
INVx2_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
AND2x2_ASAP7_75t_L g609 ( .A(n_495), .B(n_571), .Y(n_609) );
OR2x2_ASAP7_75t_L g664 ( .A(n_495), .B(n_503), .Y(n_664) );
AND2x2_ASAP7_75t_L g582 ( .A(n_502), .B(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g732 ( .A(n_502), .B(n_609), .Y(n_732) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_511), .Y(n_502) );
OR2x2_ASAP7_75t_L g569 ( .A(n_503), .B(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g600 ( .A(n_503), .Y(n_600) );
AND2x2_ASAP7_75t_L g606 ( .A(n_503), .B(n_512), .Y(n_606) );
INVx1_ASAP7_75t_L g624 ( .A(n_503), .Y(n_624) );
INVx2_ASAP7_75t_L g653 ( .A(n_503), .Y(n_653) );
INVx3_ASAP7_75t_L g629 ( .A(n_511), .Y(n_629) );
INVx2_ASAP7_75t_L g634 ( .A(n_511), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_511), .B(n_585), .Y(n_639) );
AND2x2_ASAP7_75t_L g662 ( .A(n_511), .B(n_641), .Y(n_662) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_511), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_511), .B(n_717), .Y(n_716) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g651 ( .A(n_512), .Y(n_651) );
AND2x2_ASAP7_75t_L g699 ( .A(n_512), .B(n_653), .Y(n_699) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_524), .B(n_643), .Y(n_690) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_525), .B(n_643), .Y(n_687) );
INVx1_ASAP7_75t_L g788 ( .A(n_525), .Y(n_788) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g738 ( .A(n_526), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g591 ( .A(n_527), .Y(n_591) );
OR2x2_ASAP7_75t_L g672 ( .A(n_527), .B(n_546), .Y(n_672) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g614 ( .A(n_528), .Y(n_614) );
AND2x4_ASAP7_75t_L g620 ( .A(n_528), .B(n_621), .Y(n_620) );
AOI32xp33_ASAP7_75t_L g758 ( .A1(n_535), .A2(n_661), .A3(n_759), .B1(n_761), .B2(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g707 ( .A(n_536), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .Y(n_536) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_537), .Y(n_555) );
OR2x2_ASAP7_75t_L g589 ( .A(n_537), .B(n_547), .Y(n_589) );
INVx1_ASAP7_75t_L g604 ( .A(n_537), .Y(n_604) );
AND2x2_ASAP7_75t_L g613 ( .A(n_537), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g619 ( .A(n_537), .Y(n_619) );
INVx2_ASAP7_75t_L g644 ( .A(n_537), .Y(n_644) );
AND2x2_ASAP7_75t_L g763 ( .A(n_537), .B(n_557), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_545), .B(n_596), .Y(n_683) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g556 ( .A(n_547), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g612 ( .A(n_547), .Y(n_612) );
INVx2_ASAP7_75t_L g621 ( .A(n_547), .Y(n_621) );
AND2x4_ASAP7_75t_L g643 ( .A(n_547), .B(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_547), .Y(n_735) );
AOI22x1_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_564), .B1(n_582), .B2(n_587), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_556), .B(n_713), .C(n_714), .D(n_715), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_556), .B(n_613), .Y(n_743) );
INVx4_ASAP7_75t_SL g596 ( .A(n_557), .Y(n_596) );
BUFx2_ASAP7_75t_L g659 ( .A(n_557), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_557), .B(n_604), .Y(n_722) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g684 ( .A(n_566), .B(n_633), .Y(n_684) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g607 ( .A(n_570), .B(n_585), .Y(n_607) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_571), .B(n_586), .Y(n_631) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B(n_581), .Y(n_571) );
OAI21x1_ASAP7_75t_L g626 ( .A1(n_572), .A2(n_573), .B(n_581), .Y(n_626) );
OAI21x1_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .B(n_580), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_583), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g649 ( .A(n_583), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g688 ( .A(n_584), .B(n_606), .Y(n_688) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g731 ( .A(n_586), .B(n_641), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_587), .A2(n_704), .B1(n_706), .B2(n_709), .C(n_711), .Y(n_703) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g597 ( .A(n_589), .Y(n_597) );
OR2x2_ASAP7_75t_L g697 ( .A(n_589), .B(n_636), .Y(n_697) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_598), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_593), .A2(n_719), .B1(n_723), .B2(n_726), .Y(n_718) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .Y(n_593) );
AND2x4_ASAP7_75t_L g642 ( .A(n_594), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g754 ( .A(n_594), .B(n_672), .Y(n_754) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g602 ( .A(n_596), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g618 ( .A(n_596), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g677 ( .A(n_596), .B(n_614), .Y(n_677) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_596), .Y(n_694) );
INVx1_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_596), .B(n_621), .Y(n_751) );
AND2x4_ASAP7_75t_L g658 ( .A(n_597), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g656 ( .A(n_599), .Y(n_656) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_600), .B(n_641), .Y(n_640) );
NAND2x1_ASAP7_75t_L g760 ( .A(n_600), .B(n_662), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B1(n_608), .B2(n_610), .Y(n_601) );
AND2x2_ASAP7_75t_L g627 ( .A(n_602), .B(n_620), .Y(n_627) );
INVx1_ASAP7_75t_L g668 ( .A(n_602), .Y(n_668) );
AND2x2_ASAP7_75t_L g775 ( .A(n_602), .B(n_636), .Y(n_775) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_SL g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g608 ( .A(n_606), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g748 ( .A(n_606), .Y(n_748) );
AND2x2_ASAP7_75t_L g765 ( .A(n_606), .B(n_625), .Y(n_765) );
AND2x2_ASAP7_75t_L g781 ( .A(n_606), .B(n_731), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_607), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g704 ( .A(n_607), .B(n_705), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_607), .A2(n_697), .B1(n_712), .B2(n_716), .Y(n_711) );
INVx1_ASAP7_75t_L g667 ( .A(n_609), .Y(n_667) );
AND2x2_ASAP7_75t_L g698 ( .A(n_609), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_609), .B(n_705), .Y(n_727) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g733 ( .A(n_613), .B(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_613), .A2(n_637), .B1(n_742), .B2(n_744), .Y(n_741) );
INVx3_ASAP7_75t_L g636 ( .A(n_614), .Y(n_636) );
AND2x2_ASAP7_75t_L g768 ( .A(n_614), .B(n_621), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_632), .Y(n_615) );
AOI32xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_622), .A3(n_625), .B1(n_627), .B2(n_628), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_619), .Y(n_714) );
INVx1_ASAP7_75t_L g739 ( .A(n_619), .Y(n_739) );
INVx3_ASAP7_75t_L g695 ( .A(n_620), .Y(n_695) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_623), .A2(n_771), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_770) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g747 ( .A(n_625), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g783 ( .A(n_625), .B(n_744), .Y(n_783) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g641 ( .A(n_626), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_628), .B(n_656), .Y(n_655) );
AO22x1_ASAP7_75t_L g685 ( .A1(n_628), .A2(n_686), .B1(n_688), .B2(n_689), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g789 ( .A(n_628), .B(n_656), .Y(n_789) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx2_ASAP7_75t_L g705 ( .A(n_629), .Y(n_705) );
INVx1_ASAP7_75t_L g715 ( .A(n_629), .Y(n_715) );
AND2x2_ASAP7_75t_L g635 ( .A(n_630), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_SL g717 ( .A(n_631), .Y(n_717) );
INVx1_ASAP7_75t_L g757 ( .A(n_631), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_637), .C(n_642), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR2x1p5_ASAP7_75t_L g744 ( .A(n_634), .B(n_664), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_635), .B(n_694), .Y(n_771) );
AOI31xp33_ASAP7_75t_L g654 ( .A1(n_636), .A2(n_655), .A3(n_657), .B(n_660), .Y(n_654) );
INVx4_ASAP7_75t_L g713 ( .A(n_636), .Y(n_713) );
OR2x2_ASAP7_75t_L g750 ( .A(n_636), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
AND2x4_ASAP7_75t_L g652 ( .A(n_641), .B(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_643), .Y(n_648) );
AND2x2_ASAP7_75t_L g679 ( .A(n_643), .B(n_677), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g645 ( .A(n_646), .B(n_654), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g772 ( .A(n_649), .Y(n_772) );
INVx1_ASAP7_75t_L g680 ( .A(n_650), .Y(n_680) );
AND2x4_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g710 ( .A(n_651), .Y(n_710) );
AND2x2_ASAP7_75t_L g709 ( .A(n_652), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI322xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .A3(n_669), .B1(n_673), .B2(n_676), .C1(n_678), .C2(n_680), .Y(n_666) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI211x1_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B(n_685), .C(n_691), .Y(n_681) );
INVx1_ASAP7_75t_L g786 ( .A(n_682), .Y(n_786) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g740 ( .A(n_684), .Y(n_740) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OA21x2_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_696), .B(n_698), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx2_ASAP7_75t_L g761 ( .A(n_695), .Y(n_761) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp33_ASAP7_75t_L g756 ( .A(n_699), .B(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_769), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_736), .C(n_752), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_718), .C(n_728), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_705), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g764 ( .A1(n_709), .A2(n_765), .B(n_766), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_713), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_713), .B(n_763), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_714), .B(n_788), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_715), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_725), .A2(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_732), .B(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_740), .B(n_741), .C(n_745), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_SL g755 ( .A(n_747), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_751), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_755), .B(n_758), .C(n_764), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_763), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g784 ( .A(n_763), .Y(n_784) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g780 ( .A(n_768), .Y(n_780) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_778), .C(n_785), .Y(n_769) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AOI21xp33_ASAP7_75t_SL g778 ( .A1(n_779), .A2(n_782), .B(n_784), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI21xp33_ASAP7_75t_R g785 ( .A1(n_786), .A2(n_787), .B(n_789), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g805 ( .A1(n_793), .A2(n_806), .B(n_810), .Y(n_805) );
INVxp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
BUFx12f_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx4_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AO21x1_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_805), .B(n_815), .Y(n_801) );
CKINVDCx11_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx4_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
BUFx10_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
endmodule