module fake_jpeg_30686_n_109 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_52),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_37),
.B1(n_33),
.B2(n_39),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_6),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_64),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_42),
.B(n_41),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_3),
.B(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_7),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_39),
.B1(n_43),
.B2(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_44),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_49),
.B1(n_50),
.B2(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_75),
.B1(n_67),
.B2(n_57),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_76),
.B(n_10),
.C(n_12),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_48),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_72),
.B(n_32),
.C(n_20),
.Y(n_90)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_8),
.Y(n_80)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_6),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_8),
.B(n_9),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_85),
.B1(n_90),
.B2(n_24),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_10),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_84),
.B(n_23),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_14),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_18),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_16),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_95),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_92),
.B(n_82),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_102),
.B(n_92),
.Y(n_103)
);

AOI21x1_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_79),
.B(n_100),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_93),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_79),
.B(n_91),
.C(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_89),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_31),
.Y(n_109)
);


endmodule