module fake_netlist_6_1956_n_770 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_770);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_770;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_758;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_527;
wire n_608;
wire n_261;
wire n_474;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx3_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_66),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_27),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_38),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_80),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_21),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_0),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_18),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_53),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

BUFx8_ASAP7_75t_SL g162 ( 
.A(n_96),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_86),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_84),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_42),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_32),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_93),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_67),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_19),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_7),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_110),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_22),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_63),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_68),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_69),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_24),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_56),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_82),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_94),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_19),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_138),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_5),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_106),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_59),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_142),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_0),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_1),
.Y(n_207)
);

BUFx8_ASAP7_75t_SL g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_160),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_179),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_185),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_156),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_146),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_149),
.B(n_1),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_2),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_158),
.B(n_2),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_150),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_204),
.B1(n_229),
.B2(n_186),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_197),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_214),
.B1(n_236),
.B2(n_212),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_3),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_150),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_151),
.B1(n_198),
.B2(n_152),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_151),
.B1(n_198),
.B2(n_152),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_153),
.B1(n_155),
.B2(n_200),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_153),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_155),
.Y(n_257)
);

AO22x2_ASAP7_75t_L g258 ( 
.A1(n_201),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_208),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_211),
.A2(n_195),
.B1(n_191),
.B2(n_188),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_180),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

BUFx6f_ASAP7_75t_SL g263 ( 
.A(n_201),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_211),
.A2(n_183),
.B1(n_181),
.B2(n_7),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_201),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_237),
.A2(n_216),
.B1(n_218),
.B2(n_226),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_270)
);

AO22x2_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_202),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_216),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_L g276 ( 
.A1(n_218),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_226),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_277)
);

AO22x2_ASAP7_75t_L g278 ( 
.A1(n_226),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_278)
);

AO22x2_ASAP7_75t_L g279 ( 
.A1(n_209),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_209),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_231),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_205),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_228),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_231),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_203),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_231),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_230),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_241),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_249),
.B(n_230),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_232),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_232),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_252),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_232),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_259),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_248),
.B(n_234),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_234),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_234),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_246),
.B(n_35),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_251),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_255),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_227),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_227),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_243),
.B(n_227),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_245),
.B(n_206),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_245),
.B(n_247),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_259),
.B(n_227),
.Y(n_327)
);

OR2x6_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_255),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_278),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_268),
.B(n_206),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_268),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_279),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_228),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_281),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_276),
.B(n_228),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_270),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g354 ( 
.A(n_329),
.B(n_203),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_228),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g359 ( 
.A1(n_317),
.A2(n_221),
.B(n_217),
.Y(n_359)
);

AND2x4_ASAP7_75t_SL g360 ( 
.A(n_312),
.B(n_228),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_228),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_297),
.B(n_205),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_206),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_288),
.B(n_213),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_293),
.B(n_219),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_219),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_293),
.B(n_219),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_322),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_298),
.B(n_205),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

AND2x4_ASAP7_75t_SL g377 ( 
.A(n_312),
.B(n_328),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_315),
.B(n_205),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_302),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_307),
.B(n_36),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_338),
.B(n_215),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_303),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_290),
.Y(n_386)
);

OR2x4_ASAP7_75t_L g387 ( 
.A(n_296),
.B(n_203),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_305),
.B(n_213),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g389 ( 
.A(n_330),
.B(n_203),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_305),
.B(n_215),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_314),
.B(n_39),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_304),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_315),
.B(n_205),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g394 ( 
.A(n_323),
.B(n_203),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_205),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_326),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_205),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_325),
.B(n_40),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_215),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_341),
.B(n_213),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_41),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_341),
.B(n_222),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_347),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_299),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_334),
.B(n_222),
.Y(n_407)
);

BUFx4_ASAP7_75t_SL g408 ( 
.A(n_313),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_331),
.B(n_43),
.Y(n_409)
);

BUFx4f_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_309),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_294),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_345),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_345),
.B(n_215),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_326),
.B(n_225),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_332),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_340),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_344),
.B(n_217),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_346),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_364),
.B(n_291),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_334),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_333),
.Y(n_423)
);

BUFx4f_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_374),
.B(n_342),
.Y(n_425)
);

BUFx12f_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

AND2x2_ASAP7_75t_SL g427 ( 
.A(n_365),
.B(n_349),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_410),
.B(n_328),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_335),
.Y(n_430)
);

OR2x6_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_398),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_364),
.B(n_367),
.Y(n_432)
);

OR2x6_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_350),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_404),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_339),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_343),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_44),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_372),
.B(n_343),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_367),
.B(n_222),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_370),
.B(n_327),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_372),
.B(n_217),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_398),
.B(n_217),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_370),
.B(n_384),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_398),
.B(n_224),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_417),
.Y(n_452)
);

BUFx12f_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_402),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_224),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_368),
.Y(n_458)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_410),
.B(n_221),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_353),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

BUFx12f_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_369),
.B(n_221),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_384),
.B(n_221),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_416),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_356),
.B(n_224),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_355),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_354),
.B(n_225),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_391),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_352),
.B(n_45),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_409),
.B(n_239),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_352),
.B(n_239),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_396),
.B(n_225),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_354),
.B(n_225),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_409),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_389),
.B(n_225),
.Y(n_476)
);

BUFx2_ASAP7_75t_SL g477 ( 
.A(n_435),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_427),
.A2(n_418),
.B1(n_399),
.B2(n_390),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_421),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

BUFx2_ASAP7_75t_SL g485 ( 
.A(n_439),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_444),
.Y(n_487)
);

BUFx12f_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_442),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_453),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_422),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_432),
.B(n_399),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_465),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_462),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_420),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_460),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_445),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_458),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

BUFx12f_ASAP7_75t_L g502 ( 
.A(n_425),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_436),
.B(n_418),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_434),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_464),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_461),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_475),
.B(n_396),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_448),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_448),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

NAND2x1p5_ASAP7_75t_L g518 ( 
.A(n_438),
.B(n_396),
.Y(n_518)
);

CKINVDCx6p67_ASAP7_75t_R g519 ( 
.A(n_449),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_469),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_482),
.A2(n_428),
.B1(n_436),
.B2(n_443),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_479),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_481),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_502),
.A2(n_428),
.B1(n_459),
.B2(n_433),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_509),
.A2(n_361),
.B(n_358),
.Y(n_528)
);

CKINVDCx11_ASAP7_75t_R g529 ( 
.A(n_488),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_425),
.B1(n_438),
.B2(n_433),
.Y(n_530)
);

BUFx2_ASAP7_75t_SL g531 ( 
.A(n_495),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_497),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_500),
.Y(n_533)
);

BUFx2_ASAP7_75t_SL g534 ( 
.A(n_496),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_489),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_502),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_516),
.A2(n_433),
.B1(n_423),
.B2(n_400),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_480),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_483),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_516),
.A2(n_423),
.B1(n_403),
.B2(n_407),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_SL g541 ( 
.A1(n_492),
.A2(n_472),
.B1(n_457),
.B2(n_388),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_516),
.A2(n_423),
.B1(n_429),
.B2(n_469),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_492),
.A2(n_394),
.B1(n_389),
.B2(n_449),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_500),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_478),
.A2(n_452),
.B1(n_437),
.B2(n_394),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_514),
.B(n_505),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_500),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_510),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_492),
.A2(n_449),
.B1(n_447),
.B2(n_466),
.Y(n_551)
);

CKINVDCx11_ASAP7_75t_R g552 ( 
.A(n_488),
.Y(n_552)
);

OAI21xp33_ASAP7_75t_SL g553 ( 
.A1(n_515),
.A2(n_430),
.B(n_437),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_489),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_518),
.A2(n_368),
.B(n_419),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_498),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_515),
.B(n_440),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_491),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_518),
.A2(n_452),
.B1(n_430),
.B2(n_410),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_491),
.A2(n_382),
.B1(n_471),
.B2(n_507),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_512),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_493),
.A2(n_423),
.B1(n_391),
.B2(n_447),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_523),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_541),
.A2(n_382),
.B(n_441),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_522),
.A2(n_493),
.B1(n_512),
.B2(n_509),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_530),
.A2(n_518),
.B1(n_471),
.B2(n_506),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_532),
.B(n_492),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_525),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_560),
.A2(n_531),
.B1(n_545),
.B2(n_559),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_543),
.A2(n_509),
.B1(n_487),
.B2(n_494),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_534),
.A2(n_447),
.B1(n_471),
.B2(n_506),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_526),
.Y(n_573)
);

NOR2x1_ASAP7_75t_R g574 ( 
.A(n_529),
.B(n_446),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_538),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_538),
.A2(n_447),
.B1(n_506),
.B2(n_505),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

BUFx4f_ASAP7_75t_SL g578 ( 
.A(n_558),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_536),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_527),
.A2(n_487),
.B1(n_494),
.B2(n_463),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_557),
.B(n_517),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_546),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_548),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_536),
.A2(n_505),
.B1(n_520),
.B2(n_510),
.Y(n_584)
);

AOI222xp33_ASAP7_75t_L g585 ( 
.A1(n_553),
.A2(n_440),
.B1(n_455),
.B2(n_390),
.C1(n_405),
.C2(n_239),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_540),
.A2(n_519),
.B1(n_501),
.B2(n_514),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_546),
.B(n_514),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_535),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_558),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_551),
.A2(n_519),
.B1(n_501),
.B2(n_521),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_529),
.Y(n_592)
);

INVx5_ASAP7_75t_SL g593 ( 
.A(n_546),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_549),
.A2(n_470),
.B1(n_454),
.B2(n_405),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_549),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_537),
.A2(n_542),
.B1(n_510),
.B2(n_520),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_562),
.A2(n_521),
.B1(n_520),
.B2(n_510),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_528),
.A2(n_377),
.B(n_360),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_533),
.A2(n_377),
.B(n_360),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_549),
.A2(n_387),
.B1(n_513),
.B2(n_520),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_533),
.A2(n_408),
.B(n_513),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

BUFx12f_ASAP7_75t_L g607 ( 
.A(n_552),
.Y(n_607)
);

OAI21xp33_ASAP7_75t_L g608 ( 
.A1(n_555),
.A2(n_355),
.B(n_392),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_556),
.A2(n_521),
.B1(n_520),
.B2(n_511),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_556),
.A2(n_521),
.B1(n_520),
.B2(n_511),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_585),
.B(n_521),
.C(n_510),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_563),
.B(n_550),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_570),
.A2(n_511),
.B1(n_521),
.B2(n_510),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_SL g614 ( 
.A1(n_567),
.A2(n_511),
.B1(n_513),
.B2(n_547),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_565),
.B(n_554),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_SL g616 ( 
.A1(n_564),
.A2(n_511),
.B(n_397),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_568),
.A2(n_511),
.B1(n_544),
.B2(n_547),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_581),
.B(n_554),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_580),
.A2(n_385),
.B1(n_411),
.B2(n_381),
.Y(n_619)
);

OAI21xp33_ASAP7_75t_L g620 ( 
.A1(n_580),
.A2(n_386),
.B(n_412),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_566),
.A2(n_412),
.B1(n_386),
.B2(n_419),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_569),
.B(n_539),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_566),
.A2(n_498),
.B1(n_395),
.B2(n_375),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_568),
.A2(n_581),
.B1(n_578),
.B2(n_607),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_571),
.A2(n_387),
.B1(n_555),
.B2(n_544),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_586),
.A2(n_498),
.B1(n_393),
.B2(n_378),
.Y(n_626)
);

AOI222xp33_ASAP7_75t_L g627 ( 
.A1(n_578),
.A2(n_362),
.B1(n_417),
.B2(n_499),
.C1(n_363),
.C2(n_376),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_586),
.A2(n_547),
.B1(n_544),
.B2(n_508),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_575),
.B(n_539),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_604),
.A2(n_387),
.B1(n_503),
.B2(n_500),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_591),
.A2(n_597),
.B1(n_582),
.B2(n_606),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_591),
.A2(n_597),
.B1(n_598),
.B2(n_571),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_608),
.A2(n_595),
.B(n_602),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_572),
.A2(n_503),
.B1(n_500),
.B2(n_485),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_SL g635 ( 
.A1(n_593),
.A2(n_503),
.B1(n_539),
.B2(n_477),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_588),
.A2(n_503),
.B1(n_500),
.B2(n_477),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_598),
.A2(n_468),
.B1(n_474),
.B2(n_476),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_588),
.B(n_508),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_592),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_583),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_576),
.A2(n_508),
.B1(n_363),
.B2(n_376),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_603),
.B(n_508),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_573),
.B(n_490),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_590),
.A2(n_363),
.B1(n_376),
.B2(n_490),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_584),
.A2(n_474),
.B1(n_468),
.B2(n_476),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_609),
.A2(n_485),
.B1(n_490),
.B2(n_486),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_579),
.A2(n_486),
.B1(n_484),
.B2(n_483),
.Y(n_647)
);

OA211x2_ASAP7_75t_L g648 ( 
.A1(n_611),
.A2(n_610),
.B(n_609),
.C(n_599),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_618),
.B(n_587),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_632),
.A2(n_610),
.B1(n_601),
.B2(n_593),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_622),
.B(n_605),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_616),
.A2(n_574),
.B(n_596),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_622),
.B(n_589),
.Y(n_653)
);

OA21x2_ASAP7_75t_L g654 ( 
.A1(n_640),
.A2(n_359),
.B(n_577),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_624),
.A2(n_594),
.B(n_593),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_612),
.B(n_600),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_SL g657 ( 
.A(n_639),
.B(n_594),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_631),
.B(n_594),
.C(n_486),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_614),
.B(n_620),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_SL g660 ( 
.A1(n_613),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.C(n_49),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_612),
.B(n_594),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_615),
.B(n_483),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_SL g663 ( 
.A1(n_619),
.A2(n_486),
.B(n_484),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_615),
.B(n_483),
.Y(n_664)
);

OAI221xp5_ASAP7_75t_L g665 ( 
.A1(n_634),
.A2(n_486),
.B1(n_484),
.B2(n_483),
.C(n_415),
.Y(n_665)
);

AOI221xp5_ASAP7_75t_L g666 ( 
.A1(n_633),
.A2(n_486),
.B1(n_484),
.B2(n_483),
.C(n_233),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_640),
.B(n_484),
.Y(n_667)
);

OA21x2_ASAP7_75t_L g668 ( 
.A1(n_645),
.A2(n_359),
.B(n_484),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_629),
.B(n_50),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_627),
.B(n_233),
.C(n_225),
.Y(n_670)
);

OAI211xp5_ASAP7_75t_L g671 ( 
.A1(n_633),
.A2(n_233),
.B(n_225),
.C(n_57),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_643),
.B(n_52),
.Y(n_672)
);

OAI221xp5_ASAP7_75t_L g673 ( 
.A1(n_617),
.A2(n_473),
.B1(n_233),
.B2(n_60),
.C(n_61),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_639),
.B(n_233),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_671),
.B(n_630),
.C(n_625),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_666),
.B(n_628),
.C(n_621),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_651),
.B(n_638),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_649),
.B(n_642),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_652),
.B(n_641),
.C(n_644),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_648),
.A2(n_637),
.B1(n_626),
.B2(n_623),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g681 ( 
.A(n_656),
.B(n_636),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_653),
.Y(n_682)
);

AOI211xp5_ASAP7_75t_L g683 ( 
.A1(n_660),
.A2(n_655),
.B(n_659),
.C(n_650),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_661),
.B(n_635),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_662),
.B(n_647),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_659),
.A2(n_646),
.B1(n_233),
.B2(n_62),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_658),
.B(n_233),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_664),
.B(n_54),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_667),
.B(n_58),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_668),
.B(n_64),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_657),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_668),
.B(n_70),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_682),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_677),
.Y(n_694)
);

XOR2xp5_ASAP7_75t_L g695 ( 
.A(n_681),
.B(n_669),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_677),
.Y(n_696)
);

XOR2x2_ASAP7_75t_L g697 ( 
.A(n_683),
.B(n_672),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_678),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_691),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_684),
.Y(n_700)
);

XNOR2xp5_ASAP7_75t_L g701 ( 
.A(n_684),
.B(n_670),
.Y(n_701)
);

XNOR2xp5_ASAP7_75t_L g702 ( 
.A(n_679),
.B(n_685),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_685),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_693),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_693),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_703),
.Y(n_706)
);

XOR2x2_ASAP7_75t_L g707 ( 
.A(n_697),
.B(n_675),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_694),
.Y(n_708)
);

XNOR2x1_ASAP7_75t_L g709 ( 
.A(n_707),
.B(n_702),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_704),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_705),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_707),
.A2(n_700),
.B1(n_701),
.B2(n_680),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_711),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_711),
.Y(n_715)
);

AOI322xp5_ASAP7_75t_L g716 ( 
.A1(n_713),
.A2(n_700),
.A3(n_699),
.B1(n_686),
.B2(n_696),
.C1(n_706),
.C2(n_708),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_710),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_714),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_715),
.Y(n_719)
);

NAND4xp25_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_709),
.C(n_712),
.D(n_676),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_719),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_718),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_720),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_719),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_723),
.A2(n_717),
.B1(n_695),
.B2(n_698),
.Y(n_725)
);

AOI221xp5_ASAP7_75t_L g726 ( 
.A1(n_723),
.A2(n_692),
.B1(n_673),
.B2(n_687),
.C(n_663),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_724),
.A2(n_674),
.B1(n_692),
.B2(n_687),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_722),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_721),
.B(n_690),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_722),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_723),
.A2(n_688),
.B1(n_690),
.B2(n_689),
.Y(n_731)
);

AOI221xp5_ASAP7_75t_L g732 ( 
.A1(n_723),
.A2(n_665),
.B1(n_72),
.B2(n_74),
.C(n_75),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_728),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_730),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_729),
.B(n_71),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_725),
.A2(n_668),
.B1(n_654),
.B2(n_79),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_732),
.A2(n_654),
.B1(n_78),
.B2(n_81),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_726),
.B(n_654),
.C(n_83),
.Y(n_738)
);

NOR2x1_ASAP7_75t_L g739 ( 
.A(n_731),
.B(n_77),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_727),
.Y(n_740)
);

AND5x1_ASAP7_75t_L g741 ( 
.A(n_737),
.B(n_145),
.C(n_87),
.D(n_88),
.E(n_89),
.Y(n_741)
);

NAND4xp25_ASAP7_75t_L g742 ( 
.A(n_733),
.B(n_85),
.C(n_90),
.D(n_91),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_734),
.B(n_92),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_738),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_740),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_739),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_736),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_745),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_743),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_747),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_744),
.A2(n_735),
.B1(n_104),
.B2(n_105),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_742),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_746),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_750),
.A2(n_748),
.B1(n_752),
.B2(n_753),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_753),
.A2(n_741),
.B1(n_107),
.B2(n_109),
.Y(n_755)
);

OAI22x1_ASAP7_75t_L g756 ( 
.A1(n_749),
.A2(n_103),
.B1(n_111),
.B2(n_114),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_751),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_757)
);

OA22x2_ASAP7_75t_L g758 ( 
.A1(n_750),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_750),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_759),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_754),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_758),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_756),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_761),
.A2(n_755),
.B1(n_757),
.B2(n_127),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_763),
.A2(n_123),
.B1(n_125),
.B2(n_129),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_SL g767 ( 
.A1(n_766),
.A2(n_762),
.B1(n_760),
.B2(n_765),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_767),
.Y(n_768)
);

AOI221x1_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.C(n_135),
.Y(n_769)
);

AOI211xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_136),
.B(n_139),
.C(n_141),
.Y(n_770)
);


endmodule