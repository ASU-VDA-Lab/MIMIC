module fake_jpeg_11421_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_3),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_5),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_0),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_18),
.B1(n_17),
.B2(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_32),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.B1(n_34),
.B2(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_43),
.B1(n_35),
.B2(n_21),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_31),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_51),
.C(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_16),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_32),
.B(n_16),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_57),
.C(n_50),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_44),
.B1(n_17),
.B2(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_17),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_46),
.C(n_48),
.Y(n_59)
);

AOI31xp67_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_62),
.A3(n_58),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_11),
.Y(n_64)
);

AOI221xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_52),
.B1(n_53),
.B2(n_50),
.C(n_12),
.Y(n_63)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_15),
.A3(n_13),
.B1(n_4),
.B2(n_5),
.C1(n_1),
.C2(n_2),
.Y(n_68)
);

OAI22x1_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_12),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_66),
.C(n_1),
.Y(n_69)
);

AOI221xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_68),
.B1(n_14),
.B2(n_13),
.C(n_35),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_5),
.C(n_13),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.C(n_35),
.Y(n_72)
);


endmodule