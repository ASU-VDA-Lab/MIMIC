module fake_jpeg_22785_n_258 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_14),
.B(n_20),
.C(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_21),
.B1(n_20),
.B2(n_27),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_50),
.B1(n_18),
.B2(n_22),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_16),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_51),
.Y(n_65)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_21),
.B1(n_16),
.B2(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_14),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_25),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_76),
.B1(n_46),
.B2(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_64),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_19),
.C(n_34),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_77),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_16),
.B(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_68),
.B1(n_78),
.B2(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_21),
.B1(n_22),
.B2(n_14),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_50),
.B1(n_28),
.B2(n_26),
.Y(n_93)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_71),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_18),
.B1(n_28),
.B2(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_75),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_14),
.B1(n_18),
.B2(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_82),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_54),
.B1(n_39),
.B2(n_47),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_59),
.B1(n_78),
.B2(n_67),
.Y(n_112)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_84),
.B(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_23),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_70),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_51),
.B1(n_44),
.B2(n_49),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_99),
.B1(n_69),
.B2(n_7),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_100),
.B1(n_23),
.B2(n_75),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_58),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_57),
.B1(n_44),
.B2(n_26),
.Y(n_100)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_66),
.B(n_74),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_106),
.B(n_108),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_105),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_62),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_66),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_66),
.B(n_59),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_109),
.A2(n_83),
.B1(n_84),
.B2(n_82),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_71),
.B1(n_57),
.B2(n_75),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_115),
.B1(n_120),
.B2(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_69),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_0),
.B(n_2),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_86),
.C(n_100),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_100),
.B(n_93),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_102),
.B(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_94),
.B1(n_93),
.B2(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_94),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_144),
.B(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_94),
.B1(n_93),
.B2(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_93),
.B1(n_90),
.B2(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_135),
.Y(n_150)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_140),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_83),
.B1(n_82),
.B2(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_8),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_8),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_2),
.B(n_3),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_103),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_148),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_105),
.C(n_118),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_129),
.C(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_103),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_114),
.Y(n_152)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_141),
.B1(n_125),
.B2(n_144),
.C(n_120),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_161),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_126),
.B(n_125),
.Y(n_181)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_161),
.B(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_150),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_175),
.B(n_181),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_140),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_184),
.C(n_164),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_126),
.B1(n_131),
.B2(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_186),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_141),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_182),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_155),
.B(n_159),
.C(n_156),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_125),
.B1(n_109),
.B2(n_106),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_160),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_106),
.C(n_110),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_121),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_168),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_193),
.C(n_199),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_152),
.C(n_157),
.Y(n_193)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_179),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_162),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_149),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_149),
.C(n_151),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_153),
.C(n_148),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_145),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_210),
.C(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_185),
.B1(n_181),
.B2(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_174),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_153),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_159),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_215),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_154),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_182),
.B(n_121),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_195),
.B(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_9),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_188),
.C(n_198),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_187),
.C(n_202),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_211),
.C(n_187),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_202),
.B(n_9),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_222),
.C(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_210),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_13),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_8),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_234),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_235),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_238),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_223),
.B(n_7),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_6),
.C(n_11),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_10),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_227),
.C(n_10),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_243),
.B(n_244),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_6),
.B(n_12),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_SL g251 ( 
.A1(n_246),
.A2(n_247),
.B(n_249),
.C(n_239),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_232),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_251),
.A2(n_252),
.B(n_13),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_12),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_13),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_255),
.B(n_2),
.C(n_4),
.D(n_5),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_4),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_5),
.Y(n_258)
);


endmodule