module fake_jpeg_23533_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

HAxp5_ASAP7_75t_SL g38 ( 
.A(n_19),
.B(n_0),
.CON(n_38),
.SN(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_28),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_39),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_27),
.B1(n_18),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_55),
.B1(n_57),
.B2(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_27),
.B1(n_18),
.B2(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_27),
.B1(n_21),
.B2(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_60),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_66),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_21),
.B1(n_36),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_71),
.B1(n_78),
.B2(n_30),
.Y(n_105)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_21),
.B1(n_26),
.B2(n_16),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_83),
.B1(n_43),
.B2(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_73),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_16),
.A3(n_40),
.B1(n_32),
.B2(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_1),
.B(n_2),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_22),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_68),
.B1(n_66),
.B2(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_28),
.B1(n_22),
.B2(n_30),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_15),
.B(n_75),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_104),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_96),
.B1(n_15),
.B2(n_40),
.Y(n_130)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_102),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_43),
.B1(n_46),
.B2(n_45),
.Y(n_99)
);

OAI22x1_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_100),
.B1(n_22),
.B2(n_70),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_46),
.B1(n_13),
.B2(n_8),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_34),
.C(n_33),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_40),
.C(n_61),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_40),
.B1(n_15),
.B2(n_33),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_72),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_113),
.B(n_123),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_81),
.B(n_77),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_112),
.B(n_120),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_115),
.B1(n_114),
.B2(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_122),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_79),
.B(n_78),
.Y(n_112)
);

OR2x4_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_130),
.B1(n_94),
.B2(n_90),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_88),
.C(n_86),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_40),
.Y(n_132)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_124),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_25),
.B(n_19),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_14),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_2),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_10),
.Y(n_125)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_3),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_126),
.B(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_102),
.B1(n_95),
.B2(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_136),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_110),
.B1(n_107),
.B2(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_37),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_142),
.C(n_151),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_37),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_37),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_128),
.B1(n_124),
.B2(n_119),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_15),
.B(n_4),
.C(n_5),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_146),
.B(n_111),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_85),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_34),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_34),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_153),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_148),
.B(n_145),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_133),
.C(n_136),
.Y(n_177)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_174),
.B1(n_140),
.B2(n_145),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_108),
.C(n_110),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_167),
.C(n_170),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_168),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_107),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_159),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_107),
.C(n_119),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_123),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_90),
.C(n_122),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_127),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_175),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_127),
.B1(n_125),
.B2(n_94),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_34),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_186),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_142),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_191),
.C(n_157),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_190),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_132),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_150),
.B(n_149),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_118),
.B(n_175),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_167),
.B(n_162),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_185),
.B(n_191),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_193),
.C(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_157),
.B1(n_147),
.B2(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_164),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_213),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_212),
.B1(n_12),
.B2(n_11),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_194),
.A2(n_173),
.B1(n_168),
.B2(n_70),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_193),
.B1(n_207),
.B2(n_198),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_216),
.B(n_199),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_223),
.C(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_209),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_222),
.B1(n_63),
.B2(n_4),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_178),
.B1(n_61),
.B2(n_42),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_178),
.C(n_69),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_226),
.B1(n_219),
.B2(n_227),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_230),
.B1(n_235),
.B2(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_234),
.C(n_238),
.Y(n_244)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_199),
.C(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_10),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_205),
.B1(n_200),
.B2(n_206),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_63),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_239),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_69),
.B1(n_4),
.B2(n_5),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_63),
.C(n_4),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_222),
.B1(n_225),
.B2(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_223),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_19),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_238),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_248),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_247),
.B(n_11),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_25),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_11),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_233),
.B(n_234),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_244),
.B(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_251),
.B(n_241),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_229),
.B(n_12),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_3),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_19),
.Y(n_255)
);

A2O1A1O1Ixp25_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_3),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_254),
.B1(n_256),
.B2(n_6),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_263),
.Y(n_265)
);

OAI311xp33_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_257),
.A3(n_7),
.B1(n_3),
.C1(n_25),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_266),
.A2(n_262),
.B1(n_7),
.B2(n_25),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_265),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_19),
.B(n_25),
.Y(n_269)
);


endmodule