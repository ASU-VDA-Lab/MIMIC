module real_aes_8483_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_1), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_2), .A2(n_145), .B(n_148), .C(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_3), .A2(n_173), .B(n_174), .Y(n_172) );
INVx1_ASAP7_75t_L g501 ( .A(n_4), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_5), .B(n_184), .Y(n_183) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_6), .A2(n_173), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g145 ( .A(n_7), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g248 ( .A(n_8), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_9), .B(n_41), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_9), .B(n_41), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_10), .A2(n_272), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_11), .B(n_157), .Y(n_225) );
INVx1_ASAP7_75t_L g483 ( .A(n_12), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_13), .B(n_178), .Y(n_534) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
INVx1_ASAP7_75t_L g546 ( .A(n_15), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_16), .A2(n_192), .B(n_233), .C(n_235), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_17), .B(n_184), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_18), .B(n_472), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_19), .B(n_173), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_20), .B(n_280), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_21), .A2(n_178), .B(n_209), .C(n_212), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_22), .B(n_184), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_23), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_24), .A2(n_211), .B(n_235), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_25), .B(n_157), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_26), .Y(n_139) );
INVx1_ASAP7_75t_L g190 ( .A(n_27), .Y(n_190) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_28), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_29), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_30), .B(n_157), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_31), .Y(n_453) );
INVx1_ASAP7_75t_L g277 ( .A(n_32), .Y(n_277) );
INVx1_ASAP7_75t_L g491 ( .A(n_33), .Y(n_491) );
INVx2_ASAP7_75t_L g143 ( .A(n_34), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_35), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_36), .A2(n_178), .B(n_179), .C(n_181), .Y(n_177) );
INVxp67_ASAP7_75t_L g278 ( .A(n_37), .Y(n_278) );
CKINVDCx14_ASAP7_75t_R g175 ( .A(n_38), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_39), .A2(n_148), .B(n_189), .C(n_196), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_40), .A2(n_145), .B(n_148), .C(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g490 ( .A(n_42), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_43), .A2(n_49), .B1(n_445), .B2(n_446), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_43), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_44), .A2(n_62), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_44), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_45), .A2(n_159), .B(n_246), .C(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_46), .B(n_157), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_47), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_48), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_49), .Y(n_445) );
INVx1_ASAP7_75t_L g207 ( .A(n_50), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_51), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_52), .B(n_173), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_53), .A2(n_148), .B1(n_212), .B2(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_54), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_55), .Y(n_498) );
CKINVDCx14_ASAP7_75t_R g244 ( .A(n_56), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_57), .A2(n_181), .B(n_246), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_58), .Y(n_526) );
INVx1_ASAP7_75t_L g480 ( .A(n_59), .Y(n_480) );
INVx1_ASAP7_75t_L g146 ( .A(n_60), .Y(n_146) );
INVx1_ASAP7_75t_L g136 ( .A(n_61), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_62), .Y(n_744) );
INVx1_ASAP7_75t_SL g180 ( .A(n_63), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_64), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_65), .B(n_184), .Y(n_214) );
INVx1_ASAP7_75t_L g152 ( .A(n_66), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_SL g471 ( .A1(n_67), .A2(n_181), .B(n_472), .C(n_473), .Y(n_471) );
INVxp67_ASAP7_75t_L g474 ( .A(n_68), .Y(n_474) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_70), .A2(n_173), .B(n_243), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_71), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_72), .A2(n_173), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_73), .Y(n_494) );
INVx1_ASAP7_75t_L g520 ( .A(n_74), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_75), .A2(n_272), .B(n_273), .Y(n_271) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_76), .Y(n_187) );
INVx1_ASAP7_75t_L g231 ( .A(n_77), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_78), .A2(n_145), .B(n_148), .C(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_79), .A2(n_173), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g234 ( .A(n_80), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_81), .B(n_191), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_82), .A2(n_102), .B1(n_115), .B2(n_754), .Y(n_101) );
INVx2_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
INVx1_ASAP7_75t_L g224 ( .A(n_84), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_85), .B(n_472), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_86), .A2(n_145), .B(n_148), .C(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
OR2x2_ASAP7_75t_L g448 ( .A(n_87), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g741 ( .A(n_87), .B(n_450), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_88), .A2(n_148), .B(n_151), .C(n_161), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_89), .B(n_166), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_90), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_91), .A2(n_145), .B(n_148), .C(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_92), .Y(n_538) );
INVx1_ASAP7_75t_L g470 ( .A(n_93), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_94), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_95), .B(n_191), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_96), .B(n_132), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_97), .B(n_132), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g210 ( .A(n_99), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_100), .A2(n_173), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g754 ( .A(n_104), .Y(n_754) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g450 ( .A(n_110), .B(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g458 ( .A(n_111), .B(n_450), .Y(n_458) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_111), .B(n_449), .Y(n_750) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_454), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g753 ( .A(n_119), .Y(n_753) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_447), .B(n_452), .Y(n_121) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_444), .Y(n_122) );
INVx3_ASAP7_75t_L g742 ( .A(n_123), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_123), .A2(n_457), .B1(n_740), .B2(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_399), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_336), .C(n_370), .D(n_386), .Y(n_124) );
NAND4xp25_ASAP7_75t_SL g125 ( .A(n_126), .B(n_262), .C(n_300), .D(n_316), .Y(n_125) );
AOI222xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_199), .B1(n_237), .B2(n_250), .C1(n_255), .C2(n_261), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI31xp33_ASAP7_75t_L g432 ( .A1(n_128), .A2(n_433), .A3(n_434), .B(n_436), .Y(n_432) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_167), .Y(n_128) );
AND2x2_ASAP7_75t_L g407 ( .A(n_129), .B(n_169), .Y(n_407) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_SL g254 ( .A(n_130), .Y(n_254) );
AND2x2_ASAP7_75t_L g261 ( .A(n_130), .B(n_185), .Y(n_261) );
AND2x2_ASAP7_75t_L g321 ( .A(n_130), .B(n_170), .Y(n_321) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_163), .Y(n_130) );
INVx3_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_131), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_131), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_SL g516 ( .A(n_131), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_132), .A2(n_468), .B(n_475), .Y(n_467) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g270 ( .A(n_133), .Y(n_270) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_134), .B(n_135), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_147), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_140), .A2(n_166), .B(n_187), .C(n_188), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_140), .A2(n_221), .B(n_222), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_140), .A2(n_162), .B1(n_488), .B2(n_492), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_140), .A2(n_498), .B(n_499), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_140), .A2(n_520), .B(n_521), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
AND2x4_ASAP7_75t_L g173 ( .A(n_141), .B(n_145), .Y(n_173) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx1_ASAP7_75t_L g213 ( .A(n_143), .Y(n_213) );
INVx1_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
INVx3_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
INVx1_ASAP7_75t_L g472 ( .A(n_144), .Y(n_472) );
INVx4_ASAP7_75t_SL g162 ( .A(n_145), .Y(n_162) );
BUFx3_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
INVx5_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx3_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_156), .C(n_158), .Y(n_151) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_153), .A2(n_158), .B(n_224), .C(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_154), .A2(n_155), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
INVx4_ASAP7_75t_L g178 ( .A(n_157), .Y(n_178) );
INVx2_ASAP7_75t_L g246 ( .A(n_157), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_158), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_158), .A2(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g235 ( .A(n_160), .Y(n_235) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_162), .A2(n_175), .B(n_176), .C(n_177), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g206 ( .A1(n_162), .A2(n_176), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_SL g230 ( .A1(n_162), .A2(n_176), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g243 ( .A1(n_162), .A2(n_176), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g273 ( .A1(n_162), .A2(n_176), .B(n_274), .C(n_275), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_162), .A2(n_176), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_162), .A2(n_176), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_162), .A2(n_176), .B(n_543), .C(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx1_ASAP7_75t_L g280 ( .A(n_165), .Y(n_280) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_165), .A2(n_530), .B(n_537), .Y(n_529) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g219 ( .A(n_166), .Y(n_219) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_166), .A2(n_242), .B(n_249), .Y(n_241) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_166), .A2(n_541), .B(n_547), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_167), .B(n_351), .Y(n_350) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_168), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_168), .B(n_265), .Y(n_311) );
AND2x2_ASAP7_75t_L g404 ( .A(n_168), .B(n_344), .Y(n_404) );
OAI321xp33_ASAP7_75t_L g438 ( .A1(n_168), .A2(n_254), .A3(n_411), .B1(n_439), .B2(n_441), .C(n_442), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g442 ( .A(n_168), .B(n_240), .C(n_351), .D(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_185), .Y(n_168) );
AND2x2_ASAP7_75t_L g306 ( .A(n_169), .B(n_252), .Y(n_306) );
AND2x2_ASAP7_75t_L g325 ( .A(n_169), .B(n_254), .Y(n_325) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g253 ( .A(n_170), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g281 ( .A(n_170), .B(n_185), .Y(n_281) );
AND2x2_ASAP7_75t_L g367 ( .A(n_170), .B(n_252), .Y(n_367) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_183), .Y(n_170) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_205), .B(n_214), .Y(n_204) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_171), .A2(n_229), .B(n_236), .Y(n_228) );
BUFx2_ASAP7_75t_L g272 ( .A(n_173), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_178), .B(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_182), .Y(n_535) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_184), .A2(n_478), .B(n_484), .Y(n_477) );
INVx3_ASAP7_75t_SL g252 ( .A(n_185), .Y(n_252) );
AND2x2_ASAP7_75t_L g299 ( .A(n_185), .B(n_286), .Y(n_299) );
OR2x2_ASAP7_75t_L g332 ( .A(n_185), .B(n_254), .Y(n_332) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_185), .Y(n_339) );
AND2x2_ASAP7_75t_L g368 ( .A(n_185), .B(n_253), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_185), .B(n_341), .Y(n_383) );
AND2x2_ASAP7_75t_L g415 ( .A(n_185), .B(n_407), .Y(n_415) );
AND2x2_ASAP7_75t_L g424 ( .A(n_185), .B(n_266), .Y(n_424) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_193), .C(n_194), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_191), .A2(n_211), .B1(n_277), .B2(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_191), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
INVx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_192), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_192), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_192), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_195), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_215), .Y(n_200) );
INVx1_ASAP7_75t_SL g392 ( .A(n_201), .Y(n_392) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g257 ( .A(n_202), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g239 ( .A(n_203), .B(n_217), .Y(n_239) );
AND2x2_ASAP7_75t_L g328 ( .A(n_203), .B(n_241), .Y(n_328) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g298 ( .A(n_204), .B(n_228), .Y(n_298) );
OR2x2_ASAP7_75t_L g309 ( .A(n_204), .B(n_241), .Y(n_309) );
AND2x2_ASAP7_75t_L g335 ( .A(n_204), .B(n_241), .Y(n_335) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_204), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_211), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_211), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g503 ( .A(n_212), .Y(n_503) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_215), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_215), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g308 ( .A(n_216), .B(n_309), .Y(n_308) );
AOI322xp5_ASAP7_75t_L g394 ( .A1(n_216), .A2(n_298), .A3(n_304), .B1(n_335), .B2(n_385), .C1(n_395), .C2(n_397), .Y(n_394) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_228), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_217), .B(n_240), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_217), .B(n_241), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_217), .B(n_258), .Y(n_315) );
AND2x2_ASAP7_75t_L g369 ( .A(n_217), .B(n_335), .Y(n_369) );
INVx1_ASAP7_75t_L g373 ( .A(n_217), .Y(n_373) );
AND2x2_ASAP7_75t_L g385 ( .A(n_217), .B(n_228), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_217), .B(n_257), .Y(n_417) );
INVx4_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g282 ( .A(n_218), .B(n_228), .Y(n_282) );
BUFx3_ASAP7_75t_L g296 ( .A(n_218), .Y(n_296) );
AND3x2_ASAP7_75t_L g378 ( .A(n_218), .B(n_358), .C(n_379), .Y(n_378) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_219), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_219), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_219), .B(n_538), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g238 ( .A(n_228), .B(n_239), .C(n_240), .Y(n_238) );
INVx1_ASAP7_75t_SL g258 ( .A(n_228), .Y(n_258) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_228), .Y(n_363) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g357 ( .A(n_239), .B(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g364 ( .A(n_239), .Y(n_364) );
AND2x2_ASAP7_75t_L g402 ( .A(n_240), .B(n_380), .Y(n_402) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx3_ASAP7_75t_L g283 ( .A(n_241), .Y(n_283) );
AND2x2_ASAP7_75t_L g358 ( .A(n_241), .B(n_258), .Y(n_358) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
OR2x2_ASAP7_75t_L g302 ( .A(n_252), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g421 ( .A(n_252), .B(n_321), .Y(n_421) );
AND2x2_ASAP7_75t_L g435 ( .A(n_252), .B(n_254), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_253), .B(n_266), .Y(n_376) );
AND2x2_ASAP7_75t_L g423 ( .A(n_253), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g286 ( .A(n_254), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g303 ( .A(n_254), .B(n_266), .Y(n_303) );
INVx1_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
AND2x2_ASAP7_75t_L g344 ( .A(n_254), .B(n_266), .Y(n_344) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_256), .A2(n_387), .B1(n_391), .B2(n_393), .C(n_394), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_257), .B(n_259), .Y(n_256) );
AND2x2_ASAP7_75t_L g290 ( .A(n_257), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_260), .B(n_297), .Y(n_440) );
AOI322xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_282), .A3(n_283), .B1(n_284), .B2(n_290), .C1(n_292), .C2(n_299), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_281), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_265), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_265), .B(n_331), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_265), .A2(n_281), .B(n_355), .C(n_356), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_265), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_265), .B(n_325), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_265), .B(n_407), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_265), .B(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_266), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_266), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g396 ( .A(n_266), .B(n_283), .Y(n_396) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_271), .B(n_279), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_268), .A2(n_288), .B(n_289), .Y(n_287) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_268), .A2(n_519), .B(n_525), .Y(n_518) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI21xp5_ASAP7_75t_SL g510 ( .A1(n_269), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_270), .A2(n_487), .B(n_493), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_270), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_270), .A2(n_497), .B(n_504), .Y(n_496) );
INVx1_ASAP7_75t_L g288 ( .A(n_271), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_279), .Y(n_289) );
INVx1_ASAP7_75t_L g371 ( .A(n_281), .Y(n_371) );
OAI31xp33_ASAP7_75t_L g381 ( .A1(n_281), .A2(n_306), .A3(n_382), .B(n_384), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_281), .B(n_287), .Y(n_433) );
INVx1_ASAP7_75t_SL g294 ( .A(n_282), .Y(n_294) );
AND2x2_ASAP7_75t_L g327 ( .A(n_282), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g408 ( .A(n_282), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g293 ( .A(n_283), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g318 ( .A(n_283), .Y(n_318) );
AND2x2_ASAP7_75t_L g345 ( .A(n_283), .B(n_298), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_283), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g437 ( .A(n_283), .B(n_385), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_285), .B(n_355), .Y(n_428) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g324 ( .A(n_287), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g342 ( .A(n_287), .Y(n_342) );
NAND2xp33_ASAP7_75t_SL g292 ( .A(n_293), .B(n_295), .Y(n_292) );
OAI211xp5_ASAP7_75t_SL g336 ( .A1(n_294), .A2(n_337), .B(n_343), .C(n_359), .Y(n_336) );
OR2x2_ASAP7_75t_L g411 ( .A(n_294), .B(n_392), .Y(n_411) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_296), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_296), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g317 ( .A(n_298), .B(n_318), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B(n_307), .C(n_310), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g351 ( .A(n_303), .Y(n_351) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_306), .B(n_344), .Y(n_349) );
INVx1_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g314 ( .A(n_309), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g347 ( .A(n_309), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g409 ( .A(n_309), .Y(n_409) );
AOI21xp33_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_312), .B(n_314), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_312), .A2(n_323), .B(n_326), .Y(n_322) );
AOI211xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B(n_322), .C(n_329), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_317), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_320), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_SL g333 ( .A(n_321), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_323), .A2(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_328), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g353 ( .A(n_328), .Y(n_353) );
AOI21xp33_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_333), .B(n_334), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g384 ( .A(n_335), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_341), .B(n_367), .Y(n_393) );
AND2x2_ASAP7_75t_L g406 ( .A(n_341), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g420 ( .A(n_341), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g430 ( .A(n_341), .B(n_368), .Y(n_430) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B(n_346), .C(n_354), .Y(n_343) );
INVx1_ASAP7_75t_L g390 ( .A(n_344), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B1(n_350), .B2(n_352), .Y(n_346) );
OR2x2_ASAP7_75t_L g352 ( .A(n_348), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_348), .B(n_409), .Y(n_431) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g425 ( .A(n_358), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_365), .B1(n_368), .B2(n_369), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g443 ( .A(n_363), .Y(n_443) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g389 ( .A(n_367), .Y(n_389) );
OAI211xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_372), .B(n_374), .C(n_381), .Y(n_370) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_389), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR5xp2_ASAP7_75t_L g399 ( .A(n_400), .B(n_418), .C(n_426), .D(n_432), .E(n_438), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_403), .B(n_405), .C(n_412), .Y(n_400) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_410), .Y(n_405) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_415), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B(n_425), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g441 ( .A(n_421), .Y(n_441) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2xp33_ASAP7_75t_SL g452 ( .A(n_448), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI21xp5_ASAP7_75t_SL g454 ( .A1(n_452), .A2(n_455), .B(n_752), .Y(n_454) );
OAI222xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_743), .B1(n_746), .B2(n_748), .C1(n_749), .C2(n_751), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_740), .B2(n_742), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g747 ( .A(n_459), .Y(n_747) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND4x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_658), .C(n_705), .D(n_725), .Y(n_460) );
NOR3xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_588), .C(n_613), .Y(n_461) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_506), .B(n_548), .C(n_578), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_485), .Y(n_464) );
INVx3_ASAP7_75t_SL g630 ( .A(n_465), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_465), .B(n_561), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_465), .B(n_495), .Y(n_711) );
AND2x2_ASAP7_75t_L g734 ( .A(n_465), .B(n_600), .Y(n_734) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g552 ( .A(n_467), .B(n_477), .Y(n_552) );
INVx3_ASAP7_75t_L g565 ( .A(n_467), .Y(n_565) );
AND2x2_ASAP7_75t_L g570 ( .A(n_467), .B(n_476), .Y(n_570) );
OR2x2_ASAP7_75t_L g621 ( .A(n_467), .B(n_562), .Y(n_621) );
BUFx2_ASAP7_75t_L g641 ( .A(n_467), .Y(n_641) );
AND2x2_ASAP7_75t_L g651 ( .A(n_467), .B(n_562), .Y(n_651) );
AND2x2_ASAP7_75t_L g657 ( .A(n_467), .B(n_486), .Y(n_657) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_477), .B(n_562), .Y(n_576) );
INVx2_ASAP7_75t_L g586 ( .A(n_477), .Y(n_586) );
AND2x2_ASAP7_75t_L g599 ( .A(n_477), .B(n_565), .Y(n_599) );
OR2x2_ASAP7_75t_L g610 ( .A(n_477), .B(n_562), .Y(n_610) );
AND2x2_ASAP7_75t_SL g656 ( .A(n_477), .B(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g668 ( .A(n_477), .Y(n_668) );
AND2x2_ASAP7_75t_L g714 ( .A(n_477), .B(n_486), .Y(n_714) );
INVx3_ASAP7_75t_SL g587 ( .A(n_485), .Y(n_587) );
OR2x2_ASAP7_75t_L g640 ( .A(n_485), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
INVx3_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
AND2x2_ASAP7_75t_L g629 ( .A(n_486), .B(n_496), .Y(n_629) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_486), .Y(n_697) );
AOI33xp33_ASAP7_75t_L g701 ( .A1(n_486), .A2(n_630), .A3(n_637), .B1(n_646), .B2(n_702), .B3(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g550 ( .A(n_495), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_495), .B(n_565), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_495), .B(n_625), .C(n_627), .Y(n_624) );
AND2x2_ASAP7_75t_L g650 ( .A(n_495), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_495), .B(n_657), .Y(n_660) );
AND2x2_ASAP7_75t_L g713 ( .A(n_495), .B(n_714), .Y(n_713) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g569 ( .A(n_496), .Y(n_569) );
OR2x2_ASAP7_75t_L g663 ( .A(n_496), .B(n_562), .Y(n_663) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_527), .Y(n_506) );
AOI32xp33_ASAP7_75t_L g614 ( .A1(n_507), .A2(n_615), .A3(n_617), .B1(n_619), .B2(n_622), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g687 ( .A(n_507), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g717 ( .A(n_507), .Y(n_717) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g649 ( .A(n_508), .B(n_633), .Y(n_649) );
AND2x2_ASAP7_75t_L g669 ( .A(n_508), .B(n_595), .Y(n_669) );
AND2x2_ASAP7_75t_L g737 ( .A(n_508), .B(n_655), .Y(n_737) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
INVx3_ASAP7_75t_L g558 ( .A(n_509), .Y(n_558) );
AND2x2_ASAP7_75t_L g572 ( .A(n_509), .B(n_556), .Y(n_572) );
OR2x2_ASAP7_75t_L g577 ( .A(n_509), .B(n_555), .Y(n_577) );
INVx1_ASAP7_75t_L g584 ( .A(n_509), .Y(n_584) );
AND2x2_ASAP7_75t_L g592 ( .A(n_509), .B(n_566), .Y(n_592) );
AND2x2_ASAP7_75t_L g594 ( .A(n_509), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_509), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g647 ( .A(n_509), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_509), .B(n_732), .Y(n_731) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .Y(n_509) );
INVx2_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
AND2x2_ASAP7_75t_L g602 ( .A(n_518), .B(n_528), .Y(n_602) );
AND2x2_ASAP7_75t_L g612 ( .A(n_518), .B(n_540), .Y(n_612) );
INVx2_ASAP7_75t_L g732 ( .A(n_527), .Y(n_732) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_528), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
AND2x2_ASAP7_75t_L g617 ( .A(n_528), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g633 ( .A(n_528), .B(n_596), .Y(n_633) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g581 ( .A(n_529), .Y(n_581) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g646 ( .A(n_529), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_529), .B(n_556), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g557 ( .A(n_539), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g618 ( .A(n_539), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_539), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g655 ( .A(n_539), .Y(n_655) );
INVx1_ASAP7_75t_L g688 ( .A(n_539), .Y(n_688) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g566 ( .A(n_540), .B(n_556), .Y(n_566) );
INVx1_ASAP7_75t_L g596 ( .A(n_540), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_553), .B1(n_559), .B2(n_566), .C(n_567), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_550), .B(n_570), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_550), .B(n_633), .Y(n_710) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_552), .B(n_600), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_552), .B(n_561), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_552), .B(n_575), .Y(n_704) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g626 ( .A(n_556), .Y(n_626) );
AND2x2_ASAP7_75t_L g601 ( .A(n_557), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g679 ( .A(n_557), .Y(n_679) );
AND2x2_ASAP7_75t_L g611 ( .A(n_558), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_558), .B(n_581), .Y(n_627) );
AND2x2_ASAP7_75t_L g691 ( .A(n_558), .B(n_617), .Y(n_691) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g600 ( .A(n_562), .B(n_569), .Y(n_600) );
AND2x2_ASAP7_75t_L g696 ( .A(n_563), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_565), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_566), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_566), .B(n_573), .Y(n_661) );
AND2x2_ASAP7_75t_L g681 ( .A(n_566), .B(n_581), .Y(n_681) );
AND2x2_ASAP7_75t_L g702 ( .A(n_566), .B(n_646), .Y(n_702) );
OAI32xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_571), .A3(n_573), .B1(n_574), .B2(n_577), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_SL g575 ( .A(n_569), .Y(n_575) );
NAND2x1_ASAP7_75t_L g616 ( .A(n_569), .B(n_599), .Y(n_616) );
OR2x2_ASAP7_75t_L g620 ( .A(n_569), .B(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_569), .B(n_668), .Y(n_721) );
INVx1_ASAP7_75t_L g589 ( .A(n_570), .Y(n_589) );
OAI221xp5_ASAP7_75t_SL g707 ( .A1(n_571), .A2(n_662), .B1(n_708), .B2(n_711), .C(n_712), .Y(n_707) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g579 ( .A(n_572), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g622 ( .A(n_572), .B(n_595), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_572), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g700 ( .A(n_572), .B(n_633), .Y(n_700) );
INVxp67_ASAP7_75t_L g636 ( .A(n_573), .Y(n_636) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g706 ( .A(n_575), .B(n_693), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_575), .B(n_656), .Y(n_729) );
INVx1_ASAP7_75t_L g604 ( .A(n_577), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_577), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g722 ( .A(n_577), .B(n_723), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_582), .B(n_585), .Y(n_578) );
AND2x2_ASAP7_75t_L g591 ( .A(n_580), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g675 ( .A(n_584), .B(n_595), .Y(n_675) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AND2x2_ASAP7_75t_L g693 ( .A(n_586), .B(n_651), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_586), .B(n_650), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_587), .B(n_599), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_593), .C(n_603), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_624), .B1(n_628), .B2(n_631), .C(n_634), .Y(n_623) );
AOI31xp33_ASAP7_75t_L g718 ( .A1(n_589), .A2(n_719), .A3(n_720), .B(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B1(n_599), .B2(n_601), .Y(n_593) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g719 ( .A(n_599), .Y(n_719) );
INVx1_ASAP7_75t_L g682 ( .A(n_600), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g725 ( .A1(n_602), .A2(n_726), .B(n_728), .C(n_730), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_607), .B2(n_611), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_608), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_610), .A2(n_644), .B1(n_663), .B2(n_699), .C(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g694 ( .A(n_611), .Y(n_694) );
INVx1_ASAP7_75t_L g648 ( .A(n_612), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g613 ( .A(n_614), .B(n_623), .C(n_638), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_615), .A2(n_665), .B(n_669), .Y(n_664) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_617), .B(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g724 ( .A(n_618), .Y(n_724) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g662 ( .A(n_625), .B(n_645), .Y(n_662) );
INVx1_ASAP7_75t_L g637 ( .A(n_626), .Y(n_637) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g635 ( .A(n_629), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_629), .B(n_667), .Y(n_666) );
NOR4xp25_ASAP7_75t_L g634 ( .A(n_630), .B(n_635), .C(n_636), .D(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_643), .B1(n_649), .B2(n_650), .C1(n_652), .C2(n_656), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g736 ( .A(n_640), .Y(n_736) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_652), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g712 ( .A1(n_657), .A2(n_713), .B(n_715), .Y(n_712) );
NOR4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_670), .C(n_683), .D(n_698), .Y(n_658) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_663), .C(n_664), .Y(n_659) );
INVx1_ASAP7_75t_L g739 ( .A(n_660), .Y(n_739) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_667), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
OAI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B1(n_676), .B2(n_677), .C1(n_680), .C2(n_682), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_675), .A2(n_706), .B(n_707), .C(n_718), .Y(n_705) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
OAI222xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_689), .B1(n_690), .B2(n_692), .C1(n_694), .C2(n_695), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_700), .A2(n_703), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI211xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_733), .B(n_735), .C(n_738), .Y(n_730) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g748 ( .A(n_743), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule