module fake_jpeg_20547_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx4_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_19),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_0),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_16),
.C(n_15),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_28),
.C(n_29),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_14),
.B1(n_7),
.B2(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_21),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_16),
.C(n_17),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_13),
.B(n_16),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_21),
.B(n_20),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_32),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_20),
.C(n_23),
.Y(n_37)
);

BUFx24_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_2),
.B(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_39),
.C(n_23),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.C(n_4),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_6),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_6),
.B(n_1),
.Y(n_46)
);


endmodule