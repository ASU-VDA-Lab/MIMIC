module fake_jpeg_29160_n_331 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx9p33_ASAP7_75t_R g99 ( 
.A(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_53),
.Y(n_71)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_45),
.Y(n_104)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_27),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_57),
.B1(n_23),
.B2(n_31),
.Y(n_88)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_22),
.A2(n_9),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_63),
.Y(n_76)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_61),
.B(n_26),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_28),
.Y(n_83)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_28),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_26),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_89),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_38),
.B1(n_35),
.B2(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_72),
.A2(n_77),
.B1(n_15),
.B2(n_36),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_75),
.B(n_87),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_38),
.B1(n_35),
.B2(n_18),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_37),
.B(n_34),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_78),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_40),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_81),
.B(n_85),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_87),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_40),
.B(n_31),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g87 ( 
.A(n_51),
.B(n_19),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_97),
.B1(n_27),
.B2(n_17),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_37),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_33),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_101),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_27),
.B1(n_23),
.B2(n_36),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_28),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_112),
.C(n_36),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_18),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_108),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_32),
.Y(n_108)
);

BUFx16f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx12_ASAP7_75t_R g111 ( 
.A(n_41),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_113),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_28),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_46),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_116),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g116 ( 
.A(n_66),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_48),
.B(n_28),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_19),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_124),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_93),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_139),
.B1(n_104),
.B2(n_118),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_30),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_160),
.Y(n_176)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

XOR2x1_ASAP7_75t_L g201 ( 
.A(n_136),
.B(n_141),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_36),
.B1(n_29),
.B2(n_27),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_154),
.B1(n_155),
.B2(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_164),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_78),
.A2(n_87),
.B(n_75),
.C(n_99),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_95),
.B(n_104),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_21),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_147),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_30),
.B1(n_21),
.B2(n_3),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_150),
.B1(n_86),
.B2(n_110),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_30),
.C(n_21),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_159),
.C(n_86),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_0),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_83),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_99),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_76),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_89),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_110),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_7),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_161),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_98),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_107),
.B(n_82),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_94),
.B(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_83),
.B(n_98),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_74),
.B(n_79),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_80),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_174),
.B1(n_186),
.B2(n_188),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_92),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_194),
.C(n_185),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_179),
.B(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_132),
.B(n_107),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_187),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_184),
.A2(n_192),
.B1(n_124),
.B2(n_150),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_201),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_129),
.A2(n_73),
.B1(n_82),
.B2(n_93),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_73),
.B1(n_80),
.B2(n_106),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_128),
.A2(n_115),
.B1(n_156),
.B2(n_125),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_196),
.B1(n_124),
.B2(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_115),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_131),
.B1(n_143),
.B2(n_141),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_132),
.B(n_146),
.C(n_127),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_141),
.B1(n_160),
.B2(n_144),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_143),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_152),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_135),
.B(n_145),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_176),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_136),
.B(n_141),
.C(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_218),
.Y(n_237)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_168),
.B(n_123),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_213),
.B(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_122),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_120),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_221),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_143),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_231),
.B1(n_171),
.B2(n_206),
.Y(n_242)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_181),
.B(n_126),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_179),
.C(n_183),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_163),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_234),
.B(n_191),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_180),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_227),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_229),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_192),
.A2(n_197),
.B1(n_184),
.B2(n_200),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_149),
.B1(n_134),
.B2(n_121),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_176),
.A2(n_165),
.B1(n_162),
.B2(n_140),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_235),
.Y(n_241)
);

AND2x6_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_140),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_175),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_247),
.C(n_255),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_186),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_231),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_219),
.A2(n_174),
.B1(n_187),
.B2(n_191),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_173),
.C(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_212),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_206),
.A2(n_172),
.B1(n_180),
.B2(n_148),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_172),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_223),
.C(n_209),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_258),
.C(n_260),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_205),
.C(n_211),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_216),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_259),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_269),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_267),
.A2(n_282),
.B1(n_269),
.B2(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_226),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_277),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_239),
.A2(n_212),
.B1(n_234),
.B2(n_204),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_260),
.B1(n_249),
.B2(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_245),
.A2(n_208),
.B(n_220),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_274),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

AOI221xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_229),
.B1(n_239),
.B2(n_246),
.C(n_241),
.Y(n_277)
);

AO221x1_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_236),
.B1(n_261),
.B2(n_259),
.C(n_238),
.Y(n_278)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_255),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_281),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_252),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_280),
.A2(n_257),
.B1(n_251),
.B2(n_238),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_237),
.B(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_243),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_287),
.B1(n_275),
.B2(n_263),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_293),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_249),
.B1(n_257),
.B2(n_247),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_292),
.A2(n_265),
.B1(n_282),
.B2(n_281),
.Y(n_306)
);

AOI21x1_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_236),
.B(n_271),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_300),
.B(n_306),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_265),
.C(n_266),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_305),
.C(n_284),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_264),
.B1(n_270),
.B2(n_271),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_302),
.B1(n_309),
.B2(n_306),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_266),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_276),
.Y(n_307)
);

NAND4xp25_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.C(n_262),
.D(n_292),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_268),
.Y(n_309)
);

OAI31xp33_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_294),
.A3(n_295),
.B(n_289),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_312),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_287),
.B(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.C(n_317),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_283),
.C(n_279),
.Y(n_314)
);

AOI211xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_289),
.B(n_294),
.C(n_273),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_318),
.B1(n_317),
.B2(n_312),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_303),
.B(n_305),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_320),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_278),
.B(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_310),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_325),
.C(n_323),
.Y(n_328)
);

AOI31xp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_323),
.A3(n_321),
.B(n_314),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.B(n_315),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_315),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_313),
.Y(n_331)
);


endmodule