module fake_aes_2325_n_1227 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1227);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1227;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_1198;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_1202;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_1211;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_1217;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1197;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_1200;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1201;
wire n_1191;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_1216;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1215;
wire n_286;
wire n_1174;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1078;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_1125;
wire n_773;
wire n_847;
wire n_1097;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_1094;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_1222;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_1188;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1132;
wire n_1159;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_1160;
wire n_1184;
wire n_274;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_1225;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1138;
wire n_293;
wire n_1063;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_1212;
wire n_771;
wire n_696;
wire n_735;
wire n_1091;
wire n_1203;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_1220;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1186;
wire n_864;
wire n_1167;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_1206;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_1178;
wire n_1209;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1218;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1210;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_1214;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_899;
wire n_806;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1224;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_1199;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_1221;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_1208;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_1141;
wire n_1213;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_1205;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1117;
wire n_859;
wire n_1007;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_1223;
wire n_774;
wire n_1207;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1112;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_1219;
wire n_585;
wire n_913;
wire n_1226;
wire n_845;
wire n_1190;
wire n_1204;
wire n_1025;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
INVx2_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_156), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_176), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_13), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_27), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_78), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_79), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_207), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_51), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_26), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_141), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_66), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_13), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_149), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_120), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_9), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_235), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_163), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_200), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_179), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_147), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_189), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_114), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g268 ( .A(n_86), .B(n_158), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_100), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_83), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_183), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_19), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_6), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_77), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_29), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_122), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_23), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_31), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_108), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_177), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_62), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_148), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_133), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_166), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_76), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_31), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_88), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_136), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_14), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_140), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_22), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_95), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_137), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_240), .Y(n_295) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_243), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_96), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_160), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_84), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_242), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_24), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_1), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_220), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_231), .Y(n_304) );
CKINVDCx14_ASAP7_75t_R g305 ( .A(n_101), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_97), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_57), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_144), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_19), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_150), .Y(n_310) );
INVxp33_ASAP7_75t_SL g311 ( .A(n_89), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_190), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_234), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_173), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_73), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_203), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_67), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_21), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_47), .Y(n_319) );
BUFx5_ASAP7_75t_L g320 ( .A(n_5), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_0), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_115), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_121), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_105), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_228), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_8), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_55), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_209), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_59), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_93), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_168), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_236), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_126), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_191), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_17), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_68), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_80), .Y(n_337) );
INVxp33_ASAP7_75t_SL g338 ( .A(n_132), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_216), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_103), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_18), .B(n_229), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_123), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_81), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_48), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_28), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_117), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_37), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_215), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_224), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_125), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_192), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_38), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_91), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_18), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_124), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_20), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_223), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_187), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_85), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_0), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_62), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_23), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_104), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_198), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_4), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_22), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_219), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_152), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_230), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_145), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_213), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_38), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g373 ( .A(n_221), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_24), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_50), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_193), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_33), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_169), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_170), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_43), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_217), .Y(n_381) );
INVx4_ASAP7_75t_L g382 ( .A(n_349), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_320), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_320), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_320), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_287), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_353), .B(n_1), .Y(n_387) );
OAI22xp5_ASAP7_75t_SL g388 ( .A1(n_292), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_275), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_263), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_320), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_296), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_320), .Y(n_393) );
INVx4_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_247), .B(n_2), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_305), .B(n_3), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_287), .B(n_5), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_275), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_275), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_362), .B(n_7), .Y(n_400) );
INVx4_ASAP7_75t_L g401 ( .A(n_267), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_275), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_312), .B(n_7), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_297), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_297), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_245), .A2(n_70), .B(n_69), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_362), .B(n_8), .Y(n_407) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_337), .B(n_244), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_297), .B(n_9), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_320), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_297), .B(n_10), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_248), .B(n_10), .Y(n_412) );
INVx6_ASAP7_75t_L g413 ( .A(n_267), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_355), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_249), .B(n_11), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_396), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_386), .B(n_305), .Y(n_417) );
BUFx4f_ASAP7_75t_L g418 ( .A(n_397), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_386), .B(n_373), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
INVx4_ASAP7_75t_L g422 ( .A(n_397), .Y(n_422) );
INVx4_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_382), .B(n_245), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_389), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_389), .Y(n_427) );
AND2x6_ASAP7_75t_L g428 ( .A(n_397), .B(n_294), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_413), .Y(n_429) );
AND2x6_ASAP7_75t_L g430 ( .A(n_400), .B(n_294), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_389), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_413), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_382), .B(n_277), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_382), .B(n_379), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_396), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_394), .B(n_392), .Y(n_438) );
INVx4_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_408), .B(n_265), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_389), .Y(n_441) );
AND2x6_ASAP7_75t_L g442 ( .A(n_400), .B(n_295), .Y(n_442) );
NOR2xp33_ASAP7_75t_SL g443 ( .A(n_408), .B(n_263), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_394), .B(n_262), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_400), .B(n_407), .Y(n_445) );
INVx5_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_401), .B(n_246), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_384), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_396), .B(n_354), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_385), .Y(n_450) );
INVx4_ASAP7_75t_SL g451 ( .A(n_413), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_387), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_413), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_389), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_401), .B(n_251), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_407), .A2(n_408), .B1(n_403), .B2(n_387), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_385), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_452), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_459), .A2(n_403), .B1(n_280), .B2(n_286), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_458), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_417), .B(n_395), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_417), .B(n_395), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_437), .B(n_401), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_458), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_438), .B(n_412), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_449), .B(n_390), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_437), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_420), .B(n_401), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_420), .B(n_265), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_422), .B(n_412), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_458), .Y(n_476) );
AO22x1_ASAP7_75t_L g477 ( .A1(n_449), .A2(n_390), .B1(n_311), .B2(n_338), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_422), .B(n_415), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_445), .A2(n_391), .B1(n_410), .B2(n_393), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_418), .A2(n_393), .B(n_410), .C(n_391), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_434), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_443), .A2(n_388), .B1(n_345), .B2(n_360), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_418), .B(n_252), .Y(n_484) );
INVx4_ASAP7_75t_L g485 ( .A(n_446), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_440), .A2(n_411), .B(n_409), .C(n_253), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_435), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_422), .B(n_311), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_423), .B(n_338), .Y(n_489) );
BUFx4f_ASAP7_75t_L g490 ( .A(n_428), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_443), .A2(n_280), .B1(n_286), .B2(n_284), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
NOR2x1p5_ASAP7_75t_L g493 ( .A(n_423), .B(n_274), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_458), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_423), .B(n_250), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_423), .B(n_259), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_429), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_439), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_439), .B(n_264), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_445), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_418), .A2(n_284), .B1(n_314), .B2(n_310), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_454), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_439), .B(n_269), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_418), .A2(n_320), .B1(n_260), .B2(n_273), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_428), .A2(n_276), .B1(n_279), .B2(n_257), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_454), .B(n_271), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_447), .A2(n_310), .B1(n_381), .B2(n_314), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_428), .A2(n_381), .B1(n_388), .B2(n_380), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_446), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_447), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_446), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_428), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_428), .A2(n_301), .B1(n_307), .B2(n_290), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_456), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_446), .B(n_255), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_428), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_446), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_446), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_446), .B(n_258), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_430), .A2(n_318), .B1(n_319), .B2(n_309), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_429), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_430), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_430), .A2(n_327), .B1(n_329), .B2(n_326), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_430), .B(n_288), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_430), .B(n_293), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_429), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_433), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_430), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_430), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_442), .B(n_366), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_444), .B(n_334), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_442), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_442), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_442), .B(n_375), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_442), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_442), .B(n_304), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_433), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_442), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_461), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_465), .B(n_421), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_492), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_499), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_508), .A2(n_302), .B1(n_321), .B2(n_282), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_466), .B(n_421), .Y(n_546) );
BUFx3_ASAP7_75t_L g547 ( .A(n_464), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_469), .A2(n_431), .B(n_448), .C(n_424), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_494), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_469), .A2(n_431), .B(n_448), .C(n_424), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_470), .B(n_292), .Y(n_551) );
NOR3xp33_ASAP7_75t_SL g552 ( .A(n_483), .B(n_356), .C(n_344), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_471), .A2(n_460), .B(n_450), .C(n_347), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_506), .A2(n_345), .B1(n_360), .B2(n_352), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_473), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_475), .B(n_460), .Y(n_557) );
NOR2xp67_ASAP7_75t_SL g558 ( .A(n_540), .B(n_365), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_462), .B(n_372), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_478), .A2(n_453), .B(n_406), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_474), .A2(n_361), .B(n_377), .C(n_335), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_501), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_499), .Y(n_563) );
NOR2xp33_ASAP7_75t_SL g564 ( .A(n_490), .B(n_308), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_488), .A2(n_453), .B(n_406), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_540), .Y(n_566) );
CKINVDCx16_ASAP7_75t_R g567 ( .A(n_502), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_491), .B(n_254), .Y(n_568) );
O2A1O1Ixp33_ASAP7_75t_L g569 ( .A1(n_481), .A2(n_256), .B(n_278), .C(n_254), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_536), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_480), .B(n_256), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_503), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_506), .A2(n_278), .B1(n_266), .B2(n_270), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_474), .A2(n_453), .B(n_406), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_493), .B(n_451), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_484), .A2(n_406), .B(n_457), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_477), .B(n_457), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_467), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_463), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_540), .B(n_315), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_505), .B(n_406), .C(n_374), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_511), .A2(n_341), .B(n_272), .C(n_281), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_472), .Y(n_583) );
AO32x2_ASAP7_75t_L g584 ( .A1(n_518), .A2(n_414), .A3(n_404), .B1(n_268), .B2(n_355), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_509), .B(n_341), .C(n_283), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_540), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_482), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_463), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_489), .B(n_322), .Y(n_589) );
NOR3xp33_ASAP7_75t_SL g590 ( .A(n_486), .B(n_331), .C(n_330), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_487), .Y(n_591) );
INVx4_ASAP7_75t_L g592 ( .A(n_485), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_514), .A2(n_525), .B1(n_522), .B2(n_516), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_481), .A2(n_285), .B(n_289), .C(n_261), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_489), .B(n_332), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_515), .B(n_374), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_490), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_468), .A2(n_427), .B(n_419), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_514), .A2(n_298), .B1(n_299), .B2(n_291), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_534), .B(n_343), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_468), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_476), .Y(n_602) );
AO32x2_ASAP7_75t_L g603 ( .A1(n_535), .A2(n_414), .A3(n_404), .B1(n_355), .B2(n_374), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_533), .B(n_451), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_507), .B(n_351), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_522), .A2(n_300), .B1(n_317), .B2(n_303), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_495), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_533), .B(n_324), .C(n_323), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_534), .B(n_368), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_524), .B(n_371), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_479), .B(n_325), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_525), .A2(n_333), .B1(n_336), .B2(n_328), .Y(n_612) );
AND2x2_ASAP7_75t_SL g613 ( .A(n_485), .B(n_339), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_479), .B(n_340), .Y(n_614) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_485), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_523), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_505), .B(n_11), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_530), .A2(n_537), .B1(n_531), .B2(n_513), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_498), .B(n_342), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_496), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_510), .B(n_346), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_510), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_497), .Y(n_623) );
NOR2xp67_ASAP7_75t_L g624 ( .A(n_500), .B(n_12), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_517), .A2(n_441), .B(n_432), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_504), .B(n_348), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_539), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_523), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_498), .B(n_350), .Y(n_629) );
AOI33xp33_ASAP7_75t_L g630 ( .A1(n_528), .A2(n_370), .A3(n_357), .B1(n_358), .B2(n_359), .B3(n_363), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_517), .Y(n_631) );
CKINVDCx16_ASAP7_75t_R g632 ( .A(n_526), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_528), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_512), .B(n_12), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_527), .A2(n_455), .B(n_364), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_529), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_538), .A2(n_455), .B(n_369), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_512), .Y(n_638) );
BUFx3_ASAP7_75t_L g639 ( .A(n_519), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_519), .B(n_14), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_539), .A2(n_378), .B(n_367), .C(n_376), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_520), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_520), .B(n_295), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_521), .B(n_15), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_461), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_471), .B(n_16), .Y(n_646) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_540), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_506), .A2(n_306), .B1(n_313), .B2(n_316), .Y(n_648) );
AO32x1_ASAP7_75t_L g649 ( .A1(n_524), .A2(n_399), .A3(n_398), .B1(n_405), .B2(n_402), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_465), .B(n_306), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_461), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_508), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_506), .A2(n_398), .B1(n_399), .B2(n_402), .Y(n_653) );
AO21x1_ASAP7_75t_L g654 ( .A1(n_484), .A2(n_405), .B(n_404), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_465), .B(n_16), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_465), .B(n_17), .Y(n_656) );
BUFx10_ASAP7_75t_L g657 ( .A(n_493), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_551), .B(n_20), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_569), .A2(n_405), .B(n_355), .C(n_414), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_574), .A2(n_436), .B(n_426), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_565), .A2(n_436), .B(n_426), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_587), .B(n_21), .Y(n_662) );
AO31x2_ASAP7_75t_L g663 ( .A1(n_560), .A2(n_414), .A3(n_404), .B(n_436), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_591), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_554), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_613), .A2(n_404), .B1(n_414), .B2(n_29), .Y(n_666) );
AO21x2_ASAP7_75t_L g667 ( .A1(n_581), .A2(n_414), .B(n_404), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_541), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_547), .B(n_25), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_645), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_657), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_548), .A2(n_414), .B(n_404), .C(n_436), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_557), .A2(n_436), .B(n_426), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_576), .A2(n_426), .B(n_72), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_652), .B(n_28), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_592), .B(n_71), .Y(n_676) );
BUFx2_ASAP7_75t_L g677 ( .A(n_554), .Y(n_677) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_615), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_572), .B(n_30), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_593), .A2(n_30), .B1(n_32), .B2(n_33), .Y(n_680) );
BUFx3_ASAP7_75t_L g681 ( .A(n_657), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_590), .B(n_608), .C(n_595), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_581), .A2(n_75), .B(n_74), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_559), .B(n_32), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g685 ( .A1(n_594), .A2(n_426), .B(n_35), .C(n_36), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_646), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_542), .A2(n_87), .B(n_82), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_651), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_567), .B(n_34), .Y(n_689) );
AO21x2_ASAP7_75t_L g690 ( .A1(n_654), .A2(n_92), .B(n_90), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g691 ( .A1(n_546), .A2(n_637), .B(n_635), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_571), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_552), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_555), .B(n_34), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_561), .B(n_35), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_553), .A2(n_36), .B(n_37), .C(n_39), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_568), .B(n_39), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_SL g698 ( .A1(n_582), .A2(n_143), .B(n_241), .C(n_239), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_596), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_571), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_L g701 ( .A1(n_641), .A2(n_40), .B(n_41), .C(n_42), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_592), .B(n_40), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_655), .Y(n_703) );
CKINVDCx11_ASAP7_75t_R g704 ( .A(n_615), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_656), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_545), .B(n_41), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_556), .B(n_42), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_585), .A2(n_43), .B1(n_44), .B2(n_45), .C(n_46), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_570), .B(n_44), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g710 ( .A(n_623), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_578), .A2(n_146), .B(n_238), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_630), .A2(n_45), .B(n_46), .C(n_47), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_544), .Y(n_713) );
CKINVDCx6p67_ASAP7_75t_R g714 ( .A(n_575), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g715 ( .A1(n_626), .A2(n_48), .B(n_49), .Y(n_715) );
BUFx10_ASAP7_75t_L g716 ( .A(n_575), .Y(n_716) );
BUFx3_ASAP7_75t_L g717 ( .A(n_615), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_593), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_564), .B(n_52), .Y(n_719) );
AOI221x1_ASAP7_75t_L g720 ( .A1(n_648), .A2(n_52), .B1(n_53), .B2(n_54), .C(n_55), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_566), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_604), .A2(n_154), .B(n_233), .Y(n_722) );
OAI21x1_ASAP7_75t_L g723 ( .A1(n_625), .A2(n_153), .B(n_232), .Y(n_723) );
AOI221x1_ASAP7_75t_L g724 ( .A1(n_648), .A2(n_53), .B1(n_54), .B2(n_56), .C(n_57), .Y(n_724) );
BUFx10_ASAP7_75t_L g725 ( .A(n_619), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_624), .A2(n_56), .B(n_58), .C(n_59), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_639), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_620), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_632), .B(n_58), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_573), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_583), .B(n_60), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_577), .A2(n_60), .B(n_61), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_563), .A2(n_157), .B(n_227), .Y(n_733) );
AO31x2_ASAP7_75t_L g734 ( .A1(n_573), .A2(n_599), .A3(n_653), .B(n_644), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g735 ( .A1(n_589), .A2(n_61), .B(n_63), .C(n_64), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_638), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_621), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g738 ( .A(n_564), .B(n_63), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_599), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_739) );
O2A1O1Ixp33_ASAP7_75t_L g740 ( .A1(n_650), .A2(n_65), .B(n_94), .C(n_98), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_579), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_588), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_543), .B(n_99), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_621), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_602), .Y(n_745) );
AO32x2_ASAP7_75t_L g746 ( .A1(n_653), .A2(n_102), .A3(n_106), .B1(n_107), .B2(n_109), .Y(n_746) );
NOR2x1_ASAP7_75t_R g747 ( .A(n_617), .B(n_110), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_605), .B(n_111), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_549), .B(n_112), .Y(n_749) );
AND2x4_ASAP7_75t_L g750 ( .A(n_562), .B(n_113), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_607), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_619), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_606), .A2(n_116), .B(n_118), .C(n_119), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_629), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_634), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_598), .A2(n_127), .B(n_128), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_640), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_612), .A2(n_129), .B(n_130), .C(n_131), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_629), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_601), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_566), .Y(n_761) );
AOI21xp33_ASAP7_75t_L g762 ( .A1(n_611), .A2(n_134), .B(n_135), .Y(n_762) );
O2A1O1Ixp33_ASAP7_75t_SL g763 ( .A1(n_622), .A2(n_138), .B(n_139), .C(n_142), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_L g764 ( .A1(n_614), .A2(n_151), .B(n_155), .C(n_159), .Y(n_764) );
BUFx10_ASAP7_75t_L g765 ( .A(n_586), .Y(n_765) );
CKINVDCx6p67_ASAP7_75t_R g766 ( .A(n_642), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_616), .Y(n_767) );
INVxp67_ASAP7_75t_L g768 ( .A(n_622), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_627), .B(n_161), .Y(n_769) );
AO21x1_ASAP7_75t_L g770 ( .A1(n_643), .A2(n_162), .B(n_164), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_649), .A2(n_165), .B(n_167), .Y(n_771) );
O2A1O1Ixp33_ASAP7_75t_SL g772 ( .A1(n_580), .A2(n_171), .B(n_172), .C(n_174), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g773 ( .A1(n_628), .A2(n_175), .B(n_178), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_L g774 ( .A1(n_610), .A2(n_180), .B(n_181), .C(n_182), .Y(n_774) );
CKINVDCx6p67_ASAP7_75t_R g775 ( .A(n_597), .Y(n_775) );
O2A1O1Ixp33_ASAP7_75t_L g776 ( .A1(n_600), .A2(n_184), .B(n_185), .C(n_186), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_633), .Y(n_777) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_586), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_649), .A2(n_188), .B(n_194), .Y(n_779) );
O2A1O1Ixp33_ASAP7_75t_L g780 ( .A1(n_609), .A2(n_195), .B(n_196), .C(n_197), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_636), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_584), .Y(n_782) );
INVx4_ASAP7_75t_L g783 ( .A(n_586), .Y(n_783) );
OA21x2_ASAP7_75t_L g784 ( .A1(n_661), .A2(n_649), .B(n_584), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_730), .A2(n_618), .B1(n_647), .B2(n_631), .Y(n_785) );
OA21x2_ASAP7_75t_L g786 ( .A1(n_660), .A2(n_584), .B(n_603), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_670), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_688), .Y(n_788) );
INVx4_ASAP7_75t_SL g789 ( .A(n_669), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_677), .B(n_597), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_728), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_736), .B(n_603), .Y(n_792) );
OA21x2_ASAP7_75t_L g793 ( .A1(n_782), .A2(n_558), .B(n_647), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_664), .Y(n_794) );
OA21x2_ASAP7_75t_L g795 ( .A1(n_683), .A2(n_647), .B(n_201), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_668), .Y(n_796) );
INVx2_ASAP7_75t_SL g797 ( .A(n_725), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_692), .B(n_597), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_669), .Y(n_799) );
OAI221xp5_ASAP7_75t_L g800 ( .A1(n_658), .A2(n_199), .B1(n_202), .B2(n_204), .C(n_205), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_679), .Y(n_801) );
AO31x2_ASAP7_75t_L g802 ( .A1(n_672), .A2(n_206), .A3(n_208), .B(n_210), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_679), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_684), .B(n_212), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_682), .A2(n_214), .B1(n_218), .B2(n_222), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_725), .B(n_225), .Y(n_806) );
OAI221xp5_ASAP7_75t_SL g807 ( .A1(n_739), .A2(n_706), .B1(n_708), .B2(n_665), .C(n_689), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_697), .B(n_226), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_694), .B(n_703), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_705), .B(n_752), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_680), .A2(n_718), .B1(n_729), .B2(n_686), .C(n_695), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_754), .B(n_759), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_737), .B(n_744), .Y(n_813) );
OA21x2_ASAP7_75t_L g814 ( .A1(n_723), .A2(n_779), .B(n_771), .Y(n_814) );
INVx3_ASAP7_75t_L g815 ( .A(n_717), .Y(n_815) );
AO21x2_ASAP7_75t_L g816 ( .A1(n_667), .A2(n_659), .B(n_711), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_702), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_710), .B(n_714), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_673), .A2(n_691), .B(n_667), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_768), .B(n_731), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_769), .A2(n_743), .B(n_698), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_760), .Y(n_822) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_704), .Y(n_823) );
A2O1A1Ixp33_ASAP7_75t_L g824 ( .A1(n_715), .A2(n_701), .B(n_748), .C(n_685), .Y(n_824) );
AND2x4_ASAP7_75t_L g825 ( .A(n_727), .B(n_750), .Y(n_825) );
AO31x2_ASAP7_75t_L g826 ( .A1(n_770), .A2(n_720), .A3(n_724), .B(n_712), .Y(n_826) );
BUFx3_ASAP7_75t_L g827 ( .A(n_766), .Y(n_827) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_678), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_662), .B(n_707), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_713), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_702), .B(n_739), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_750), .A2(n_763), .B(n_722), .Y(n_832) );
OA21x2_ASAP7_75t_L g833 ( .A1(n_687), .A2(n_773), .B(n_733), .Y(n_833) );
OR2x6_ASAP7_75t_L g834 ( .A(n_671), .B(n_681), .Y(n_834) );
A2O1A1Ixp33_ASAP7_75t_L g835 ( .A1(n_715), .A2(n_740), .B(n_675), .C(n_749), .Y(n_835) );
OAI221xp5_ASAP7_75t_L g836 ( .A1(n_696), .A2(n_709), .B1(n_735), .B2(n_726), .C(n_666), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_755), .A2(n_757), .B1(n_693), .B2(n_699), .Y(n_837) );
A2O1A1Ixp33_ASAP7_75t_L g838 ( .A1(n_732), .A2(n_738), .B(n_780), .C(n_776), .Y(n_838) );
AOI21xp33_ASAP7_75t_L g839 ( .A1(n_747), .A2(n_764), .B(n_719), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_716), .B(n_777), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_741), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_734), .B(n_747), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_734), .B(n_751), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_678), .B(n_676), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_742), .A2(n_745), .B1(n_781), .B2(n_767), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_690), .A2(n_756), .B(n_774), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_716), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_775), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_678), .Y(n_849) );
AOI321xp33_ASAP7_75t_L g850 ( .A1(n_753), .A2(n_758), .A3(n_762), .B1(n_734), .B2(n_746), .C(n_690), .Y(n_850) );
AND2x4_ASAP7_75t_L g851 ( .A(n_783), .B(n_778), .Y(n_851) );
BUFx6f_ASAP7_75t_L g852 ( .A(n_721), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_783), .A2(n_721), .B1(n_761), .B2(n_778), .Y(n_853) );
A2O1A1Ixp33_ASAP7_75t_L g854 ( .A1(n_721), .A2(n_761), .B(n_778), .C(n_746), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g855 ( .A1(n_772), .A2(n_761), .B(n_663), .Y(n_855) );
OAI21x1_ASAP7_75t_SL g856 ( .A1(n_746), .A2(n_765), .B(n_663), .Y(n_856) );
AO31x2_ASAP7_75t_L g857 ( .A1(n_765), .A2(n_782), .A3(n_672), .B(n_661), .Y(n_857) );
BUFx8_ASAP7_75t_SL g858 ( .A(n_681), .Y(n_858) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_704), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_704), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_728), .B(n_452), .Y(n_861) );
OR2x6_ASAP7_75t_L g862 ( .A(n_669), .B(n_508), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_677), .B(n_587), .Y(n_863) );
AO31x2_ASAP7_75t_L g864 ( .A1(n_782), .A2(n_672), .A3(n_661), .B(n_660), .Y(n_864) );
BUFx12f_ASAP7_75t_L g865 ( .A(n_704), .Y(n_865) );
INVx4_ASAP7_75t_L g866 ( .A(n_704), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_670), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_677), .B(n_587), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g869 ( .A1(n_692), .A2(n_700), .B(n_682), .C(n_658), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_660), .A2(n_661), .B(n_574), .Y(n_870) );
OAI21xp5_ASAP7_75t_L g871 ( .A1(n_691), .A2(n_550), .B(n_548), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_668), .Y(n_872) );
AND2x4_ASAP7_75t_L g873 ( .A(n_692), .B(n_587), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_L g874 ( .A1(n_692), .A2(n_700), .B(n_682), .C(n_658), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_692), .B(n_700), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_677), .A2(n_483), .B1(n_551), .B2(n_730), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_728), .B(n_452), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_692), .B(n_700), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_668), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g880 ( .A1(n_677), .A2(n_508), .B1(n_443), .B2(n_730), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_668), .Y(n_881) );
INVx1_ASAP7_75t_SL g882 ( .A(n_704), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_670), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_704), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_728), .B(n_452), .Y(n_885) );
OAI21x1_ASAP7_75t_L g886 ( .A1(n_660), .A2(n_661), .B(n_674), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g887 ( .A1(n_660), .A2(n_661), .B(n_574), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_728), .B(n_452), .Y(n_888) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_660), .A2(n_661), .B(n_574), .Y(n_889) );
INVx3_ASAP7_75t_L g890 ( .A(n_717), .Y(n_890) );
BUFx2_ASAP7_75t_L g891 ( .A(n_728), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_677), .A2(n_551), .B1(n_483), .B2(n_554), .C(n_555), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_670), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_660), .A2(n_661), .B(n_574), .Y(n_894) );
OR2x6_ASAP7_75t_L g895 ( .A(n_669), .B(n_508), .Y(n_895) );
OR2x6_ASAP7_75t_L g896 ( .A(n_669), .B(n_508), .Y(n_896) );
AND2x4_ASAP7_75t_L g897 ( .A(n_692), .B(n_587), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_692), .B(n_700), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_677), .A2(n_508), .B1(n_443), .B2(n_730), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_794), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_791), .B(n_891), .Y(n_901) );
AO21x2_ASAP7_75t_L g902 ( .A1(n_870), .A2(n_894), .B(n_889), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_787), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_788), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_892), .B(n_876), .Y(n_905) );
AO21x2_ASAP7_75t_L g906 ( .A1(n_887), .A2(n_819), .B(n_856), .Y(n_906) );
NAND2x1p5_ASAP7_75t_L g907 ( .A(n_827), .B(n_825), .Y(n_907) );
AO31x2_ASAP7_75t_L g908 ( .A1(n_854), .A2(n_843), .A3(n_842), .B(n_835), .Y(n_908) );
AND2x4_ASAP7_75t_L g909 ( .A(n_789), .B(n_851), .Y(n_909) );
OR2x6_ASAP7_75t_L g910 ( .A(n_831), .B(n_825), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_867), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_883), .Y(n_912) );
BUFx2_ASAP7_75t_L g913 ( .A(n_789), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_893), .Y(n_914) );
OA21x2_ASAP7_75t_L g915 ( .A1(n_886), .A2(n_855), .B(n_846), .Y(n_915) );
OR2x2_ASAP7_75t_L g916 ( .A(n_872), .B(n_879), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_796), .Y(n_917) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_873), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_822), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_881), .B(n_875), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_862), .A2(n_896), .B1(n_895), .B2(n_799), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_810), .Y(n_922) );
BUFx3_ASAP7_75t_L g923 ( .A(n_884), .Y(n_923) );
BUFx2_ASAP7_75t_L g924 ( .A(n_834), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_875), .B(n_878), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_878), .B(n_898), .Y(n_926) );
AND2x4_ASAP7_75t_L g927 ( .A(n_851), .B(n_849), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_898), .B(n_830), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_813), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_841), .B(n_813), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_873), .B(n_897), .Y(n_931) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_869), .B(n_874), .C(n_807), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_897), .B(n_861), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_812), .Y(n_934) );
OR2x6_ASAP7_75t_L g935 ( .A(n_862), .B(n_895), .Y(n_935) );
INVx1_ASAP7_75t_SL g936 ( .A(n_858), .Y(n_936) );
OR2x6_ASAP7_75t_L g937 ( .A(n_862), .B(n_895), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_896), .B(n_863), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_896), .B(n_868), .Y(n_939) );
AO21x2_ASAP7_75t_L g940 ( .A1(n_871), .A2(n_824), .B(n_816), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_880), .A2(n_899), .B1(n_811), .B2(n_837), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g942 ( .A1(n_809), .A2(n_877), .B1(n_885), .B2(n_888), .C(n_836), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_834), .Y(n_943) );
OR2x6_ASAP7_75t_L g944 ( .A(n_785), .B(n_817), .Y(n_944) );
OR2x2_ASAP7_75t_L g945 ( .A(n_829), .B(n_803), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_792), .B(n_845), .Y(n_946) );
AO21x2_ASAP7_75t_L g947 ( .A1(n_816), .A2(n_821), .B(n_832), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_801), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_840), .Y(n_949) );
INVxp67_ASAP7_75t_L g950 ( .A(n_834), .Y(n_950) );
OAI21xp5_ASAP7_75t_L g951 ( .A1(n_838), .A2(n_839), .B(n_820), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_804), .B(n_790), .Y(n_952) );
AOI211xp5_ASAP7_75t_L g953 ( .A1(n_839), .A2(n_882), .B(n_785), .C(n_847), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_797), .B(n_798), .Y(n_954) );
NAND4xp25_ASAP7_75t_L g955 ( .A(n_818), .B(n_882), .C(n_866), .D(n_850), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_848), .B(n_815), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_890), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_890), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_864), .Y(n_959) );
OR2x2_ASAP7_75t_L g960 ( .A(n_823), .B(n_859), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_786), .Y(n_961) );
OAI21xp5_ASAP7_75t_L g962 ( .A1(n_808), .A2(n_800), .B(n_844), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_815), .B(n_849), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_828), .B(n_852), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_806), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_852), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_852), .Y(n_967) );
INVx3_ASAP7_75t_L g968 ( .A(n_828), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_823), .Y(n_969) );
OR2x6_ASAP7_75t_L g970 ( .A(n_828), .B(n_866), .Y(n_970) );
OAI21xp33_ASAP7_75t_L g971 ( .A1(n_805), .A2(n_860), .B(n_853), .Y(n_971) );
BUFx3_ASAP7_75t_L g972 ( .A(n_823), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_784), .Y(n_973) );
AND2x4_ASAP7_75t_L g974 ( .A(n_857), .B(n_802), .Y(n_974) );
OR2x6_ASAP7_75t_L g975 ( .A(n_859), .B(n_865), .Y(n_975) );
OR2x6_ASAP7_75t_L g976 ( .A(n_793), .B(n_795), .Y(n_976) );
AOI221xp5_ASAP7_75t_L g977 ( .A1(n_826), .A2(n_857), .B1(n_784), .B2(n_833), .C(n_814), .Y(n_977) );
BUFx3_ASAP7_75t_L g978 ( .A(n_793), .Y(n_978) );
AND2x4_ASAP7_75t_L g979 ( .A(n_826), .B(n_814), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_833), .B(n_795), .Y(n_980) );
INVx3_ASAP7_75t_L g981 ( .A(n_828), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_961), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_925), .B(n_946), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_925), .B(n_946), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_926), .B(n_938), .Y(n_985) );
OAI321xp33_ASAP7_75t_L g986 ( .A1(n_932), .A2(n_955), .A3(n_941), .B1(n_937), .B2(n_935), .C(n_951), .Y(n_986) );
BUFx2_ASAP7_75t_L g987 ( .A(n_978), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_938), .B(n_939), .Y(n_988) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_923), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_973), .Y(n_990) );
BUFx2_ASAP7_75t_L g991 ( .A(n_978), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_920), .B(n_928), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_920), .B(n_928), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_930), .B(n_939), .Y(n_994) );
BUFx2_ASAP7_75t_L g995 ( .A(n_964), .Y(n_995) );
OR2x2_ASAP7_75t_L g996 ( .A(n_935), .B(n_937), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_930), .B(n_940), .Y(n_997) );
AOI21xp5_ASAP7_75t_L g998 ( .A1(n_902), .A2(n_915), .B(n_976), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_940), .B(n_935), .Y(n_999) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_964), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_929), .B(n_903), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_940), .B(n_937), .Y(n_1002) );
INVx4_ASAP7_75t_L g1003 ( .A(n_909), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_919), .B(n_904), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_911), .B(n_912), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_964), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_902), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_914), .B(n_917), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_952), .B(n_910), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1010 ( .A1(n_902), .A2(n_915), .B(n_976), .Y(n_1010) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_924), .Y(n_1011) );
INVx4_ASAP7_75t_L g1012 ( .A(n_909), .Y(n_1012) );
INVx2_ASAP7_75t_SL g1013 ( .A(n_909), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_910), .B(n_945), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_918), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_952), .B(n_910), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_910), .B(n_979), .Y(n_1017) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_945), .B(n_933), .Y(n_1018) );
NOR2x1_ASAP7_75t_L g1019 ( .A(n_913), .B(n_943), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_922), .B(n_944), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_979), .B(n_931), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_901), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_944), .B(n_916), .Y(n_1023) );
AO21x2_ASAP7_75t_L g1024 ( .A1(n_947), .A2(n_906), .B(n_980), .Y(n_1024) );
INVx2_ASAP7_75t_SL g1025 ( .A(n_968), .Y(n_1025) );
AO21x2_ASAP7_75t_L g1026 ( .A1(n_947), .A2(n_906), .B(n_980), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_944), .B(n_934), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_944), .B(n_942), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_979), .B(n_931), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1030 ( .A(n_968), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_954), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_900), .B(n_948), .Y(n_1032) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_968), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_992), .B(n_921), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_992), .B(n_905), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1005), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_993), .B(n_953), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1005), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_982), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_985), .B(n_949), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_993), .B(n_954), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_983), .B(n_965), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_997), .B(n_959), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1008), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_983), .B(n_950), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1008), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_994), .B(n_963), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1004), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1004), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_984), .B(n_958), .Y(n_1050) );
INVx5_ASAP7_75t_L g1051 ( .A(n_1003), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1032), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1032), .Y(n_1053) );
AND2x4_ASAP7_75t_L g1054 ( .A(n_1017), .B(n_906), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1001), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1001), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_994), .B(n_963), .Y(n_1057) );
NAND4xp25_ASAP7_75t_L g1058 ( .A(n_1028), .B(n_971), .C(n_956), .D(n_923), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_985), .B(n_960), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_984), .B(n_969), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1031), .Y(n_1061) );
INVxp67_ASAP7_75t_L g1062 ( .A(n_987), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1018), .B(n_957), .Y(n_1063) );
INVx2_ASAP7_75t_SL g1064 ( .A(n_1019), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_987), .Y(n_1065) );
OAI31xp33_ASAP7_75t_L g1066 ( .A1(n_1028), .A2(n_907), .A3(n_936), .B(n_972), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1018), .B(n_927), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1021), .B(n_972), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1015), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_988), .B(n_970), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1021), .B(n_927), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_988), .B(n_970), .Y(n_1072) );
AND2x4_ASAP7_75t_L g1073 ( .A(n_1017), .B(n_997), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1022), .B(n_927), .Y(n_1074) );
NAND2x1p5_ASAP7_75t_L g1075 ( .A(n_1003), .B(n_981), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_999), .B(n_974), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1009), .B(n_907), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1029), .B(n_908), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1011), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1009), .B(n_970), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1011), .Y(n_1081) );
INVxp67_ASAP7_75t_L g1082 ( .A(n_991), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_999), .B(n_974), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_986), .B(n_970), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1016), .B(n_966), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1020), .B(n_967), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1002), .B(n_908), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1020), .B(n_977), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1002), .B(n_908), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_991), .Y(n_1090) );
NOR2x1_ASAP7_75t_L g1091 ( .A(n_1019), .B(n_975), .Y(n_1091) );
INVx1_ASAP7_75t_SL g1092 ( .A(n_1068), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1061), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1044), .B(n_1027), .Y(n_1094) );
NOR2x2_ASAP7_75t_L g1095 ( .A(n_1091), .B(n_975), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1048), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1049), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1078), .B(n_1024), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1046), .B(n_1027), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1078), .B(n_1026), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1101 ( .A(n_1051), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1052), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1043), .B(n_1026), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1039), .Y(n_1104) );
NAND2x1p5_ASAP7_75t_L g1105 ( .A(n_1051), .B(n_1012), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1053), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1041), .B(n_1014), .Y(n_1107) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1039), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1043), .B(n_1026), .Y(n_1109) );
INVxp67_ASAP7_75t_L g1110 ( .A(n_1059), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1087), .B(n_1026), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1112 ( .A(n_1065), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1069), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1036), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1087), .B(n_1024), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1073), .B(n_1023), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1055), .B(n_1014), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_1065), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1089), .B(n_1024), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1073), .B(n_1023), .Y(n_1120) );
INVxp67_ASAP7_75t_SL g1121 ( .A(n_1090), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1056), .B(n_990), .Y(n_1122) );
OR2x6_ASAP7_75t_L g1123 ( .A(n_1064), .B(n_996), .Y(n_1123) );
INVx3_ASAP7_75t_L g1124 ( .A(n_1051), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1089), .B(n_1024), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1038), .Y(n_1126) );
INVx2_ASAP7_75t_SL g1127 ( .A(n_1051), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1086), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1035), .B(n_990), .Y(n_1129) );
INVxp67_ASAP7_75t_SL g1130 ( .A(n_1090), .Y(n_1130) );
NAND2x1_ASAP7_75t_L g1131 ( .A(n_1064), .B(n_1003), .Y(n_1131) );
INVxp67_ASAP7_75t_L g1132 ( .A(n_1060), .Y(n_1132) );
INVxp67_ASAP7_75t_L g1133 ( .A(n_1112), .Y(n_1133) );
NAND2xp5_ASAP7_75t_SL g1134 ( .A(n_1124), .B(n_1066), .Y(n_1134) );
INVxp67_ASAP7_75t_L g1135 ( .A(n_1118), .Y(n_1135) );
INVx1_ASAP7_75t_SL g1136 ( .A(n_1092), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1128), .B(n_1042), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_1131), .A2(n_986), .B(n_1084), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1128), .B(n_1088), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1123), .B(n_1054), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_1121), .Y(n_1141) );
OAI32xp33_ASAP7_75t_L g1142 ( .A1(n_1105), .A2(n_1058), .A3(n_1070), .B1(n_1072), .B2(n_1037), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1103), .B(n_1050), .Y(n_1143) );
NOR2x1_ASAP7_75t_L g1144 ( .A(n_1124), .B(n_975), .Y(n_1144) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1104), .Y(n_1145) );
INVx1_ASAP7_75t_SL g1146 ( .A(n_1095), .Y(n_1146) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_1123), .B(n_1054), .Y(n_1147) );
AOI22x1_ASAP7_75t_L g1148 ( .A1(n_1105), .A2(n_1003), .B1(n_1012), .B2(n_1075), .Y(n_1148) );
INVx1_ASAP7_75t_SL g1149 ( .A(n_1105), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1098), .B(n_1047), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1104), .Y(n_1151) );
AND2x4_ASAP7_75t_L g1152 ( .A(n_1123), .B(n_1054), .Y(n_1152) );
AND2x4_ASAP7_75t_L g1153 ( .A(n_1123), .B(n_1073), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1126), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1098), .B(n_1057), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1100), .B(n_1045), .Y(n_1156) );
OAI21xp5_ASAP7_75t_L g1157 ( .A1(n_1131), .A2(n_1084), .B(n_989), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1100), .B(n_1079), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1108), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1126), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1103), .B(n_1081), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1108), .Y(n_1162) );
OAI21xp33_ASAP7_75t_SL g1163 ( .A1(n_1146), .A2(n_1101), .B(n_1127), .Y(n_1163) );
A2O1A1Ixp33_ASAP7_75t_L g1164 ( .A1(n_1144), .A2(n_1124), .B(n_1101), .C(n_1127), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1139), .B(n_1111), .Y(n_1165) );
INVx2_ASAP7_75t_L g1166 ( .A(n_1145), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1154), .Y(n_1167) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_1136), .A2(n_1132), .B1(n_1116), .B2(n_1120), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1160), .Y(n_1169) );
OAI32xp33_ASAP7_75t_L g1170 ( .A1(n_1134), .A2(n_1110), .A3(n_1072), .B1(n_1012), .B2(n_1116), .Y(n_1170) );
AOI21xp5_ASAP7_75t_L g1171 ( .A1(n_1134), .A2(n_1130), .B(n_1062), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1161), .Y(n_1172) );
AOI322xp5_ASAP7_75t_L g1173 ( .A1(n_1150), .A2(n_1115), .A3(n_1125), .B1(n_1111), .B2(n_1119), .C1(n_1109), .C2(n_1113), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1155), .B(n_1115), .Y(n_1174) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_1148), .A2(n_1120), .B1(n_1012), .B2(n_1107), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_1148), .A2(n_996), .B1(n_1034), .B2(n_1040), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1143), .B(n_1109), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1161), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1141), .Y(n_1179) );
NOR3xp33_ASAP7_75t_L g1180 ( .A(n_1142), .B(n_1093), .C(n_962), .Y(n_1180) );
INVxp67_ASAP7_75t_L g1181 ( .A(n_1133), .Y(n_1181) );
INVx1_ASAP7_75t_SL g1182 ( .A(n_1149), .Y(n_1182) );
AOI211xp5_ASAP7_75t_L g1183 ( .A1(n_1163), .A2(n_1142), .B(n_1157), .C(n_1138), .Y(n_1183) );
OAI21xp5_ASAP7_75t_SL g1184 ( .A1(n_1164), .A2(n_1153), .B(n_1147), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_1180), .A2(n_1147), .B1(n_1140), .B2(n_1152), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1173), .B(n_1119), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1179), .Y(n_1187) );
A2O1A1Ixp33_ASAP7_75t_L g1188 ( .A1(n_1164), .A2(n_1153), .B(n_1152), .C(n_1147), .Y(n_1188) );
AOI211xp5_ASAP7_75t_L g1189 ( .A1(n_1170), .A2(n_1152), .B(n_1140), .C(n_1153), .Y(n_1189) );
NAND2xp5_ASAP7_75t_SL g1190 ( .A(n_1175), .B(n_1140), .Y(n_1190) );
AOI321xp33_ASAP7_75t_L g1191 ( .A1(n_1170), .A2(n_1125), .A3(n_1137), .B1(n_1074), .B2(n_1158), .C(n_1117), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_1181), .A2(n_1067), .B1(n_1077), .B2(n_1083), .Y(n_1192) );
AOI21xp5_ASAP7_75t_L g1193 ( .A1(n_1176), .A2(n_1135), .B(n_1129), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_1168), .A2(n_1143), .B1(n_1156), .B2(n_1062), .Y(n_1194) );
OAI211xp5_ASAP7_75t_L g1195 ( .A1(n_1171), .A2(n_1063), .B(n_1080), .C(n_1082), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_1186), .A2(n_1178), .B1(n_1172), .B2(n_1165), .C(n_1169), .Y(n_1196) );
NAND3xp33_ASAP7_75t_SL g1197 ( .A(n_1183), .B(n_1182), .C(n_1075), .Y(n_1197) );
O2A1O1Ixp33_ASAP7_75t_L g1198 ( .A1(n_1188), .A2(n_975), .B(n_1167), .C(n_1174), .Y(n_1198) );
OAI211xp5_ASAP7_75t_L g1199 ( .A1(n_1189), .A2(n_1177), .B(n_1114), .C(n_1082), .Y(n_1199) );
AOI21xp5_ASAP7_75t_L g1200 ( .A1(n_1184), .A2(n_1166), .B(n_1122), .Y(n_1200) );
NOR2xp33_ASAP7_75t_R g1201 ( .A(n_1187), .B(n_1013), .Y(n_1201) );
OAI211xp5_ASAP7_75t_SL g1202 ( .A1(n_1185), .A2(n_1097), .B(n_1106), .C(n_1096), .Y(n_1202) );
OAI221xp5_ASAP7_75t_L g1203 ( .A1(n_1191), .A2(n_1097), .B1(n_1102), .B2(n_1106), .C(n_1096), .Y(n_1203) );
NOR3x1_ASAP7_75t_L g1204 ( .A(n_1190), .B(n_1013), .C(n_1099), .Y(n_1204) );
NOR3xp33_ASAP7_75t_L g1205 ( .A(n_1197), .B(n_1195), .C(n_1194), .Y(n_1205) );
AOI211xp5_ASAP7_75t_L g1206 ( .A1(n_1199), .A2(n_1193), .B(n_1177), .C(n_1102), .Y(n_1206) );
AOI211xp5_ASAP7_75t_L g1207 ( .A1(n_1198), .A2(n_1010), .B(n_998), .C(n_1094), .Y(n_1207) );
OAI211xp5_ASAP7_75t_L g1208 ( .A1(n_1196), .A2(n_1192), .B(n_998), .C(n_1010), .Y(n_1208) );
NOR3xp33_ASAP7_75t_L g1209 ( .A(n_1202), .B(n_1166), .C(n_981), .Y(n_1209) );
NAND3xp33_ASAP7_75t_SL g1210 ( .A(n_1201), .B(n_1192), .C(n_1033), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_1205), .A2(n_1203), .B1(n_1200), .B2(n_1204), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_1208), .A2(n_1162), .B1(n_1159), .B2(n_1151), .C(n_1145), .Y(n_1212) );
NAND5xp2_ASAP7_75t_L g1213 ( .A(n_1207), .B(n_1000), .C(n_995), .D(n_1006), .E(n_1071), .Y(n_1213) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1209), .Y(n_1214) );
NAND3xp33_ASAP7_75t_L g1215 ( .A(n_1206), .B(n_1007), .C(n_1162), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1216 ( .A(n_1214), .Y(n_1216) );
AND2x4_ASAP7_75t_L g1217 ( .A(n_1211), .B(n_1159), .Y(n_1217) );
OR4x1_ASAP7_75t_L g1218 ( .A(n_1213), .B(n_1210), .C(n_1025), .D(n_1030), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1215), .Y(n_1219) );
NOR3xp33_ASAP7_75t_L g1220 ( .A(n_1216), .B(n_1219), .C(n_1217), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1217), .Y(n_1221) );
OAI22xp33_ASAP7_75t_SL g1222 ( .A1(n_1221), .A2(n_1218), .B1(n_1212), .B2(n_1007), .Y(n_1222) );
INVx3_ASAP7_75t_L g1223 ( .A(n_1220), .Y(n_1223) );
AOI221xp5_ASAP7_75t_L g1224 ( .A1(n_1223), .A2(n_1218), .B1(n_1007), .B2(n_1030), .C(n_1025), .Y(n_1224) );
INVxp67_ASAP7_75t_L g1225 ( .A(n_1224), .Y(n_1225) );
NAND2x2_ASAP7_75t_L g1226 ( .A(n_1225), .B(n_1222), .Y(n_1226) );
AOI22xp5_ASAP7_75t_L g1227 ( .A1(n_1226), .A2(n_1076), .B1(n_1083), .B2(n_1085), .Y(n_1227) );
endmodule