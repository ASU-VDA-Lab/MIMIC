module fake_jpeg_15995_n_392 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_392);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_392;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_33),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_45),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_19),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_37),
.B1(n_41),
.B2(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_70),
.A2(n_110),
.B1(n_48),
.B2(n_42),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_75),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_28),
.B1(n_35),
.B2(n_16),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_15),
.B1(n_24),
.B2(n_26),
.Y(n_122)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_39),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_63),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_101),
.A2(n_106),
.B(n_0),
.Y(n_142)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_61),
.A2(n_15),
.B1(n_22),
.B2(n_31),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_113),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_43),
.A2(n_31),
.B1(n_24),
.B2(n_22),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_40),
.B(n_35),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_23),
.B(n_15),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_45),
.B(n_23),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_46),
.B(n_21),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_116),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_38),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_107),
.B1(n_57),
.B2(n_105),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_119),
.A2(n_130),
.B1(n_95),
.B2(n_93),
.Y(n_179)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_33),
.B(n_26),
.C(n_30),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_121),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_122),
.A2(n_155),
.B1(n_163),
.B2(n_168),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_123),
.A2(n_8),
.B(n_135),
.Y(n_212)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_129),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_81),
.A2(n_53),
.B1(n_56),
.B2(n_47),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_24),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_135),
.Y(n_184)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_71),
.B(n_30),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_134),
.B(n_140),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_18),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_148),
.Y(n_174)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_62),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_18),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_147),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_161),
.B(n_165),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_143),
.A2(n_151),
.B1(n_152),
.B2(n_5),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_145),
.B(n_156),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_34),
.C(n_19),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_97),
.A2(n_19),
.B1(n_13),
.B2(n_12),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_84),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_83),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_107),
.B(n_0),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_162),
.Y(n_202)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

NAND2x1_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_0),
.Y(n_161)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_93),
.A2(n_8),
.B(n_4),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_86),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_172),
.Y(n_228)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_173),
.B(n_183),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_175),
.B(n_192),
.Y(n_235)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_186),
.B1(n_187),
.B2(n_160),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_199),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_89),
.B1(n_82),
.B2(n_117),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_145),
.A2(n_89),
.B1(n_82),
.B2(n_117),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_5),
.B(n_7),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_188),
.A2(n_133),
.B(n_162),
.Y(n_245)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_137),
.A2(n_5),
.B(n_8),
.C(n_94),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_R g216 ( 
.A(n_191),
.B(n_212),
.C(n_161),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_142),
.A2(n_94),
.B1(n_98),
.B2(n_115),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_166),
.B1(n_132),
.B2(n_144),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_149),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_98),
.B(n_115),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_182),
.C(n_190),
.Y(n_227)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_138),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_207),
.B(n_208),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_138),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_127),
.B(n_8),
.Y(n_210)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_139),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_213),
.Y(n_244)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_216),
.A2(n_218),
.B(n_245),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_182),
.B(n_140),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_169),
.C(n_195),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_121),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_236),
.B1(n_215),
.B2(n_178),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_220),
.A2(n_222),
.B1(n_229),
.B2(n_250),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_147),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_221),
.A2(n_230),
.B(n_255),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_137),
.B1(n_167),
.B2(n_149),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_128),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_240),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_203),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_154),
.B1(n_125),
.B2(n_159),
.Y(n_229)
);

XOR2x2_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_157),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_156),
.C(n_157),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_231),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_232),
.A2(n_246),
.B1(n_181),
.B2(n_173),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_183),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_122),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_241),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_200),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_251),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_148),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_181),
.B1(n_196),
.B2(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_191),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_171),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_253),
.Y(n_261)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_247),
.B1(n_240),
.B2(n_220),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_257),
.A2(n_264),
.B1(n_269),
.B2(n_282),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_262),
.B1(n_249),
.B2(n_237),
.Y(n_298)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_230),
.A3(n_245),
.B1(n_217),
.B2(n_221),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_263),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_179),
.B1(n_187),
.B2(n_178),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_223),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_221),
.A2(n_195),
.B1(n_171),
.B2(n_197),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_276),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_222),
.A2(n_197),
.B1(n_203),
.B2(n_180),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_277),
.B(n_279),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_172),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_276),
.Y(n_306)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_213),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_211),
.B(n_201),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_236),
.A2(n_218),
.B1(n_224),
.B2(n_228),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_226),
.A2(n_224),
.B(n_232),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_288),
.B(n_239),
.Y(n_302)
);

NAND2x1_ASAP7_75t_SL g286 ( 
.A(n_246),
.B(n_256),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_241),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_226),
.A2(n_242),
.B(n_234),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_243),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_286),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_297),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_293),
.A2(n_302),
.B(n_292),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_298),
.A2(n_293),
.B1(n_294),
.B2(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_266),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_307),
.Y(n_332)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_267),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_268),
.C(n_257),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_R g311 ( 
.A1(n_290),
.A2(n_277),
.B1(n_279),
.B2(n_274),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_311),
.B(n_269),
.CI(n_312),
.CON(n_333),
.SN(n_333)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_313),
.Y(n_327)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_314),
.Y(n_338)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_315),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_280),
.A2(n_285),
.B(n_288),
.C(n_287),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_316),
.A2(n_302),
.B(n_303),
.Y(n_340)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_317),
.A2(n_318),
.B1(n_286),
.B2(n_282),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_261),
.B(n_281),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_325),
.C(n_296),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_310),
.B(n_290),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_324),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_308),
.B(n_280),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_264),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_270),
.B1(n_287),
.B2(n_275),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_326),
.A2(n_337),
.B1(n_303),
.B2(n_301),
.Y(n_350)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_270),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_336),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_296),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_340),
.B(n_301),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_312),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_291),
.C(n_300),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_351),
.C(n_355),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_332),
.Y(n_342)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_295),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_352),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_349),
.A2(n_335),
.B(n_338),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_336),
.B(n_329),
.Y(n_366)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_328),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_354),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_340),
.A2(n_309),
.B1(n_313),
.B2(n_317),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_356),
.A2(n_358),
.B1(n_327),
.B2(n_339),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_314),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_351),
.C(n_325),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_315),
.B1(n_326),
.B2(n_328),
.Y(n_358)
);

AO21x1_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_346),
.B(n_333),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_367),
.C(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_331),
.C(n_347),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_333),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_343),
.A2(n_349),
.B(n_355),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_369),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_372),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_373),
.A2(n_369),
.B1(n_366),
.B2(n_360),
.Y(n_381)
);

AOI21xp33_ASAP7_75t_L g374 ( 
.A1(n_361),
.A2(n_341),
.B(n_329),
.Y(n_374)
);

AOI21xp33_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_376),
.B(n_364),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_345),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_377),
.A2(n_370),
.B1(n_354),
.B2(n_368),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_375),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_381),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_371),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_382),
.B(n_381),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_362),
.Y(n_386)
);

NOR3xp33_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_386),
.C(n_363),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_359),
.B(n_384),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_388),
.A2(n_379),
.B1(n_360),
.B2(n_372),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_389),
.A2(n_373),
.B(n_345),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_367),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_324),
.Y(n_392)
);


endmodule