module real_aes_10062_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1873;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_1225;
wire n_951;
wire n_1199;
wire n_875;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_1383;
wire n_552;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_948;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1800;
wire n_1435;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1802;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_1838;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_1617;
wire n_525;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_1457;
wire n_719;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_0), .A2(n_173), .B1(n_672), .B2(n_674), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_0), .A2(n_173), .B1(n_682), .B2(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_1), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_1), .A2(n_9), .B1(n_870), .B2(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g1084 ( .A(n_2), .Y(n_1084) );
AOI22xp5_ASAP7_75t_L g1578 ( .A1(n_3), .A2(n_366), .B1(n_1564), .B2(n_1567), .Y(n_1578) );
CKINVDCx5p33_ASAP7_75t_R g1814 ( .A(n_4), .Y(n_1814) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_5), .A2(n_246), .B1(n_504), .B2(n_676), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_5), .A2(n_246), .B1(n_558), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_6), .A2(n_185), .B1(n_558), .B2(n_692), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_6), .A2(n_185), .B1(n_478), .B2(n_483), .Y(n_830) );
AOI22xp33_ASAP7_75t_SL g1353 ( .A1(n_7), .A2(n_18), .B1(n_1103), .B2(n_1354), .Y(n_1353) );
INVxp67_ASAP7_75t_SL g1376 ( .A(n_7), .Y(n_1376) );
INVx1_ASAP7_75t_L g840 ( .A(n_8), .Y(n_840) );
INVx1_ASAP7_75t_L g849 ( .A(n_9), .Y(n_849) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_10), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_10), .A2(n_76), .B1(n_1281), .B2(n_1282), .Y(n_1280) );
AOI22xp33_ASAP7_75t_SL g1502 ( .A1(n_11), .A2(n_310), .B1(n_1270), .B2(n_1362), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_11), .A2(n_310), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
INVxp33_ASAP7_75t_SL g1349 ( .A(n_12), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_12), .A2(n_340), .B1(n_1043), .B2(n_1362), .Y(n_1361) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_13), .Y(n_572) );
INVx1_ASAP7_75t_L g1198 ( .A(n_14), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_14), .A2(n_223), .B1(n_1211), .B2(n_1212), .Y(n_1210) );
INVx1_ASAP7_75t_L g1393 ( .A(n_15), .Y(n_1393) );
AOI22xp33_ASAP7_75t_SL g1408 ( .A1(n_15), .A2(n_81), .B1(n_827), .B2(n_1409), .Y(n_1408) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_16), .A2(n_320), .B1(n_692), .B2(n_693), .Y(n_691) );
INVxp67_ASAP7_75t_L g710 ( .A(n_16), .Y(n_710) );
INVxp67_ASAP7_75t_SL g1345 ( .A(n_17), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_17), .A2(n_234), .B1(n_855), .B2(n_906), .Y(n_1372) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_18), .Y(n_1377) );
INVx1_ASAP7_75t_L g1499 ( .A(n_19), .Y(n_1499) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_19), .A2(n_68), .B1(n_702), .B2(n_1222), .Y(n_1506) );
AOI22xp5_ASAP7_75t_L g1864 ( .A1(n_20), .A2(n_1865), .B1(n_1866), .B2(n_1867), .Y(n_1864) );
CKINVDCx5p33_ASAP7_75t_R g1865 ( .A(n_20), .Y(n_1865) );
INVx1_ASAP7_75t_L g839 ( .A(n_21), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_21), .A2(n_73), .B1(n_827), .B2(n_865), .Y(n_873) );
INVxp33_ASAP7_75t_SL g1490 ( .A(n_22), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_22), .A2(n_112), .B1(n_1107), .B2(n_1174), .Y(n_1513) );
INVxp33_ASAP7_75t_L g1299 ( .A(n_23), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_23), .A2(n_41), .B1(n_688), .B2(n_746), .Y(n_1326) );
INVx1_ASAP7_75t_L g942 ( .A(n_24), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_24), .A2(n_343), .B1(n_386), .B2(n_401), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g1579 ( .A1(n_25), .A2(n_314), .B1(n_1557), .B2(n_1575), .Y(n_1579) );
XOR2x2_ASAP7_75t_L g1336 ( .A(n_26), .B(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g984 ( .A(n_27), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_28), .A2(n_89), .B1(n_496), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_28), .A2(n_89), .B1(n_777), .B2(n_779), .Y(n_776) );
CKINVDCx16_ASAP7_75t_R g1555 ( .A(n_29), .Y(n_1555) );
AOI22xp33_ASAP7_75t_SL g1403 ( .A1(n_30), .A2(n_272), .B1(n_504), .B2(n_676), .Y(n_1403) );
AOI22xp33_ASAP7_75t_SL g1412 ( .A1(n_30), .A2(n_272), .B1(n_589), .B2(n_1413), .Y(n_1412) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_31), .A2(n_416), .B(n_420), .C(n_425), .Y(n_415) );
INVx1_ASAP7_75t_L g509 ( .A(n_31), .Y(n_509) );
OAI222xp33_ASAP7_75t_L g1185 ( .A1(n_32), .A2(n_94), .B1(n_241), .B2(n_844), .C1(n_847), .C2(n_1186), .Y(n_1185) );
AOI22xp33_ASAP7_75t_SL g1221 ( .A1(n_32), .A2(n_201), .B1(n_1222), .B2(n_1224), .Y(n_1221) );
INVx1_ASAP7_75t_L g731 ( .A(n_33), .Y(n_731) );
INVx1_ASAP7_75t_L g911 ( .A(n_34), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g924 ( .A1(n_34), .A2(n_211), .B1(n_549), .B2(n_692), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_35), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_36), .Y(n_1026) );
INVx1_ASAP7_75t_L g659 ( .A(n_37), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_37), .A2(n_40), .B1(n_704), .B2(n_705), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g1461 ( .A1(n_38), .A2(n_100), .B1(n_805), .B2(n_1266), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_38), .A2(n_100), .B1(n_1211), .B2(n_1282), .Y(n_1470) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_39), .Y(n_531) );
INVx1_ASAP7_75t_L g661 ( .A(n_40), .Y(n_661) );
INVx1_ASAP7_75t_L g1294 ( .A(n_41), .Y(n_1294) );
INVx1_ASAP7_75t_L g978 ( .A(n_42), .Y(n_978) );
INVx1_ASAP7_75t_L g1194 ( .A(n_43), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_43), .A2(n_196), .B1(n_805), .B2(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1382 ( .A(n_44), .Y(n_1382) );
AOI22xp33_ASAP7_75t_SL g1417 ( .A1(n_44), .A2(n_170), .B1(n_549), .B2(n_692), .Y(n_1417) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_45), .Y(n_632) );
INVx1_ASAP7_75t_L g585 ( .A(n_46), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_46), .A2(n_199), .B1(n_478), .B2(n_483), .Y(n_634) );
INVxp33_ASAP7_75t_L g1781 ( .A(n_47), .Y(n_1781) );
AOI221xp5_ASAP7_75t_L g1829 ( .A1(n_47), .A2(n_98), .B1(n_779), .B2(n_878), .C(n_1830), .Y(n_1829) );
AOI22xp33_ASAP7_75t_SL g1796 ( .A1(n_48), .A2(n_174), .B1(n_757), .B2(n_1797), .Y(n_1796) );
AOI22xp33_ASAP7_75t_L g1843 ( .A1(n_48), .A2(n_174), .B1(n_1511), .B2(n_1844), .Y(n_1843) );
INVx1_ASAP7_75t_L g1487 ( .A(n_49), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_50), .A2(n_95), .B1(n_870), .B2(n_1314), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_50), .A2(n_95), .B1(n_954), .B2(n_1273), .Y(n_1324) );
XNOR2xp5_ASAP7_75t_L g561 ( .A(n_51), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g1522 ( .A(n_52), .Y(n_1522) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_53), .A2(n_250), .B1(n_805), .B2(n_806), .C(n_807), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_53), .A2(n_250), .B1(n_549), .B2(n_692), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g1563 ( .A1(n_54), .A2(n_168), .B1(n_1564), .B2(n_1567), .Y(n_1563) );
INVx1_ASAP7_75t_L g663 ( .A(n_55), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_56), .A2(n_242), .B1(n_1226), .B2(n_1266), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_56), .A2(n_242), .B1(n_1211), .B2(n_1273), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1657 ( .A1(n_57), .A2(n_225), .B1(n_1551), .B2(n_1617), .Y(n_1657) );
INVxp33_ASAP7_75t_L g1458 ( .A(n_58), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_58), .A2(n_306), .B1(n_882), .B2(n_1008), .Y(n_1472) );
AOI22xp33_ASAP7_75t_SL g1799 ( .A1(n_59), .A2(n_330), .B1(n_1800), .B2(n_1801), .Y(n_1799) );
AOI221xp5_ASAP7_75t_L g1837 ( .A1(n_59), .A2(n_330), .B1(n_1838), .B2(n_1839), .C(n_1841), .Y(n_1837) );
INVxp67_ASAP7_75t_SL g1497 ( .A(n_60), .Y(n_1497) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_60), .A2(n_304), .B1(n_1362), .B2(n_1366), .Y(n_1505) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_61), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_62), .A2(n_207), .B1(n_678), .B2(n_827), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_62), .A2(n_207), .B1(n_672), .B2(n_674), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_63), .A2(n_138), .B1(n_1564), .B2(n_1567), .Y(n_1573) );
AO221x2_ASAP7_75t_L g1581 ( .A1(n_64), .A2(n_263), .B1(n_1557), .B2(n_1575), .C(n_1582), .Y(n_1581) );
CKINVDCx16_ASAP7_75t_R g1558 ( .A(n_65), .Y(n_1558) );
AOI22xp33_ASAP7_75t_SL g1802 ( .A1(n_66), .A2(n_134), .B1(n_1797), .B2(n_1800), .Y(n_1802) );
INVxp67_ASAP7_75t_SL g1817 ( .A(n_66), .Y(n_1817) );
AOI22xp5_ASAP7_75t_SL g1594 ( .A1(n_67), .A2(n_245), .B1(n_1551), .B2(n_1557), .Y(n_1594) );
INVxp33_ASAP7_75t_SL g1494 ( .A(n_68), .Y(n_1494) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_69), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_69), .A2(n_83), .B1(n_549), .B2(n_785), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_70), .A2(n_120), .B1(n_478), .B2(n_483), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_70), .A2(n_111), .B1(n_1068), .B2(n_1069), .Y(n_1067) );
INVxp67_ASAP7_75t_SL g1876 ( .A(n_71), .Y(n_1876) );
AOI22xp33_ASAP7_75t_L g1887 ( .A1(n_71), .A2(n_230), .B1(n_766), .B2(n_806), .Y(n_1887) );
INVx1_ASAP7_75t_L g820 ( .A(n_72), .Y(n_820) );
INVx1_ASAP7_75t_L g842 ( .A(n_73), .Y(n_842) );
INVx1_ASAP7_75t_L g853 ( .A(n_74), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_74), .A2(n_266), .B1(n_790), .B2(n_882), .Y(n_881) );
OAI211xp5_ASAP7_75t_L g796 ( .A1(n_75), .A2(n_420), .B(n_797), .C(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g814 ( .A(n_75), .Y(n_814) );
INVxp33_ASAP7_75t_SL g1259 ( .A(n_76), .Y(n_1259) );
AO22x2_ASAP7_75t_L g1238 ( .A1(n_77), .A2(n_1239), .B1(n_1284), .B2(n_1285), .Y(n_1238) );
CKINVDCx14_ASAP7_75t_R g1284 ( .A(n_77), .Y(n_1284) );
INVx1_ASAP7_75t_L g1385 ( .A(n_78), .Y(n_1385) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_78), .A2(n_187), .B1(n_590), .B2(n_1323), .Y(n_1416) );
OAI211xp5_ASAP7_75t_L g1422 ( .A1(n_78), .A2(n_474), .B(n_1423), .C(n_1424), .Y(n_1422) );
CKINVDCx5p33_ASAP7_75t_R g1193 ( .A(n_79), .Y(n_1193) );
INVx1_ASAP7_75t_L g1087 ( .A(n_80), .Y(n_1087) );
INVx1_ASAP7_75t_L g1397 ( .A(n_81), .Y(n_1397) );
OAI211xp5_ASAP7_75t_L g1428 ( .A1(n_81), .A2(n_420), .B(n_1429), .C(n_1430), .Y(n_1428) );
INVx1_ASAP7_75t_L g1081 ( .A(n_82), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_82), .A2(n_176), .B1(n_745), .B2(n_1103), .Y(n_1110) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_83), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g1803 ( .A1(n_84), .A2(n_121), .B1(n_757), .B2(n_1801), .Y(n_1803) );
INVxp67_ASAP7_75t_L g1836 ( .A(n_84), .Y(n_1836) );
INVx1_ASAP7_75t_L g1246 ( .A(n_85), .Y(n_1246) );
INVx1_ASAP7_75t_L g975 ( .A(n_86), .Y(n_975) );
INVx1_ASAP7_75t_L g1138 ( .A(n_87), .Y(n_1138) );
INVx1_ASAP7_75t_L g1394 ( .A(n_88), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_88), .A2(n_345), .B1(n_870), .B2(n_1407), .Y(n_1406) );
AO22x2_ASAP7_75t_L g1019 ( .A1(n_90), .A2(n_1020), .B1(n_1021), .B2(n_1071), .Y(n_1019) );
INVxp67_ASAP7_75t_L g1071 ( .A(n_90), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1655 ( .A1(n_90), .A2(n_221), .B1(n_1564), .B2(n_1656), .Y(n_1655) );
CKINVDCx5p33_ASAP7_75t_R g961 ( .A(n_91), .Y(n_961) );
INVxp33_ASAP7_75t_SL g1095 ( .A(n_92), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_92), .A2(n_161), .B1(n_496), .B2(n_1049), .Y(n_1116) );
INVxp67_ASAP7_75t_SL g1250 ( .A(n_93), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_93), .A2(n_319), .B1(n_522), .B2(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1202 ( .A(n_94), .Y(n_1202) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_96), .A2(n_275), .B1(n_522), .B2(n_524), .C(n_528), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_96), .A2(n_275), .B1(n_548), .B2(n_549), .Y(n_547) );
CKINVDCx14_ASAP7_75t_R g1583 ( .A(n_97), .Y(n_1583) );
INVxp33_ASAP7_75t_SL g1792 ( .A(n_98), .Y(n_1792) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_99), .A2(n_257), .B1(n_478), .B2(n_483), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_99), .A2(n_257), .B1(n_548), .B2(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g438 ( .A(n_101), .Y(n_438) );
BUFx2_ASAP7_75t_L g490 ( .A(n_101), .Y(n_490) );
INVx1_ASAP7_75t_L g518 ( .A(n_101), .Y(n_518) );
OR2x2_ASAP7_75t_L g1774 ( .A(n_101), .B(n_1775), .Y(n_1774) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_102), .A2(n_199), .B1(n_587), .B2(n_590), .Y(n_586) );
OAI211xp5_ASAP7_75t_L g628 ( .A1(n_102), .A2(n_474), .B(n_629), .C(n_630), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_103), .A2(n_262), .B1(n_1277), .B2(n_1303), .Y(n_1352) );
INVxp67_ASAP7_75t_SL g1371 ( .A(n_103), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_104), .A2(n_365), .B1(n_1211), .B2(n_1358), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_104), .A2(n_365), .B1(n_1362), .B2(n_1366), .Y(n_1365) );
INVxp67_ASAP7_75t_SL g1243 ( .A(n_105), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_105), .A2(n_323), .B1(n_733), .B2(n_855), .Y(n_1256) );
AO22x2_ASAP7_75t_L g1180 ( .A1(n_106), .A2(n_1181), .B1(n_1182), .B2(n_1235), .Y(n_1180) );
INVx1_ASAP7_75t_L g1235 ( .A(n_106), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_107), .A2(n_297), .B1(n_1172), .B2(n_1303), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_107), .A2(n_297), .B1(n_702), .B2(n_1159), .Y(n_1368) );
INVx1_ASAP7_75t_L g893 ( .A(n_108), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_108), .A2(n_368), .B1(n_498), .B2(n_504), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_109), .A2(n_332), .B1(n_757), .B2(n_760), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_109), .A2(n_332), .B1(n_689), .B2(n_774), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_110), .Y(n_464) );
INVx1_ASAP7_75t_L g1030 ( .A(n_111), .Y(n_1030) );
INVx1_ASAP7_75t_L g1486 ( .A(n_112), .Y(n_1486) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_113), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_114), .A2(n_367), .B1(n_688), .B2(n_689), .Y(n_687) );
INVxp33_ASAP7_75t_L g712 ( .A(n_114), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_115), .A2(n_261), .B1(n_396), .B2(n_409), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_115), .A2(n_261), .B1(n_496), .B2(n_767), .C(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g623 ( .A(n_116), .Y(n_623) );
OAI211xp5_ASAP7_75t_SL g638 ( .A1(n_116), .A2(n_639), .B(n_641), .C(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g1009 ( .A(n_117), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_118), .A2(n_126), .B1(n_847), .B2(n_898), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_118), .A2(n_126), .B1(n_855), .B2(n_906), .Y(n_905) );
INVxp67_ASAP7_75t_SL g1132 ( .A(n_119), .Y(n_1132) );
AOI22xp33_ASAP7_75t_SL g1155 ( .A1(n_119), .A2(n_249), .B1(n_805), .B2(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1066 ( .A(n_120), .Y(n_1066) );
INVxp33_ASAP7_75t_L g1849 ( .A(n_121), .Y(n_1849) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_122), .A2(n_148), .B1(n_1106), .B2(n_1109), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_122), .A2(n_148), .B1(n_1049), .B2(n_1082), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_123), .A2(n_281), .B1(n_1008), .B2(n_1107), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_123), .A2(n_281), .B1(n_1232), .B2(n_1233), .Y(n_1231) );
INVx1_ASAP7_75t_L g808 ( .A(n_124), .Y(n_808) );
INVx1_ASAP7_75t_L g1002 ( .A(n_125), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1404 ( .A1(n_127), .A2(n_162), .B1(n_698), .B2(n_866), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_127), .A2(n_162), .B1(n_790), .B2(n_882), .Y(n_1411) );
INVx1_ASAP7_75t_L g1789 ( .A(n_128), .Y(n_1789) );
INVxp33_ASAP7_75t_SL g1078 ( .A(n_129), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_129), .A2(n_178), .B1(n_1102), .B2(n_1112), .Y(n_1111) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_130), .Y(n_529) );
INVx1_ASAP7_75t_L g987 ( .A(n_131), .Y(n_987) );
OAI22xp33_ASAP7_75t_SL g1015 ( .A1(n_131), .A2(n_232), .B1(n_466), .B2(n_478), .Y(n_1015) );
AO22x2_ASAP7_75t_L g645 ( .A1(n_132), .A2(n_646), .B1(n_715), .B2(n_716), .Y(n_645) );
INVx1_ASAP7_75t_L g715 ( .A(n_132), .Y(n_715) );
INVx1_ASAP7_75t_L g801 ( .A(n_133), .Y(n_801) );
INVxp33_ASAP7_75t_L g1852 ( .A(n_134), .Y(n_1852) );
INVxp33_ASAP7_75t_SL g1455 ( .A(n_135), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_135), .A2(n_233), .B1(n_1212), .B2(n_1474), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1892 ( .A1(n_136), .A2(n_270), .B1(n_774), .B2(n_1303), .Y(n_1892) );
INVxp67_ASAP7_75t_SL g1897 ( .A(n_136), .Y(n_1897) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_137), .A2(n_218), .B1(n_1176), .B2(n_1212), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_137), .A2(n_218), .B1(n_1226), .B2(n_1228), .Y(n_1225) );
XOR2xp5_ASAP7_75t_L g926 ( .A(n_138), .B(n_927), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_139), .A2(n_327), .B1(n_548), .B2(n_549), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_139), .A2(n_327), .B1(n_504), .B2(n_676), .Y(n_696) );
INVx1_ASAP7_75t_L g1300 ( .A(n_140), .Y(n_1300) );
INVx1_ASAP7_75t_L g1880 ( .A(n_141), .Y(n_1880) );
OAI22xp5_ASAP7_75t_L g1898 ( .A1(n_141), .A2(n_321), .B1(n_704), .B2(n_705), .Y(n_1898) );
INVxp33_ASAP7_75t_L g739 ( .A(n_142), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_142), .A2(n_198), .B1(n_757), .B2(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_SL g1462 ( .A1(n_143), .A2(n_317), .B1(n_1222), .B2(n_1224), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_143), .A2(n_317), .B1(n_1008), .B2(n_1277), .Y(n_1469) );
INVxp33_ASAP7_75t_SL g1442 ( .A(n_144), .Y(n_1442) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_144), .A2(n_359), .B1(n_1226), .B2(n_1465), .Y(n_1464) );
INVxp67_ASAP7_75t_SL g1776 ( .A(n_145), .Y(n_1776) );
OAI22xp33_ASAP7_75t_L g1821 ( .A1(n_145), .A2(n_181), .B1(n_1822), .B2(n_1826), .Y(n_1821) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_146), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_146), .A2(n_229), .B1(n_678), .B2(n_682), .Y(n_677) );
INVx1_ASAP7_75t_L g998 ( .A(n_147), .Y(n_998) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_147), .A2(n_154), .B1(n_386), .B2(n_396), .Y(n_1004) );
INVx1_ASAP7_75t_L g726 ( .A(n_149), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_150), .A2(n_224), .B1(n_574), .B2(n_576), .Y(n_573) );
INVx1_ASAP7_75t_L g604 ( .A(n_150), .Y(n_604) );
INVxp33_ASAP7_75t_L g1310 ( .A(n_151), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_151), .A2(n_342), .B1(n_698), .B2(n_760), .Y(n_1320) );
INVx1_ASAP7_75t_L g940 ( .A(n_152), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_152), .A2(n_307), .B1(n_396), .B2(n_409), .Y(n_963) );
AOI22xp5_ASAP7_75t_L g1479 ( .A1(n_153), .A2(n_1480), .B1(n_1516), .B2(n_1517), .Y(n_1479) );
INVxp67_ASAP7_75t_L g1516 ( .A(n_153), .Y(n_1516) );
AOI22xp5_ASAP7_75t_SL g1593 ( .A1(n_153), .A2(n_177), .B1(n_1564), .B2(n_1567), .Y(n_1593) );
INVx1_ASAP7_75t_L g1001 ( .A(n_154), .Y(n_1001) );
INVxp33_ASAP7_75t_SL g653 ( .A(n_155), .Y(n_653) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_155), .A2(n_337), .B1(n_504), .B2(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1541 ( .A(n_156), .Y(n_1541) );
INVxp33_ASAP7_75t_SL g1128 ( .A(n_157), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_157), .A2(n_313), .B1(n_443), .B2(n_1159), .Y(n_1158) );
INVxp33_ASAP7_75t_SL g1872 ( .A(n_158), .Y(n_1872) );
AOI22xp33_ASAP7_75t_L g1888 ( .A1(n_158), .A2(n_203), .B1(n_757), .B2(n_1145), .Y(n_1888) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_159), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_160), .A2(n_256), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_160), .A2(n_256), .B1(n_590), .B2(n_876), .Y(n_875) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_161), .Y(n_1097) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_163), .Y(n_729) );
INVx1_ASAP7_75t_L g1448 ( .A(n_164), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1453 ( .A1(n_164), .A2(n_300), .B1(n_705), .B2(n_733), .Y(n_1453) );
OAI211xp5_ASAP7_75t_L g1034 ( .A1(n_165), .A2(n_420), .B(n_639), .C(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1055 ( .A(n_165), .Y(n_1055) );
CKINVDCx16_ASAP7_75t_R g1548 ( .A(n_166), .Y(n_1548) );
INVx1_ASAP7_75t_L g951 ( .A(n_167), .Y(n_951) );
OAI22xp33_ASAP7_75t_SL g969 ( .A1(n_167), .A2(n_184), .B1(n_466), .B2(n_478), .Y(n_969) );
INVxp33_ASAP7_75t_SL g1340 ( .A(n_169), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_169), .A2(n_182), .B1(n_702), .B2(n_758), .Y(n_1363) );
INVx1_ASAP7_75t_L g1383 ( .A(n_170), .Y(n_1383) );
INVx1_ASAP7_75t_L g1542 ( .A(n_171), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_171), .B(n_1540), .Y(n_1547) );
INVxp33_ASAP7_75t_SL g1253 ( .A(n_172), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_172), .A2(n_346), .B1(n_656), .B2(n_1277), .Y(n_1276) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_175), .Y(n_1387) );
INVxp67_ASAP7_75t_SL g1079 ( .A(n_176), .Y(n_1079) );
INVxp33_ASAP7_75t_SL g1086 ( .A(n_178), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_179), .A2(n_190), .B1(n_386), .B2(n_396), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_179), .A2(n_324), .B1(n_496), .B2(n_502), .C(n_505), .Y(n_495) );
INVx2_ASAP7_75t_L g448 ( .A(n_180), .Y(n_448) );
INVxp67_ASAP7_75t_SL g1778 ( .A(n_181), .Y(n_1778) );
INVxp67_ASAP7_75t_SL g1343 ( .A(n_182), .Y(n_1343) );
INVxp33_ASAP7_75t_L g1441 ( .A(n_183), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_183), .A2(n_350), .B1(n_682), .B2(n_1232), .Y(n_1467) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_184), .A2(n_299), .B1(n_558), .B2(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g393 ( .A(n_186), .Y(n_393) );
BUFx3_ASAP7_75t_L g399 ( .A(n_186), .Y(n_399) );
INVx1_ASAP7_75t_L g1389 ( .A(n_187), .Y(n_1389) );
INVx1_ASAP7_75t_L g1144 ( .A(n_188), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_188), .A2(n_265), .B1(n_1172), .B2(n_1174), .Y(n_1171) );
INVx1_ASAP7_75t_L g1137 ( .A(n_189), .Y(n_1137) );
INVx1_ASAP7_75t_L g506 ( .A(n_190), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_191), .A2(n_252), .B1(n_504), .B2(n_676), .Y(n_914) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_191), .A2(n_252), .B1(n_558), .B2(n_692), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_192), .A2(n_356), .B1(n_386), .B2(n_396), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_192), .A2(n_356), .B1(n_496), .B2(n_1049), .C(n_1052), .Y(n_1048) );
AOI22xp33_ASAP7_75t_SL g1153 ( .A1(n_193), .A2(n_371), .B1(n_443), .B2(n_758), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_193), .A2(n_371), .B1(n_746), .B2(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g889 ( .A(n_194), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_194), .A2(n_326), .B1(n_678), .B2(n_827), .Y(n_918) );
INVxp33_ASAP7_75t_L g735 ( .A(n_195), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_195), .A2(n_255), .B1(n_774), .B2(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g1191 ( .A(n_196), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1886 ( .A1(n_197), .A2(n_248), .B1(n_496), .B2(n_502), .Y(n_1886) );
AOI22xp33_ASAP7_75t_L g1890 ( .A1(n_197), .A2(n_248), .B1(n_1176), .B2(n_1511), .Y(n_1890) );
INVx1_ASAP7_75t_L g744 ( .A(n_198), .Y(n_744) );
INVx1_ASAP7_75t_L g1131 ( .A(n_200), .Y(n_1131) );
INVx1_ASAP7_75t_L g1190 ( .A(n_201), .Y(n_1190) );
AOI22xp33_ASAP7_75t_SL g1884 ( .A1(n_202), .A2(n_369), .B1(n_757), .B2(n_1885), .Y(n_1884) );
AOI22xp33_ASAP7_75t_SL g1891 ( .A1(n_202), .A2(n_369), .B1(n_746), .B2(n_1164), .Y(n_1891) );
INVx1_ASAP7_75t_L g1878 ( .A(n_203), .Y(n_1878) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_204), .A2(n_302), .B1(n_1102), .B2(n_1103), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_204), .A2(n_302), .B1(n_496), .B2(n_1043), .Y(n_1115) );
INVx1_ASAP7_75t_L g1295 ( .A(n_205), .Y(n_1295) );
XNOR2xp5_ASAP7_75t_L g382 ( .A(n_206), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g988 ( .A(n_208), .Y(n_988) );
OAI211xp5_ASAP7_75t_SL g1013 ( .A1(n_208), .A2(n_474), .B(n_967), .C(n_1014), .Y(n_1013) );
AO22x2_ASAP7_75t_L g1287 ( .A1(n_209), .A2(n_1288), .B1(n_1328), .B2(n_1329), .Y(n_1287) );
INVx1_ASAP7_75t_L g1328 ( .A(n_209), .Y(n_1328) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_210), .A2(n_303), .B1(n_386), .B2(n_401), .Y(n_795) );
INVx1_ASAP7_75t_L g829 ( .A(n_210), .Y(n_829) );
INVx1_ASAP7_75t_L g909 ( .A(n_211), .Y(n_909) );
INVx1_ASAP7_75t_L g436 ( .A(n_212), .Y(n_436) );
INVx1_ASAP7_75t_L g1813 ( .A(n_212), .Y(n_1813) );
INVxp33_ASAP7_75t_SL g1141 ( .A(n_213), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_213), .A2(n_247), .B1(n_576), .B2(n_1176), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_214), .A2(n_217), .B1(n_702), .B2(n_758), .Y(n_1503) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_214), .A2(n_217), .B1(n_1277), .B2(n_1303), .Y(n_1508) );
INVx1_ASAP7_75t_L g1785 ( .A(n_215), .Y(n_1785) );
INVxp67_ASAP7_75t_L g860 ( .A(n_216), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_216), .A2(n_309), .B1(n_549), .B2(n_692), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g1620 ( .A(n_219), .Y(n_1620) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_220), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_220), .A2(n_349), .B1(n_558), .B2(n_589), .Y(n_949) );
INVx1_ASAP7_75t_L g615 ( .A(n_222), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_222), .A2(n_226), .B1(n_386), .B2(n_396), .Y(n_636) );
INVx1_ASAP7_75t_L g1197 ( .A(n_223), .Y(n_1197) );
INVx1_ASAP7_75t_L g598 ( .A(n_224), .Y(n_598) );
INVx1_ASAP7_75t_L g611 ( .A(n_226), .Y(n_611) );
CKINVDCx14_ASAP7_75t_R g792 ( .A(n_227), .Y(n_792) );
INVx1_ASAP7_75t_L g800 ( .A(n_228), .Y(n_800) );
INVxp33_ASAP7_75t_SL g649 ( .A(n_229), .Y(n_649) );
INVxp33_ASAP7_75t_SL g1873 ( .A(n_230), .Y(n_1873) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_231), .A2(n_324), .B1(n_401), .B2(n_409), .Y(n_400) );
INVx1_ASAP7_75t_L g469 ( .A(n_231), .Y(n_469) );
INVx1_ASAP7_75t_L g990 ( .A(n_232), .Y(n_990) );
INVxp67_ASAP7_75t_SL g1456 ( .A(n_233), .Y(n_1456) );
INVxp67_ASAP7_75t_SL g1346 ( .A(n_234), .Y(n_1346) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_235), .Y(n_1046) );
INVxp33_ASAP7_75t_L g1291 ( .A(n_236), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_236), .A2(n_333), .B1(n_584), .B2(n_954), .Y(n_1327) );
INVxp33_ASAP7_75t_L g1309 ( .A(n_237), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_237), .A2(n_293), .B1(n_1219), .B2(n_1319), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_238), .A2(n_362), .B1(n_760), .B2(n_865), .Y(n_1316) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_238), .A2(n_362), .B1(n_674), .B2(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g932 ( .A(n_239), .Y(n_932) );
INVx1_ASAP7_75t_L g1875 ( .A(n_240), .Y(n_1875) );
INVx1_ASAP7_75t_L g1201 ( .A(n_241), .Y(n_1201) );
INVx1_ASAP7_75t_L g1348 ( .A(n_243), .Y(n_1348) );
INVxp33_ASAP7_75t_SL g1249 ( .A(n_244), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_244), .A2(n_258), .B1(n_702), .B2(n_1232), .Y(n_1268) );
INVxp33_ASAP7_75t_SL g1142 ( .A(n_247), .Y(n_1142) );
INVxp33_ASAP7_75t_SL g1129 ( .A(n_249), .Y(n_1129) );
INVx1_ASAP7_75t_L g810 ( .A(n_251), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_253), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_254), .A2(n_259), .B1(n_401), .B2(n_409), .Y(n_1037) );
INVx1_ASAP7_75t_L g1053 ( .A(n_254), .Y(n_1053) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_255), .Y(n_730) );
INVx1_ASAP7_75t_L g1242 ( .A(n_258), .Y(n_1242) );
INVx1_ASAP7_75t_L g1031 ( .A(n_259), .Y(n_1031) );
INVx1_ASAP7_75t_L g1093 ( .A(n_260), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_260), .A2(n_308), .B1(n_682), .B2(n_806), .Y(n_1117) );
INVxp67_ASAP7_75t_SL g1374 ( .A(n_262), .Y(n_1374) );
INVx1_ASAP7_75t_L g991 ( .A(n_264), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_264), .A2(n_277), .B1(n_471), .B2(n_483), .Y(n_1012) );
INVxp33_ASAP7_75t_SL g1147 ( .A(n_265), .Y(n_1147) );
INVxp33_ASAP7_75t_L g857 ( .A(n_266), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_267), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g1543 ( .A(n_268), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1862 ( .A1(n_268), .A2(n_1863), .B1(n_1904), .B2(n_1908), .Y(n_1862) );
INVx1_ASAP7_75t_L g1083 ( .A(n_269), .Y(n_1083) );
INVxp33_ASAP7_75t_L g1903 ( .A(n_270), .Y(n_1903) );
INVx1_ASAP7_75t_L g395 ( .A(n_271), .Y(n_395) );
BUFx3_ASAP7_75t_L g408 ( .A(n_271), .Y(n_408) );
INVx1_ASAP7_75t_L g821 ( .A(n_273), .Y(n_821) );
AO221x2_ASAP7_75t_L g1616 ( .A1(n_274), .A2(n_347), .B1(n_1617), .B2(n_1618), .C(n_1619), .Y(n_1616) );
INVx1_ASAP7_75t_L g582 ( .A(n_276), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_276), .A2(n_339), .B1(n_466), .B2(n_471), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_277), .A2(n_286), .B1(n_401), .B2(n_409), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1574 ( .A1(n_278), .A2(n_279), .B1(n_1557), .B2(n_1575), .Y(n_1574) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_280), .Y(n_493) );
INVx1_ASAP7_75t_L g520 ( .A(n_280), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g1775 ( .A(n_280), .B(n_354), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1784 ( .A(n_280), .B(n_462), .Y(n_1784) );
AOI221xp5_ASAP7_75t_SL g1042 ( .A1(n_282), .A2(n_290), .B1(n_1043), .B2(n_1044), .C(n_1045), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_282), .A2(n_290), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
AO22x2_ASAP7_75t_L g1124 ( .A1(n_283), .A2(n_1125), .B1(n_1178), .B2(n_1179), .Y(n_1124) );
INVx1_ASAP7_75t_L g1178 ( .A(n_283), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_284), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_285), .A2(n_328), .B1(n_902), .B2(n_1232), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_285), .A2(n_328), .B1(n_1008), .B2(n_1107), .Y(n_1275) );
INVx1_ASAP7_75t_L g999 ( .A(n_286), .Y(n_999) );
XNOR2xp5_ASAP7_75t_L g970 ( .A(n_287), .B(n_971), .Y(n_970) );
INVx2_ASAP7_75t_L g390 ( .A(n_288), .Y(n_390) );
OR2x2_ASAP7_75t_L g1820 ( .A(n_288), .B(n_1813), .Y(n_1820) );
INVx1_ASAP7_75t_L g835 ( .A(n_289), .Y(n_835) );
INVx1_ASAP7_75t_L g1204 ( .A(n_291), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_291), .A2(n_296), .B1(n_1107), .B2(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1444 ( .A(n_292), .Y(n_1444) );
INVxp33_ASAP7_75t_L g1307 ( .A(n_293), .Y(n_1307) );
INVx1_ASAP7_75t_L g1010 ( .A(n_294), .Y(n_1010) );
INVxp33_ASAP7_75t_SL g1483 ( .A(n_295), .Y(n_1483) );
AOI22xp33_ASAP7_75t_SL g1514 ( .A1(n_295), .A2(n_298), .B1(n_1354), .B2(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1200 ( .A(n_296), .Y(n_1200) );
INVxp33_ASAP7_75t_SL g1484 ( .A(n_298), .Y(n_1484) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_299), .A2(n_343), .B1(n_471), .B2(n_483), .Y(n_965) );
INVx1_ASAP7_75t_L g1449 ( .A(n_300), .Y(n_1449) );
CKINVDCx5p33_ASAP7_75t_R g1047 ( .A(n_301), .Y(n_1047) );
INVx1_ASAP7_75t_L g813 ( .A(n_303), .Y(n_813) );
INVxp33_ASAP7_75t_SL g1495 ( .A(n_304), .Y(n_1495) );
AOI22xp5_ASAP7_75t_SL g1569 ( .A1(n_305), .A2(n_311), .B1(n_1551), .B2(n_1557), .Y(n_1569) );
INVxp67_ASAP7_75t_SL g1452 ( .A(n_306), .Y(n_1452) );
INVx1_ASAP7_75t_L g938 ( .A(n_307), .Y(n_938) );
INVxp33_ASAP7_75t_SL g1091 ( .A(n_308), .Y(n_1091) );
INVx1_ASAP7_75t_L g858 ( .A(n_309), .Y(n_858) );
AO22x2_ASAP7_75t_L g1378 ( .A1(n_312), .A2(n_1379), .B1(n_1418), .B2(n_1419), .Y(n_1378) );
INVxp67_ASAP7_75t_L g1418 ( .A(n_312), .Y(n_1418) );
INVx1_ASAP7_75t_L g1134 ( .A(n_313), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_315), .A2(n_353), .B1(n_805), .B2(n_1151), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_315), .A2(n_353), .B1(n_1167), .B2(n_1169), .Y(n_1166) );
INVx1_ASAP7_75t_L g952 ( .A(n_316), .Y(n_952) );
OAI211xp5_ASAP7_75t_SL g966 ( .A1(n_316), .A2(n_474), .B(n_967), .C(n_968), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_318), .A2(n_351), .B1(n_844), .B2(n_847), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_318), .A2(n_351), .B1(n_704), .B2(n_855), .Y(n_854) );
INVxp67_ASAP7_75t_SL g1247 ( .A(n_319), .Y(n_1247) );
INVxp33_ASAP7_75t_L g708 ( .A(n_320), .Y(n_708) );
INVx1_ASAP7_75t_L g1881 ( .A(n_321), .Y(n_1881) );
INVx1_ASAP7_75t_L g908 ( .A(n_322), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_322), .A2(n_358), .B1(n_672), .B2(n_790), .Y(n_923) );
INVxp67_ASAP7_75t_SL g1244 ( .A(n_323), .Y(n_1244) );
CKINVDCx5p33_ASAP7_75t_R g1390 ( .A(n_325), .Y(n_1390) );
INVx1_ASAP7_75t_L g896 ( .A(n_326), .Y(n_896) );
INVx1_ASAP7_75t_L g722 ( .A(n_329), .Y(n_722) );
INVx1_ASAP7_75t_L g1488 ( .A(n_331), .Y(n_1488) );
INVxp33_ASAP7_75t_L g1292 ( .A(n_333), .Y(n_1292) );
INVx1_ASAP7_75t_L g981 ( .A(n_334), .Y(n_981) );
INVx1_ASAP7_75t_L g1297 ( .A(n_335), .Y(n_1297) );
INVxp67_ASAP7_75t_SL g740 ( .A(n_336), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_336), .A2(n_357), .B1(n_766), .B2(n_767), .Y(n_765) );
INVxp33_ASAP7_75t_SL g664 ( .A(n_337), .Y(n_664) );
HB1xp67_ASAP7_75t_L g1524 ( .A(n_338), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_338), .B(n_1522), .Y(n_1538) );
AND3x2_ASAP7_75t_L g1554 ( .A(n_338), .B(n_1522), .C(n_1541), .Y(n_1554) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_339), .A2(n_364), .B1(n_401), .B2(n_409), .Y(n_637) );
INVxp33_ASAP7_75t_SL g1341 ( .A(n_340), .Y(n_1341) );
INVx2_ASAP7_75t_L g450 ( .A(n_341), .Y(n_450) );
INVx1_ASAP7_75t_L g1305 ( .A(n_342), .Y(n_1305) );
INVx1_ASAP7_75t_L g1491 ( .A(n_344), .Y(n_1491) );
INVx1_ASAP7_75t_L g1399 ( .A(n_345), .Y(n_1399) );
INVxp67_ASAP7_75t_SL g1255 ( .A(n_346), .Y(n_1255) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_348), .Y(n_430) );
INVxp67_ASAP7_75t_SL g934 ( .A(n_349), .Y(n_934) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_350), .Y(n_1447) );
INVx1_ASAP7_75t_L g931 ( .A(n_352), .Y(n_931) );
INVx1_ASAP7_75t_L g453 ( .A(n_354), .Y(n_453) );
INVx2_ASAP7_75t_L g462 ( .A(n_354), .Y(n_462) );
XNOR2xp5_ASAP7_75t_L g885 ( .A(n_355), .B(n_886), .Y(n_885) );
INVxp67_ASAP7_75t_SL g742 ( .A(n_357), .Y(n_742) );
INVx1_ASAP7_75t_L g901 ( .A(n_358), .Y(n_901) );
INVxp33_ASAP7_75t_L g1445 ( .A(n_359), .Y(n_1445) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_360), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_361), .Y(n_433) );
AO22x2_ASAP7_75t_L g1073 ( .A1(n_363), .A2(n_1074), .B1(n_1075), .B2(n_1118), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_363), .Y(n_1074) );
INVx1_ASAP7_75t_L g620 ( .A(n_364), .Y(n_620) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_367), .Y(n_701) );
INVx1_ASAP7_75t_L g894 ( .A(n_368), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g1893 ( .A1(n_370), .A2(n_373), .B1(n_1065), .B2(n_1894), .Y(n_1893) );
INVxp33_ASAP7_75t_L g1900 ( .A(n_370), .Y(n_1900) );
INVx1_ASAP7_75t_L g944 ( .A(n_372), .Y(n_944) );
INVxp67_ASAP7_75t_SL g1901 ( .A(n_373), .Y(n_1901) );
AO22x1_ASAP7_75t_L g1436 ( .A1(n_374), .A2(n_1437), .B1(n_1438), .B2(n_1475), .Y(n_1436) );
INVxp67_ASAP7_75t_L g1437 ( .A(n_374), .Y(n_1437) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_1518), .B(n_1528), .Y(n_375) );
XNOR2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_1120), .Y(n_376) );
XNOR2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_718), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
XOR2x2_ASAP7_75t_SL g379 ( .A(n_380), .B(n_559), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND3x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_439), .C(n_494), .Y(n_383) );
OAI31xp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_400), .A3(n_415), .B(n_434), .Y(n_384) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_391), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x6_ASAP7_75t_L g397 ( .A(n_388), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
AND2x2_ASAP7_75t_L g798 ( .A(n_388), .B(n_674), .Y(n_798) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x6_ASAP7_75t_L g431 ( .A(n_389), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_390), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
AND2x2_ASAP7_75t_L g541 ( .A(n_390), .B(n_436), .Y(n_541) );
INVx2_ASAP7_75t_L g553 ( .A(n_390), .Y(n_553) );
INVx2_ASAP7_75t_L g544 ( .A(n_391), .Y(n_544) );
BUFx2_ASAP7_75t_L g568 ( .A(n_391), .Y(n_568) );
INVx1_ASAP7_75t_L g581 ( .A(n_391), .Y(n_581) );
INVx1_ASAP7_75t_L g983 ( .A(n_391), .Y(n_983) );
OR2x2_ASAP7_75t_L g1851 ( .A(n_391), .B(n_1820), .Y(n_1851) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
AND2x2_ASAP7_75t_L g419 ( .A(n_392), .B(n_394), .Y(n_419) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g414 ( .A(n_393), .B(n_408), .Y(n_414) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g398 ( .A(n_395), .B(n_399), .Y(n_398) );
CKINVDCx6p67_ASAP7_75t_R g396 ( .A(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_397), .A2(n_649), .B1(n_650), .B2(n_653), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_397), .A2(n_650), .B1(n_739), .B2(n_740), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_397), .A2(n_410), .B1(n_849), .B2(n_850), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_397), .A2(n_410), .B1(n_893), .B2(n_894), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_397), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_397), .A2(n_650), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_397), .A2(n_890), .B1(n_1190), .B2(n_1191), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_397), .A2(n_650), .B1(n_1249), .B2(n_1250), .Y(n_1248) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_397), .A2(n_890), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
AOI221xp5_ASAP7_75t_L g1339 ( .A1(n_397), .A2(n_421), .B1(n_650), .B2(n_1340), .C(n_1341), .Y(n_1339) );
AOI22xp5_ASAP7_75t_SL g1392 ( .A1(n_397), .A2(n_890), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_397), .A2(n_890), .B1(n_1441), .B2(n_1442), .Y(n_1440) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_397), .A2(n_650), .B1(n_1494), .B2(n_1495), .Y(n_1493) );
AOI22xp33_ASAP7_75t_L g1871 ( .A1(n_397), .A2(n_650), .B1(n_1872), .B2(n_1873), .Y(n_1871) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_398), .Y(n_548) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_398), .Y(n_589) );
BUFx3_ASAP7_75t_L g692 ( .A(n_398), .Y(n_692) );
INVx2_ASAP7_75t_SL g879 ( .A(n_398), .Y(n_879) );
BUFx6f_ASAP7_75t_L g954 ( .A(n_398), .Y(n_954) );
BUFx6f_ASAP7_75t_L g977 ( .A(n_398), .Y(n_977) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_398), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1474 ( .A(n_398), .Y(n_1474) );
BUFx2_ASAP7_75t_L g1510 ( .A(n_398), .Y(n_1510) );
BUFx2_ASAP7_75t_L g1838 ( .A(n_398), .Y(n_1838) );
INVx2_ASAP7_75t_L g406 ( .A(n_399), .Y(n_406) );
AND2x2_ASAP7_75t_L g424 ( .A(n_399), .B(n_408), .Y(n_424) );
INVx4_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_402), .A2(n_410), .B1(n_663), .B2(n_664), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_402), .A2(n_410), .B1(n_726), .B2(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_SL g838 ( .A1(n_402), .A2(n_650), .B1(n_839), .B2(n_840), .Y(n_838) );
AOI22xp5_ASAP7_75t_SL g888 ( .A1(n_402), .A2(n_889), .B1(n_890), .B2(n_891), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_402), .A2(n_410), .B1(n_1087), .B2(n_1091), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_402), .A2(n_410), .B1(n_1131), .B2(n_1132), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_402), .A2(n_410), .B1(n_1193), .B2(n_1194), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_402), .A2(n_410), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1306 ( .A1(n_402), .A2(n_410), .B1(n_421), .B2(n_1300), .C(n_1307), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_402), .A2(n_410), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
AOI22xp5_ASAP7_75t_L g1398 ( .A1(n_402), .A2(n_410), .B1(n_1390), .B2(n_1399), .Y(n_1398) );
AOI22xp33_ASAP7_75t_L g1443 ( .A1(n_402), .A2(n_410), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_402), .A2(n_410), .B1(n_1491), .B2(n_1497), .Y(n_1496) );
AOI22xp33_ASAP7_75t_L g1874 ( .A1(n_402), .A2(n_410), .B1(n_1875), .B2(n_1876), .Y(n_1874) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
AND2x4_ASAP7_75t_L g426 ( .A(n_403), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_SL g660 ( .A(n_403), .B(n_427), .Y(n_660) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx6_ASAP7_75t_L g652 ( .A(n_405), .Y(n_652) );
INVx2_ASAP7_75t_L g673 ( .A(n_405), .Y(n_673) );
BUFx2_ASAP7_75t_L g882 ( .A(n_405), .Y(n_882) );
AND2x2_ASAP7_75t_L g1810 ( .A(n_405), .B(n_1811), .Y(n_1810) );
AND2x4_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
INVx1_ASAP7_75t_L g429 ( .A(n_407), .Y(n_429) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x6_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
AND2x4_ASAP7_75t_L g650 ( .A(n_411), .B(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_L g890 ( .A(n_411), .B(n_651), .Y(n_890) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g845 ( .A(n_412), .B(n_846), .Y(n_845) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_413), .Y(n_549) );
INVx2_ASAP7_75t_L g577 ( .A(n_413), .Y(n_577) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_413), .Y(n_584) );
INVx1_ASAP7_75t_L g1274 ( .A(n_413), .Y(n_1274) );
INVx1_ASAP7_75t_L g1283 ( .A(n_413), .Y(n_1283) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_414), .Y(n_558) );
INVx2_ASAP7_75t_L g695 ( .A(n_414), .Y(n_695) );
INVx1_ASAP7_75t_L g780 ( .A(n_414), .Y(n_780) );
INVx1_ASAP7_75t_L g1414 ( .A(n_414), .Y(n_1414) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_417), .A2(n_543), .B1(n_951), .B2(n_952), .C(n_953), .Y(n_950) );
INVx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g546 ( .A(n_419), .Y(n_546) );
BUFx4f_ASAP7_75t_L g556 ( .A(n_419), .Y(n_556) );
INVx1_ASAP7_75t_L g571 ( .A(n_419), .Y(n_571) );
INVx1_ASAP7_75t_L g1188 ( .A(n_419), .Y(n_1188) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_420), .B(n_648), .C(n_654), .D(n_662), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g957 ( .A(n_420), .B(n_958), .Y(n_957) );
NAND2xp5_ASAP7_75t_SL g1006 ( .A(n_420), .B(n_1007), .Y(n_1006) );
NAND4xp25_ASAP7_75t_SL g1240 ( .A(n_420), .B(n_1241), .C(n_1245), .D(n_1248), .Y(n_1240) );
NAND4xp25_ASAP7_75t_SL g1492 ( .A(n_420), .B(n_1493), .C(n_1496), .D(n_1498), .Y(n_1492) );
CKINVDCx8_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
INVx5_ASAP7_75t_L g641 ( .A(n_421), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_421), .B(n_1185), .Y(n_1184) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g591 ( .A(n_423), .Y(n_591) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_423), .Y(n_674) );
INVx2_ASAP7_75t_L g690 ( .A(n_423), .Y(n_690) );
BUFx6f_ASAP7_75t_L g1304 ( .A(n_423), .Y(n_1304) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_424), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_430), .B1(n_431), .B2(n_433), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_426), .A2(n_431), .B1(n_631), .B2(n_632), .Y(n_642) );
BUFx4f_ASAP7_75t_L g747 ( .A(n_426), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_426), .A2(n_431), .B1(n_800), .B2(n_801), .Y(n_799) );
AOI222xp33_ASAP7_75t_L g1241 ( .A1(n_426), .A2(n_431), .B1(n_590), .B2(n_1242), .C1(n_1243), .C2(n_1244), .Y(n_1241) );
AOI22xp33_ASAP7_75t_SL g1430 ( .A1(n_426), .A2(n_431), .B1(n_1386), .B2(n_1387), .Y(n_1430) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g846 ( .A(n_428), .Y(n_846) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g1825 ( .A(n_429), .Y(n_1825) );
AOI222xp33_ASAP7_75t_SL g441 ( .A1(n_430), .A2(n_433), .B1(n_442), .B2(n_443), .C1(n_451), .C2(n_455), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_431), .A2(n_655), .B1(n_656), .B2(n_659), .C1(n_660), .C2(n_661), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g743 ( .A1(n_431), .A2(n_729), .B1(n_731), .B2(n_744), .C1(n_745), .C2(n_747), .Y(n_743) );
INVx3_ASAP7_75t_L g847 ( .A(n_431), .Y(n_847) );
AOI222xp33_ASAP7_75t_L g958 ( .A1(n_431), .A2(n_845), .B1(n_944), .B2(n_959), .C1(n_961), .C2(n_962), .Y(n_958) );
AOI222xp33_ASAP7_75t_L g1007 ( .A1(n_431), .A2(n_845), .B1(n_1002), .B2(n_1008), .C1(n_1009), .C2(n_1010), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_431), .A2(n_747), .B1(n_1026), .B2(n_1028), .Y(n_1035) );
AOI222xp33_ASAP7_75t_L g1092 ( .A1(n_431), .A2(n_745), .B1(n_747), .B2(n_1083), .C1(n_1084), .C2(n_1093), .Y(n_1092) );
AOI222xp33_ASAP7_75t_L g1133 ( .A1(n_431), .A2(n_747), .B1(n_1134), .B2(n_1135), .C1(n_1137), .C2(n_1138), .Y(n_1133) );
AOI222xp33_ASAP7_75t_L g1302 ( .A1(n_431), .A2(n_660), .B1(n_1295), .B2(n_1297), .C1(n_1303), .C2(n_1305), .Y(n_1302) );
AOI222xp33_ASAP7_75t_L g1342 ( .A1(n_431), .A2(n_660), .B1(n_1343), .B2(n_1344), .C1(n_1345), .C2(n_1346), .Y(n_1342) );
AOI222xp33_ASAP7_75t_L g1395 ( .A1(n_431), .A2(n_747), .B1(n_1386), .B2(n_1387), .C1(n_1396), .C2(n_1397), .Y(n_1395) );
AOI222xp33_ASAP7_75t_L g1446 ( .A1(n_431), .A2(n_660), .B1(n_790), .B2(n_1447), .C1(n_1448), .C2(n_1449), .Y(n_1446) );
AOI222xp33_ASAP7_75t_L g1498 ( .A1(n_431), .A2(n_660), .B1(n_689), .B2(n_1487), .C1(n_1488), .C2(n_1499), .Y(n_1498) );
AOI222xp33_ASAP7_75t_L g1877 ( .A1(n_431), .A2(n_747), .B1(n_1878), .B2(n_1879), .C1(n_1880), .C2(n_1881), .Y(n_1877) );
BUFx3_ASAP7_75t_L g1828 ( .A(n_432), .Y(n_1828) );
AOI211x1_ASAP7_75t_L g646 ( .A1(n_434), .A2(n_647), .B(n_665), .C(n_699), .Y(n_646) );
OAI31xp33_ASAP7_75t_L g794 ( .A1(n_434), .A2(n_795), .A3(n_796), .B(n_802), .Y(n_794) );
AOI211xp5_ASAP7_75t_L g836 ( .A1(n_434), .A2(n_837), .B(n_851), .C(n_861), .Y(n_836) );
AOI211xp5_ASAP7_75t_L g886 ( .A1(n_434), .A2(n_887), .B(n_899), .C(n_912), .Y(n_886) );
OAI31xp33_ASAP7_75t_SL g955 ( .A1(n_434), .A2(n_956), .A3(n_957), .B(n_963), .Y(n_955) );
OAI31xp33_ASAP7_75t_L g1003 ( .A1(n_434), .A2(n_1004), .A3(n_1005), .B(n_1006), .Y(n_1003) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
AND2x4_ASAP7_75t_L g643 ( .A(n_435), .B(n_437), .Y(n_643) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g552 ( .A(n_436), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g1855 ( .A(n_437), .Y(n_1855) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g536 ( .A(n_438), .Y(n_536) );
OR2x6_ASAP7_75t_L g595 ( .A(n_438), .B(n_596), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_477), .B(n_488), .Y(n_439) );
NAND3xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_463), .C(n_474), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_442), .A2(n_464), .B1(n_543), .B2(n_555), .C(n_557), .Y(n_554) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g1082 ( .A(n_444), .Y(n_1082) );
INVx1_ASAP7_75t_L g1145 ( .A(n_444), .Y(n_1145) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g1293 ( .A1(n_445), .A2(n_455), .B1(n_1294), .B2(n_1295), .C1(n_1296), .C2(n_1297), .Y(n_1293) );
AND2x4_ASAP7_75t_L g1779 ( .A(n_445), .B(n_1773), .Y(n_1779) );
HB1xp67_ASAP7_75t_L g1801 ( .A(n_445), .Y(n_1801) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g475 ( .A(n_446), .B(n_476), .Y(n_475) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_446), .Y(n_682) );
BUFx3_ASAP7_75t_L g761 ( .A(n_446), .Y(n_761) );
BUFx3_ASAP7_75t_L g827 ( .A(n_446), .Y(n_827) );
INVx1_ASAP7_75t_L g867 ( .A(n_446), .Y(n_867) );
BUFx6f_ASAP7_75t_L g904 ( .A(n_446), .Y(n_904) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g458 ( .A(n_448), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_448), .B(n_450), .Y(n_468) );
INVx2_ASAP7_75t_L g482 ( .A(n_448), .Y(n_482) );
AND2x4_ASAP7_75t_L g487 ( .A(n_448), .B(n_449), .Y(n_487) );
AND2x2_ASAP7_75t_L g681 ( .A(n_448), .B(n_450), .Y(n_681) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g454 ( .A(n_450), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_450), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g501 ( .A(n_450), .Y(n_501) );
INVx1_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_451), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_630) );
INVx2_ASAP7_75t_L g704 ( .A(n_451), .Y(n_704) );
INVx2_ASAP7_75t_L g733 ( .A(n_451), .Y(n_733) );
AOI222xp33_ASAP7_75t_L g825 ( .A1(n_451), .A2(n_633), .B1(n_800), .B2(n_801), .C1(n_821), .C2(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g906 ( .A(n_451), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_451), .A2(n_633), .B1(n_961), .B2(n_962), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_451), .A2(n_633), .B1(n_1009), .B2(n_1010), .Y(n_1014) );
AOI222xp33_ASAP7_75t_L g1025 ( .A1(n_451), .A2(n_633), .B1(n_682), .B2(n_1026), .C1(n_1027), .C2(n_1028), .Y(n_1025) );
AOI222xp33_ASAP7_75t_L g1080 ( .A1(n_451), .A2(n_633), .B1(n_1081), .B2(n_1082), .C1(n_1083), .C2(n_1084), .Y(n_1080) );
AOI222xp33_ASAP7_75t_L g1485 ( .A1(n_451), .A2(n_455), .B1(n_904), .B2(n_1486), .C1(n_1487), .C2(n_1488), .Y(n_1485) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
OR2x6_ASAP7_75t_L g466 ( .A(n_452), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g537 ( .A(n_453), .B(n_492), .Y(n_537) );
OR2x2_ASAP7_75t_L g705 ( .A(n_453), .B(n_457), .Y(n_705) );
OR2x2_ASAP7_75t_L g855 ( .A(n_453), .B(n_457), .Y(n_855) );
HB1xp67_ASAP7_75t_L g1772 ( .A(n_454), .Y(n_1772) );
AOI222xp33_ASAP7_75t_L g1199 ( .A1(n_455), .A2(n_732), .B1(n_1082), .B2(n_1200), .C1(n_1201), .C2(n_1202), .Y(n_1199) );
AOI222xp33_ASAP7_75t_L g1384 ( .A1(n_455), .A2(n_732), .B1(n_760), .B2(n_1385), .C1(n_1386), .C2(n_1387), .Y(n_1384) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_459), .Y(n_455) );
AND2x4_ASAP7_75t_L g633 ( .A(n_456), .B(n_459), .Y(n_633) );
AND2x4_ASAP7_75t_L g1777 ( .A(n_456), .B(n_1773), .Y(n_1777) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_458), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g533 ( .A(n_458), .B(n_514), .Y(n_533) );
INVxp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g476 ( .A(n_460), .Y(n_476) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_461), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g473 ( .A(n_462), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_469), .B2(n_470), .Y(n_463) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_465), .A2(n_663), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_465), .A2(n_709), .B1(n_735), .B2(n_736), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_465), .A2(n_470), .B1(n_820), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_465), .A2(n_707), .B1(n_857), .B2(n_858), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_465), .A2(n_707), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_465), .A2(n_713), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_465), .A2(n_470), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_465), .A2(n_713), .B1(n_1131), .B2(n_1147), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_465), .A2(n_470), .B1(n_1193), .B2(n_1204), .Y(n_1203) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_465), .A2(n_713), .B1(n_1246), .B2(n_1253), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_465), .A2(n_713), .B1(n_1299), .B2(n_1300), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1373 ( .A1(n_465), .A2(n_470), .B1(n_1348), .B2(n_1374), .Y(n_1373) );
AOI22xp5_ASAP7_75t_L g1388 ( .A1(n_465), .A2(n_470), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
AOI22xp33_ASAP7_75t_SL g1457 ( .A1(n_465), .A2(n_713), .B1(n_1444), .B2(n_1458), .Y(n_1457) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_465), .A2(n_470), .B1(n_1490), .B2(n_1491), .Y(n_1489) );
AOI22xp33_ASAP7_75t_L g1902 ( .A1(n_465), .A2(n_713), .B1(n_1875), .B2(n_1903), .Y(n_1902) );
INVx8_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g1526 ( .A(n_466), .B(n_1527), .Y(n_1526) );
OR2x6_ASAP7_75t_L g471 ( .A(n_467), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g508 ( .A(n_467), .Y(n_508) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_467), .Y(n_530) );
INVx2_ASAP7_75t_SL g607 ( .A(n_467), .Y(n_607) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_467), .Y(n_809) );
OR2x2_ASAP7_75t_L g1807 ( .A(n_467), .B(n_1774), .Y(n_1807) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_470), .A2(n_707), .B1(n_726), .B2(n_727), .Y(n_725) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx5_ASAP7_75t_L g713 ( .A(n_471), .Y(n_713) );
INVx1_ASAP7_75t_L g479 ( .A(n_472), .Y(n_479) );
AND2x4_ASAP7_75t_L g484 ( .A(n_472), .B(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g707 ( .A(n_472), .B(n_499), .Y(n_707) );
AND2x4_ASAP7_75t_L g709 ( .A(n_472), .B(n_485), .Y(n_709) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g596 ( .A(n_473), .B(n_493), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_474), .B(n_725), .C(n_728), .D(n_734), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_474), .B(n_825), .C(n_828), .Y(n_824) );
NAND3xp33_ASAP7_75t_L g1024 ( .A(n_474), .B(n_1025), .C(n_1029), .Y(n_1024) );
NAND4xp25_ASAP7_75t_L g1076 ( .A(n_474), .B(n_1077), .C(n_1080), .D(n_1085), .Y(n_1076) );
NAND4xp25_ASAP7_75t_SL g1139 ( .A(n_474), .B(n_1140), .C(n_1143), .D(n_1146), .Y(n_1139) );
NAND4xp25_ASAP7_75t_SL g1195 ( .A(n_474), .B(n_1196), .C(n_1199), .D(n_1203), .Y(n_1195) );
NAND4xp25_ASAP7_75t_L g1289 ( .A(n_474), .B(n_1290), .C(n_1293), .D(n_1298), .Y(n_1289) );
NAND4xp25_ASAP7_75t_L g1380 ( .A(n_474), .B(n_1381), .C(n_1384), .D(n_1388), .Y(n_1380) );
NAND4xp25_ASAP7_75t_L g1481 ( .A(n_474), .B(n_1482), .C(n_1485), .D(n_1489), .Y(n_1481) );
CKINVDCx11_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
AOI211xp5_ASAP7_75t_L g700 ( .A1(n_475), .A2(n_701), .B(n_702), .C(n_703), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g852 ( .A1(n_475), .A2(n_826), .B(n_853), .C(n_854), .Y(n_852) );
AOI211xp5_ASAP7_75t_L g900 ( .A1(n_475), .A2(n_901), .B(n_902), .C(n_905), .Y(n_900) );
AOI211xp5_ASAP7_75t_L g1254 ( .A1(n_475), .A2(n_866), .B(n_1255), .C(n_1256), .Y(n_1254) );
AOI211xp5_ASAP7_75t_L g1370 ( .A1(n_475), .A2(n_760), .B(n_1371), .C(n_1372), .Y(n_1370) );
AOI211xp5_ASAP7_75t_L g1451 ( .A1(n_475), .A2(n_702), .B(n_1452), .C(n_1453), .Y(n_1451) );
AOI211xp5_ASAP7_75t_L g1896 ( .A1(n_475), .A2(n_760), .B(n_1897), .C(n_1898), .Y(n_1896) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g601 ( .A(n_481), .Y(n_601) );
INVx1_ASAP7_75t_L g614 ( .A(n_481), .Y(n_614) );
AND2x4_ASAP7_75t_L g499 ( .A(n_482), .B(n_500), .Y(n_499) );
INVx5_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_484), .A2(n_713), .B1(n_840), .B2(n_860), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_484), .A2(n_713), .B1(n_891), .B2(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_484), .A2(n_707), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_484), .A2(n_707), .B1(n_1197), .B2(n_1198), .Y(n_1196) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_484), .A2(n_707), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
AOI22xp5_ASAP7_75t_L g1381 ( .A1(n_484), .A2(n_707), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_484), .A2(n_707), .B1(n_1483), .B2(n_1484), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1899 ( .A1(n_484), .A2(n_707), .B1(n_1900), .B2(n_1901), .Y(n_1899) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_486), .Y(n_872) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_487), .Y(n_504) );
INVx3_ASAP7_75t_L g527 ( .A(n_487), .Y(n_527) );
INVx1_ASAP7_75t_L g1220 ( .A(n_487), .Y(n_1220) );
OAI31xp33_ASAP7_75t_SL g626 ( .A1(n_488), .A2(n_627), .A3(n_628), .B(n_634), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_488), .A2(n_724), .B1(n_737), .B2(n_748), .C(n_750), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_488), .A2(n_824), .B(n_830), .Y(n_823) );
OAI31xp33_ASAP7_75t_SL g964 ( .A1(n_488), .A2(n_965), .A3(n_966), .B(n_969), .Y(n_964) );
OAI31xp33_ASAP7_75t_SL g1011 ( .A1(n_488), .A2(n_1012), .A3(n_1013), .B(n_1015), .Y(n_1011) );
O2A1O1Ixp33_ASAP7_75t_L g1022 ( .A1(n_488), .A2(n_1023), .B(n_1024), .C(n_1032), .Y(n_1022) );
AOI221x1_ASAP7_75t_L g1075 ( .A1(n_488), .A2(n_643), .B1(n_1076), .B2(n_1088), .C(n_1098), .Y(n_1075) );
AOI221x1_ASAP7_75t_L g1125 ( .A1(n_488), .A2(n_1040), .B1(n_1126), .B2(n_1139), .C(n_1148), .Y(n_1125) );
AOI221x1_ASAP7_75t_L g1182 ( .A1(n_488), .A2(n_1040), .B1(n_1183), .B2(n_1195), .C(n_1205), .Y(n_1182) );
AOI221x1_ASAP7_75t_L g1288 ( .A1(n_488), .A2(n_643), .B1(n_1289), .B2(n_1301), .C(n_1311), .Y(n_1288) );
AOI221x1_ASAP7_75t_L g1379 ( .A1(n_488), .A2(n_1040), .B1(n_1380), .B2(n_1391), .C(n_1400), .Y(n_1379) );
OAI31xp33_ASAP7_75t_L g1420 ( .A1(n_488), .A2(n_1421), .A3(n_1422), .B(n_1425), .Y(n_1420) );
AOI221xp5_ASAP7_75t_L g1480 ( .A1(n_488), .A2(n_643), .B1(n_1481), .B2(n_1492), .C(n_1500), .Y(n_1480) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
AOI31xp33_ASAP7_75t_SL g1369 ( .A1(n_489), .A2(n_1370), .A3(n_1373), .B(n_1375), .Y(n_1369) );
AOI31xp33_ASAP7_75t_L g1450 ( .A1(n_489), .A2(n_1451), .A3(n_1454), .B(n_1457), .Y(n_1450) );
AOI31xp33_ASAP7_75t_L g1895 ( .A1(n_489), .A2(n_1896), .A3(n_1899), .B(n_1902), .Y(n_1895) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x4_ASAP7_75t_L g551 ( .A(n_490), .B(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g686 ( .A(n_490), .B(n_552), .Y(n_686) );
OR2x2_ASAP7_75t_L g714 ( .A(n_490), .B(n_491), .Y(n_714) );
AND2x4_ASAP7_75t_L g1809 ( .A(n_490), .B(n_1810), .Y(n_1809) );
INVxp67_ASAP7_75t_L g1527 ( .A(n_491), .Y(n_1527) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_515), .B1(n_521), .B2(n_534), .C(n_538), .Y(n_494) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g1782 ( .A(n_498), .B(n_1783), .Y(n_1782) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g523 ( .A(n_499), .Y(n_523) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_499), .Y(n_676) );
BUFx2_ASAP7_75t_L g766 ( .A(n_499), .Y(n_766) );
BUFx2_ASAP7_75t_L g805 ( .A(n_499), .Y(n_805) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_499), .Y(n_870) );
INVx1_ASAP7_75t_L g1227 ( .A(n_499), .Y(n_1227) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g768 ( .A(n_504), .Y(n_768) );
BUFx3_ASAP7_75t_L g806 ( .A(n_504), .Y(n_806) );
INVx2_ASAP7_75t_SL g1152 ( .A(n_504), .Y(n_1152) );
INVx4_ASAP7_75t_L g1157 ( .A(n_504), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_509), .B2(n_510), .Y(n_505) );
OAI22xp33_ASAP7_75t_SL g812 ( .A1(n_507), .A2(n_532), .B1(n_813), .B2(n_814), .Y(n_812) );
OAI22xp5_ASAP7_75t_SL g1045 ( .A1(n_507), .A2(n_510), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx3_ASAP7_75t_L g629 ( .A(n_512), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_512), .A2(n_530), .B1(n_931), .B2(n_932), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g994 ( .A1(n_512), .A2(n_606), .B1(n_981), .B2(n_984), .Y(n_994) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_515), .A2(n_534), .B1(n_804), .B2(n_811), .C(n_815), .Y(n_803) );
AOI33xp33_ASAP7_75t_L g1883 ( .A1(n_515), .A2(n_762), .A3(n_1884), .B1(n_1886), .B2(n_1887), .B3(n_1888), .Y(n_1883) );
INVx6_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx5_ASAP7_75t_L g625 ( .A(n_516), .Y(n_625) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_519), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g1783 ( .A(n_518), .B(n_1784), .Y(n_1783) );
INVx2_ASAP7_75t_L g684 ( .A(n_519), .Y(n_684) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g1319 ( .A(n_523), .Y(n_1319) );
INVx1_ASAP7_75t_L g1362 ( .A(n_523), .Y(n_1362) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g603 ( .A(n_525), .Y(n_603) );
OAI22xp33_ASAP7_75t_SL g933 ( .A1(n_525), .A2(n_934), .B1(n_935), .B2(n_936), .Y(n_933) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g619 ( .A(n_526), .Y(n_619) );
INVx2_ASAP7_75t_L g1267 ( .A(n_526), .Y(n_1267) );
INVx2_ASAP7_75t_L g1466 ( .A(n_526), .Y(n_1466) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g755 ( .A(n_527), .Y(n_755) );
BUFx6f_ASAP7_75t_L g1315 ( .A(n_527), .Y(n_1315) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g542 ( .A1(n_529), .A2(n_531), .B1(n_543), .B2(n_545), .C(n_547), .Y(n_542) );
INVx1_ASAP7_75t_L g609 ( .A(n_532), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g807 ( .A1(n_532), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_532), .A2(n_606), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g622 ( .A(n_533), .Y(n_622) );
INVx2_ASAP7_75t_L g943 ( .A(n_533), .Y(n_943) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI33xp33_ASAP7_75t_L g685 ( .A1(n_535), .A2(n_686), .A3(n_687), .B1(n_691), .B2(n_696), .B3(n_697), .Y(n_685) );
INVx2_ASAP7_75t_L g763 ( .A(n_535), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g862 ( .A(n_535), .B(n_863), .C(n_864), .Y(n_862) );
NAND3xp33_ASAP7_75t_L g913 ( .A(n_535), .B(n_914), .C(n_915), .Y(n_913) );
AOI33xp33_ASAP7_75t_L g1215 ( .A1(n_535), .A2(n_625), .A3(n_1216), .B1(n_1221), .B2(n_1225), .B3(n_1231), .Y(n_1215) );
NAND3xp33_ASAP7_75t_L g1312 ( .A(n_535), .B(n_1313), .C(n_1316), .Y(n_1312) );
NAND3xp33_ASAP7_75t_L g1402 ( .A(n_535), .B(n_1403), .C(n_1404), .Y(n_1402) );
NAND3xp33_ASAP7_75t_L g1460 ( .A(n_535), .B(n_1461), .C(n_1462), .Y(n_1460) );
NAND3xp33_ASAP7_75t_L g1501 ( .A(n_535), .B(n_1502), .C(n_1503), .Y(n_1501) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OR2x2_ASAP7_75t_L g539 ( .A(n_536), .B(n_540), .Y(n_539) );
OR2x6_ASAP7_75t_L g565 ( .A(n_536), .B(n_540), .Y(n_565) );
OR2x2_ASAP7_75t_L g668 ( .A(n_536), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g683 ( .A(n_536), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g1263 ( .A(n_536), .B(n_537), .Y(n_1263) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_539), .A2(n_542), .B1(n_550), .B2(n_554), .Y(n_538) );
OAI22xp5_ASAP7_75t_SL g815 ( .A1(n_539), .A2(n_550), .B1(n_816), .B2(n_819), .Y(n_815) );
OAI33xp33_ASAP7_75t_L g973 ( .A1(n_539), .A2(n_974), .A3(n_980), .B1(n_986), .B2(n_989), .B3(n_992), .Y(n_973) );
INVx1_ASAP7_75t_L g1842 ( .A(n_540), .Y(n_1842) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g669 ( .A(n_541), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_543), .A2(n_545), .B1(n_1046), .B2(n_1047), .C(n_1060), .Y(n_1059) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g817 ( .A(n_544), .Y(n_817) );
INVx2_ASAP7_75t_L g948 ( .A(n_544), .Y(n_948) );
OAI221xp5_ASAP7_75t_L g816 ( .A1(n_545), .A2(n_808), .B1(n_810), .B2(n_817), .C(n_818), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_545), .A2(n_817), .B1(n_820), .B2(n_821), .C(n_822), .Y(n_819) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_545), .A2(n_1027), .B1(n_1064), .B2(n_1066), .C(n_1067), .Y(n_1063) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g640 ( .A(n_546), .Y(n_640) );
INVx2_ASAP7_75t_SL g575 ( .A(n_548), .Y(n_575) );
INVx1_ASAP7_75t_L g778 ( .A(n_548), .Y(n_778) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_548), .Y(n_1061) );
AND2x4_ASAP7_75t_L g1818 ( .A(n_548), .B(n_1819), .Y(n_1818) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_550), .A2(n_565), .B1(n_566), .B2(n_578), .Y(n_564) );
INVx1_ASAP7_75t_L g783 ( .A(n_550), .Y(n_783) );
OAI22xp5_ASAP7_75t_SL g946 ( .A1(n_550), .A2(n_668), .B1(n_947), .B2(n_950), .Y(n_946) );
OAI22xp5_ASAP7_75t_SL g1058 ( .A1(n_550), .A2(n_565), .B1(n_1059), .B2(n_1063), .Y(n_1058) );
INVx4_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx4f_ASAP7_75t_L g1177 ( .A(n_551), .Y(n_1177) );
BUFx4f_ASAP7_75t_L g1207 ( .A(n_551), .Y(n_1207) );
INVx1_ASAP7_75t_L g1832 ( .A(n_552), .Y(n_1832) );
AND2x4_ASAP7_75t_L g1811 ( .A(n_553), .B(n_1812), .Y(n_1811) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g985 ( .A(n_556), .Y(n_985) );
INVx1_ASAP7_75t_L g979 ( .A(n_558), .Y(n_979) );
BUFx6f_ASAP7_75t_L g1062 ( .A(n_558), .Y(n_1062) );
INVx1_ASAP7_75t_L g1070 ( .A(n_558), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1515 ( .A(n_558), .Y(n_1515) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_644), .B1(n_645), .B2(n_717), .Y(n_560) );
INVx1_ASAP7_75t_L g717 ( .A(n_561), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_626), .C(n_635), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_592), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_565), .Y(n_781) );
INVx2_ASAP7_75t_L g1100 ( .A(n_565), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g1359 ( .A(n_565), .Y(n_1359) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_569), .B2(n_572), .C(n_573), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_567), .A2(n_572), .B1(n_606), .B2(n_608), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g1830 ( .A1(n_568), .A2(n_1186), .B1(n_1785), .B2(n_1789), .C(n_1831), .Y(n_1830) );
OAI221xp5_ASAP7_75t_L g947 ( .A1(n_569), .A2(n_931), .B1(n_932), .B2(n_948), .C(n_949), .Y(n_947) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_577), .A2(n_778), .B1(n_990), .B2(n_991), .Y(n_989) );
INVx1_ASAP7_75t_L g1169 ( .A(n_577), .Y(n_1169) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B1(n_583), .B2(n_585), .C(n_586), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx3_ASAP7_75t_L g1065 ( .A(n_589), .Y(n_1065) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_589), .Y(n_1102) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI33xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_597), .A3(n_605), .B1(n_610), .B2(n_616), .B3(n_624), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI33xp33_ASAP7_75t_L g929 ( .A1(n_595), .A2(n_930), .A3(n_933), .B1(n_937), .B2(n_941), .B3(n_945), .Y(n_929) );
OAI33xp33_ASAP7_75t_L g993 ( .A1(n_595), .A2(n_945), .A3(n_994), .B1(n_995), .B2(n_996), .B3(n_1000), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_602), .B2(n_604), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_606), .A2(n_611), .B1(n_612), .B2(n_615), .Y(n_610) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g1423 ( .A(n_609), .Y(n_1423) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g935 ( .A(n_614), .Y(n_935) );
INVx1_ASAP7_75t_L g997 ( .A(n_614), .Y(n_997) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B1(n_621), .B2(n_623), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g967 ( .A(n_622), .Y(n_967) );
INVx1_ASAP7_75t_L g1057 ( .A(n_624), .Y(n_1057) );
CKINVDCx8_ASAP7_75t_R g624 ( .A(n_625), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g764 ( .A(n_625), .B(n_765), .C(n_769), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g1154 ( .A(n_625), .B(n_1155), .C(n_1158), .Y(n_1154) );
AOI33xp33_ASAP7_75t_L g1261 ( .A1(n_625), .A2(n_1262), .A3(n_1264), .B1(n_1265), .B2(n_1268), .B3(n_1269), .Y(n_1261) );
NAND3xp33_ASAP7_75t_L g1360 ( .A(n_625), .B(n_1361), .C(n_1363), .Y(n_1360) );
NAND3xp33_ASAP7_75t_L g1463 ( .A(n_625), .B(n_1464), .C(n_1467), .Y(n_1463) );
NAND3xp33_ASAP7_75t_L g1504 ( .A(n_625), .B(n_1505), .C(n_1506), .Y(n_1504) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_629), .Y(n_1056) );
AOI222xp33_ASAP7_75t_L g728 ( .A1(n_633), .A2(n_702), .B1(n_729), .B2(n_730), .C1(n_731), .C2(n_732), .Y(n_728) );
AOI222xp33_ASAP7_75t_L g1143 ( .A1(n_633), .A2(n_732), .B1(n_1137), .B2(n_1138), .C1(n_1144), .C2(n_1145), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1424 ( .A1(n_633), .A2(n_1296), .B1(n_1386), .B2(n_1387), .Y(n_1424) );
OAI31xp33_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_637), .A3(n_638), .B(n_643), .Y(n_635) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g737 ( .A(n_641), .B(n_738), .C(n_741), .D(n_743), .Y(n_737) );
NAND4xp25_ASAP7_75t_L g837 ( .A(n_641), .B(n_838), .C(n_841), .D(n_848), .Y(n_837) );
NAND4xp25_ASAP7_75t_L g887 ( .A(n_641), .B(n_888), .C(n_892), .D(n_895), .Y(n_887) );
BUFx2_ASAP7_75t_L g1089 ( .A(n_641), .Y(n_1089) );
NAND4xp25_ASAP7_75t_L g1391 ( .A(n_641), .B(n_1392), .C(n_1395), .D(n_1398), .Y(n_1391) );
NAND4xp25_ASAP7_75t_SL g1439 ( .A(n_641), .B(n_1440), .C(n_1443), .D(n_1446), .Y(n_1439) );
NAND4xp25_ASAP7_75t_SL g1870 ( .A(n_641), .B(n_1871), .C(n_1874), .D(n_1877), .Y(n_1870) );
INVx1_ASAP7_75t_L g749 ( .A(n_643), .Y(n_749) );
BUFx6f_ASAP7_75t_L g1040 ( .A(n_643), .Y(n_1040) );
AOI211x1_ASAP7_75t_SL g1239 ( .A1(n_643), .A2(n_1240), .B(n_1251), .C(n_1260), .Y(n_1239) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g716 ( .A(n_646), .Y(n_716) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_650), .Y(n_1096) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g775 ( .A(n_652), .Y(n_775) );
INVx1_ASAP7_75t_L g876 ( .A(n_652), .Y(n_876) );
INVx2_ASAP7_75t_L g1108 ( .A(n_652), .Y(n_1108) );
BUFx6f_ASAP7_75t_L g1165 ( .A(n_652), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_652), .Y(n_1173) );
INVx2_ASAP7_75t_SL g1279 ( .A(n_652), .Y(n_1279) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx4f_ASAP7_75t_L g746 ( .A(n_658), .Y(n_746) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_658), .Y(n_790) );
INVx2_ASAP7_75t_SL g960 ( .A(n_658), .Y(n_960) );
BUFx3_ASAP7_75t_L g1174 ( .A(n_658), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1835 ( .A(n_658), .B(n_1819), .Y(n_1835) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_685), .Y(n_665) );
AOI33xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .A3(n_671), .B1(n_675), .B2(n_677), .B3(n_683), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g874 ( .A(n_667), .B(n_875), .C(n_877), .Y(n_874) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_667), .B(n_920), .C(n_921), .Y(n_919) );
AOI33xp33_ASAP7_75t_L g1206 ( .A1(n_667), .A2(n_1207), .A3(n_1208), .B1(n_1210), .B2(n_1213), .B3(n_1214), .Y(n_1206) );
NAND3xp33_ASAP7_75t_L g1321 ( .A(n_667), .B(n_1322), .C(n_1324), .Y(n_1321) );
NAND3xp33_ASAP7_75t_L g1410 ( .A(n_667), .B(n_1411), .C(n_1412), .Y(n_1410) );
NAND3xp33_ASAP7_75t_L g1468 ( .A(n_667), .B(n_1469), .C(n_1470), .Y(n_1468) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g688 ( .A(n_673), .Y(n_688) );
HB1xp67_ASAP7_75t_L g1396 ( .A(n_674), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g1879 ( .A(n_674), .Y(n_1879) );
BUFx3_ASAP7_75t_L g1800 ( .A(n_676), .Y(n_1800) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g698 ( .A(n_679), .Y(n_698) );
INVx2_ASAP7_75t_L g865 ( .A(n_679), .Y(n_865) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_680), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1409 ( .A(n_680), .Y(n_1409) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx3_ASAP7_75t_L g759 ( .A(n_681), .Y(n_759) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_682), .Y(n_702) );
INVx2_ASAP7_75t_SL g771 ( .A(n_682), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g868 ( .A(n_683), .B(n_869), .C(n_873), .Y(n_868) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_683), .B(n_917), .C(n_918), .Y(n_916) );
INVx1_ASAP7_75t_L g945 ( .A(n_683), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g1317 ( .A(n_683), .B(n_1318), .C(n_1320), .Y(n_1317) );
NAND3xp33_ASAP7_75t_L g1405 ( .A(n_683), .B(n_1406), .C(n_1408), .Y(n_1405) );
NAND3xp33_ASAP7_75t_L g880 ( .A(n_686), .B(n_881), .C(n_883), .Y(n_880) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_686), .B(n_923), .C(n_924), .Y(n_922) );
INVx1_ASAP7_75t_L g992 ( .A(n_686), .Y(n_992) );
AOI33xp33_ASAP7_75t_L g1271 ( .A1(n_686), .A2(n_1100), .A3(n_1272), .B1(n_1275), .B2(n_1276), .B3(n_1280), .Y(n_1271) );
NAND3xp33_ASAP7_75t_L g1325 ( .A(n_686), .B(n_1326), .C(n_1327), .Y(n_1325) );
NAND3xp33_ASAP7_75t_L g1415 ( .A(n_686), .B(n_1416), .C(n_1417), .Y(n_1415) );
NAND3xp33_ASAP7_75t_L g1471 ( .A(n_686), .B(n_1472), .C(n_1473), .Y(n_1471) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_688), .Y(n_1112) );
INVx1_ASAP7_75t_L g1136 ( .A(n_689), .Y(n_1136) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx3_ASAP7_75t_L g1008 ( .A(n_690), .Y(n_1008) );
INVx2_ASAP7_75t_SL g786 ( .A(n_692), .Y(n_786) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g1104 ( .A(n_694), .Y(n_1104) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g1854 ( .A(n_695), .B(n_1820), .Y(n_1854) );
INVx1_ASAP7_75t_L g1894 ( .A(n_695), .Y(n_1894) );
AOI31xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_706), .A3(n_711), .B(n_714), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_707), .A2(n_709), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_707), .A2(n_709), .B1(n_1291), .B2(n_1292), .Y(n_1290) );
AOI22xp5_ASAP7_75t_SL g1375 ( .A1(n_707), .A2(n_709), .B1(n_1376), .B2(n_1377), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_707), .A2(n_709), .B1(n_1455), .B2(n_1456), .Y(n_1454) );
AOI31xp33_ASAP7_75t_L g851 ( .A1(n_714), .A2(n_852), .A3(n_856), .B(n_859), .Y(n_851) );
AOI31xp33_ASAP7_75t_L g899 ( .A1(n_714), .A2(n_900), .A3(n_907), .B(n_910), .Y(n_899) );
AOI31xp33_ASAP7_75t_L g1251 ( .A1(n_714), .A2(n_1252), .A3(n_1254), .B(n_1257), .Y(n_1251) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_1018), .Y(n_718) );
XNOR2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_831), .Y(n_719) );
XNOR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_791), .Y(n_720) );
XNOR2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AOI31xp33_ASAP7_75t_L g1338 ( .A1(n_749), .A2(n_1339), .A3(n_1342), .B(n_1347), .Y(n_1338) );
NAND4xp25_ASAP7_75t_L g750 ( .A(n_751), .B(n_764), .C(n_772), .D(n_782), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_756), .C(n_762), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g939 ( .A(n_755), .Y(n_939) );
BUFx3_ASAP7_75t_L g1043 ( .A(n_755), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1794 ( .A(n_755), .B(n_1783), .Y(n_1794) );
BUFx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_759), .Y(n_1161) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_759), .Y(n_1223) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g1234 ( .A(n_761), .Y(n_1234) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_762), .A2(n_1042), .B1(n_1048), .B2(n_1057), .C(n_1058), .Y(n_1041) );
AOI33xp33_ASAP7_75t_L g1113 ( .A1(n_762), .A2(n_1057), .A3(n_1114), .B1(n_1115), .B2(n_1116), .B3(n_1117), .Y(n_1113) );
NAND3xp33_ASAP7_75t_L g1149 ( .A(n_762), .B(n_1150), .C(n_1153), .Y(n_1149) );
AOI33xp33_ASAP7_75t_L g1795 ( .A1(n_762), .A2(n_1057), .A3(n_1796), .B1(n_1799), .B2(n_1802), .B3(n_1803), .Y(n_1795) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_766), .Y(n_1044) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_SL g1885 ( .A(n_771), .Y(n_1885) );
NAND3xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .C(n_781), .Y(n_772) );
BUFx3_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_775), .Y(n_1068) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g1511 ( .A(n_780), .Y(n_1511) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_781), .B(n_1163), .C(n_1166), .Y(n_1162) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .C(n_787), .Y(n_782) );
AOI33xp33_ASAP7_75t_L g1099 ( .A1(n_783), .A2(n_1100), .A3(n_1101), .B1(n_1105), .B2(n_1110), .B3(n_1111), .Y(n_1099) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_790), .Y(n_1109) );
BUFx2_ASAP7_75t_SL g1344 ( .A(n_790), .Y(n_1344) );
XNOR2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g1582 ( .A1(n_792), .A2(n_1537), .B1(n_1546), .B2(n_1583), .Y(n_1582) );
NAND3x1_ASAP7_75t_SL g793 ( .A(n_794), .B(n_803), .C(n_823), .Y(n_793) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_798), .A2(n_842), .B(n_843), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_798), .A2(n_896), .B(n_897), .Y(n_895) );
INVx1_ASAP7_75t_L g1054 ( .A(n_806), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g941 ( .A1(n_809), .A2(n_942), .B1(n_943), .B2(n_944), .Y(n_941) );
BUFx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x6_ASAP7_75t_L g1787 ( .A(n_827), .B(n_1783), .Y(n_1787) );
XOR2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_925), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B1(n_884), .B2(n_885), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g898 ( .A(n_845), .Y(n_898) );
NAND4xp25_ASAP7_75t_L g861 ( .A(n_862), .B(n_868), .C(n_874), .D(n_880), .Y(n_861) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_SL g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_L g1281 ( .A(n_879), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g1844 ( .A(n_882), .Y(n_1844) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_SL g903 ( .A(n_904), .Y(n_903) );
HB1xp67_ASAP7_75t_L g1224 ( .A(n_904), .Y(n_1224) );
INVx1_ASAP7_75t_L g1296 ( .A(n_906), .Y(n_1296) );
NAND4xp25_ASAP7_75t_L g912 ( .A(n_913), .B(n_916), .C(n_919), .D(n_922), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_970), .B1(n_1016), .B2(n_1017), .Y(n_925) );
INVx1_ASAP7_75t_L g1016 ( .A(n_926), .Y(n_1016) );
NAND3xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_955), .C(n_964), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_946), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_935), .A2(n_938), .B1(n_939), .B2(n_940), .Y(n_937) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_935), .A2(n_939), .B1(n_975), .B2(n_978), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_939), .A2(n_997), .B1(n_998), .B2(n_999), .Y(n_996) );
INVx2_ASAP7_75t_L g1168 ( .A(n_954), .Y(n_1168) );
BUFx3_ASAP7_75t_L g1354 ( .A(n_954), .Y(n_1354) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g1209 ( .A(n_960), .Y(n_1209) );
INVx1_ASAP7_75t_L g1017 ( .A(n_970), .Y(n_1017) );
NAND3xp33_ASAP7_75t_L g971 ( .A(n_972), .B(n_1003), .C(n_1011), .Y(n_971) );
NOR2xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_993), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_976), .B1(n_978), .B2(n_979), .Y(n_974) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
BUFx4f_ASAP7_75t_L g1211 ( .A(n_977), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B1(n_984), .B2(n_985), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_982), .A2(n_985), .B1(n_987), .B2(n_988), .Y(n_986) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1008), .Y(n_1840) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1072), .B1(n_1073), .B2(n_1119), .Y(n_1018) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1019), .Y(n_1119) );
INVx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1041), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1036), .B(n_1039), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
OAI31xp33_ASAP7_75t_L g1426 ( .A1(n_1040), .A2(n_1427), .A3(n_1428), .B(n_1431), .Y(n_1426) );
AOI211xp5_ASAP7_75t_L g1438 ( .A1(n_1040), .A2(n_1439), .B(n_1450), .C(n_1459), .Y(n_1438) );
AOI211x1_ASAP7_75t_SL g1869 ( .A1(n_1040), .A2(n_1870), .B(n_1882), .C(n_1895), .Y(n_1869) );
CKINVDCx5p33_ASAP7_75t_R g1798 ( .A(n_1043), .Y(n_1798) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
OAI22xp33_ASAP7_75t_SL g1052 ( .A1(n_1053), .A2(n_1054), .B1(n_1055), .B2(n_1056), .Y(n_1052) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx2_ASAP7_75t_SL g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1075), .Y(n_1118) );
NAND4xp25_ASAP7_75t_SL g1088 ( .A(n_1089), .B(n_1090), .C(n_1092), .D(n_1094), .Y(n_1088) );
NAND4xp25_ASAP7_75t_L g1126 ( .A(n_1089), .B(n_1127), .C(n_1130), .D(n_1133), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1113), .Y(n_1098) );
INVx2_ASAP7_75t_SL g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1104), .Y(n_1212) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
XOR2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1332), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
AO22x2_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1236), .B1(n_1237), .B2(n_1331), .Y(n_1122) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1123), .Y(n_1331) );
XNOR2xp5_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1180), .Y(n_1123) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1125), .Y(n_1179) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
NAND4xp25_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1154), .C(n_1162), .D(n_1170), .Y(n_1148) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
BUFx2_ASAP7_75t_L g1232 ( .A(n_1161), .Y(n_1232) );
AND2x4_ASAP7_75t_L g1791 ( .A(n_1161), .B(n_1783), .Y(n_1791) );
INVx4_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1165), .Y(n_1323) );
INVx2_ASAP7_75t_SL g1167 ( .A(n_1168), .Y(n_1167) );
NAND3xp33_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1175), .C(n_1177), .Y(n_1170) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
NAND3xp33_ASAP7_75t_L g1512 ( .A(n_1177), .B(n_1513), .C(n_1514), .Y(n_1512) );
AOI33xp33_ASAP7_75t_L g1889 ( .A1(n_1177), .A2(n_1359), .A3(n_1890), .B1(n_1891), .B2(n_1892), .B3(n_1893), .Y(n_1889) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
NAND3xp33_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1189), .C(n_1192), .Y(n_1183) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1429 ( .A(n_1188), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1215), .Y(n_1205) );
NAND3xp33_ASAP7_75t_L g1351 ( .A(n_1207), .B(n_1352), .C(n_1353), .Y(n_1351) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1220), .Y(n_1230) );
BUFx2_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1230), .Y(n_1367) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
AOI22xp5_ASAP7_75t_L g1237 ( .A1(n_1238), .A2(n_1286), .B1(n_1287), .B2(n_1330), .Y(n_1237) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1238), .Y(n_1330) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1239), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1271), .Y(n_1260) );
BUFx2_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
NAND3xp33_ASAP7_75t_L g1364 ( .A(n_1263), .B(n_1365), .C(n_1368), .Y(n_1364) );
INVx2_ASAP7_75t_SL g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1267), .Y(n_1270) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1274), .Y(n_1358) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
OAI22xp33_ASAP7_75t_L g1619 ( .A1(n_1284), .A2(n_1620), .B1(n_1621), .B2(n_1622), .Y(n_1619) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1288), .Y(n_1329) );
NAND3xp33_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1306), .C(n_1308), .Y(n_1301) );
BUFx6f_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
AND2x4_ASAP7_75t_L g1845 ( .A(n_1304), .B(n_1846), .Y(n_1845) );
NAND4xp25_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1317), .C(n_1321), .D(n_1325), .Y(n_1311) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx3_ASAP7_75t_L g1407 ( .A(n_1315), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_1333), .A2(n_1334), .B1(n_1477), .B2(n_1478), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_1335), .A2(n_1434), .B1(n_1435), .B2(n_1476), .Y(n_1334) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1335), .Y(n_1476) );
OAI22x1_ASAP7_75t_L g1335 ( .A1(n_1336), .A2(n_1378), .B1(n_1432), .B2(n_1433), .Y(n_1335) );
INVx2_ASAP7_75t_L g1432 ( .A(n_1336), .Y(n_1432) );
NOR3xp33_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1350), .C(n_1369), .Y(n_1337) );
NAND4xp25_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1355), .C(n_1360), .D(n_1364), .Y(n_1350) );
NAND3xp33_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1357), .C(n_1359), .Y(n_1355) );
NAND3xp33_ASAP7_75t_L g1507 ( .A(n_1359), .B(n_1508), .C(n_1509), .Y(n_1507) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1378), .Y(n_1433) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1381), .Y(n_1425) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1388), .Y(n_1421) );
INVxp67_ASAP7_75t_L g1427 ( .A(n_1392), .Y(n_1427) );
INVxp67_ASAP7_75t_L g1431 ( .A(n_1398), .Y(n_1431) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
NAND3xp33_ASAP7_75t_L g1419 ( .A(n_1401), .B(n_1420), .C(n_1426), .Y(n_1419) );
AND4x1_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1405), .C(n_1410), .D(n_1415), .Y(n_1401) );
INVx2_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1438), .Y(n_1475) );
NAND4xp25_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1463), .C(n_1468), .D(n_1471), .Y(n_1459) );
INVx2_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
HB1xp67_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1480), .Y(n_1517) );
NAND4xp25_ASAP7_75t_SL g1500 ( .A(n_1501), .B(n_1504), .C(n_1507), .D(n_1512), .Y(n_1500) );
BUFx3_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
AND2x4_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1525), .Y(n_1519) );
AND2x4_ASAP7_75t_L g1861 ( .A(n_1520), .B(n_1526), .Y(n_1861) );
NOR2xp33_ASAP7_75t_SL g1520 ( .A(n_1521), .B(n_1523), .Y(n_1520) );
INVx1_ASAP7_75t_SL g1907 ( .A(n_1521), .Y(n_1907) );
NAND2xp5_ASAP7_75t_L g1910 ( .A(n_1521), .B(n_1523), .Y(n_1910) );
HB1xp67_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1906 ( .A(n_1523), .B(n_1907), .Y(n_1906) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
OAI221xp5_ASAP7_75t_L g1528 ( .A1(n_1529), .A2(n_1764), .B1(n_1766), .B2(n_1856), .C(n_1862), .Y(n_1528) );
AOI311xp33_ASAP7_75t_L g1529 ( .A1(n_1530), .A2(n_1623), .A3(n_1651), .B(n_1658), .C(n_1730), .Y(n_1529) );
OAI211xp5_ASAP7_75t_L g1530 ( .A1(n_1531), .A2(n_1559), .B(n_1584), .C(n_1610), .Y(n_1530) );
A2O1A1Ixp33_ASAP7_75t_L g1584 ( .A1(n_1531), .A2(n_1585), .B(n_1589), .C(n_1595), .Y(n_1584) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_1532), .B(n_1676), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1532), .B(n_1652), .Y(n_1757) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx2_ASAP7_75t_SL g1600 ( .A(n_1533), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1533), .B(n_1592), .Y(n_1634) );
AND2x4_ASAP7_75t_L g1648 ( .A(n_1533), .B(n_1591), .Y(n_1648) );
NAND2xp5_ASAP7_75t_L g1673 ( .A(n_1533), .B(n_1652), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1533), .B(n_1680), .Y(n_1679) );
NOR2xp33_ASAP7_75t_L g1721 ( .A(n_1533), .B(n_1680), .Y(n_1721) );
HB1xp67_ASAP7_75t_L g1748 ( .A(n_1533), .Y(n_1748) );
CKINVDCx5p33_ASAP7_75t_R g1533 ( .A(n_1534), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1534), .B(n_1592), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1534), .B(n_1591), .Y(n_1686) );
OR2x2_ASAP7_75t_L g1534 ( .A(n_1535), .B(n_1549), .Y(n_1534) );
OAI22xp5_ASAP7_75t_L g1535 ( .A1(n_1536), .A2(n_1543), .B1(n_1544), .B2(n_1548), .Y(n_1535) );
BUFx3_ASAP7_75t_L g1621 ( .A(n_1536), .Y(n_1621) );
BUFx6f_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
OR2x2_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1539), .Y(n_1537) );
OR2x2_ASAP7_75t_L g1546 ( .A(n_1538), .B(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1538), .Y(n_1566) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1539), .Y(n_1565) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1542), .Y(n_1539) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1542), .Y(n_1553) );
XOR2x2_ASAP7_75t_L g1767 ( .A(n_1543), .B(n_1768), .Y(n_1767) );
HB1xp67_ASAP7_75t_L g1622 ( .A(n_1544), .Y(n_1622) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1547), .Y(n_1568) );
OAI22xp5_ASAP7_75t_L g1549 ( .A1(n_1550), .A2(n_1555), .B1(n_1556), .B2(n_1558), .Y(n_1549) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
BUFx3_ASAP7_75t_L g1618 ( .A(n_1551), .Y(n_1618) );
AND2x4_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1554), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1552), .B(n_1554), .Y(n_1575) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
AND2x4_ASAP7_75t_L g1557 ( .A(n_1553), .B(n_1554), .Y(n_1557) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1556), .Y(n_1617) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
OR2x2_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1570), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1560), .B(n_1587), .Y(n_1586) );
OAI321xp33_ASAP7_75t_SL g1671 ( .A1(n_1560), .A2(n_1672), .A3(n_1673), .B1(n_1674), .B2(n_1675), .C(n_1677), .Y(n_1671) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_1560), .B(n_1602), .Y(n_1683) );
INVx2_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1561), .B(n_1576), .Y(n_1670) );
NAND2xp5_ASAP7_75t_SL g1705 ( .A(n_1561), .B(n_1706), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1561), .B(n_1634), .Y(n_1736) );
BUFx2_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1562), .B(n_1599), .Y(n_1598) );
INVx2_ASAP7_75t_L g1606 ( .A(n_1562), .Y(n_1606) );
NAND2xp5_ASAP7_75t_L g1626 ( .A(n_1562), .B(n_1627), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1644 ( .A(n_1562), .B(n_1632), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1562), .B(n_1588), .Y(n_1663) );
INVx2_ASAP7_75t_L g1680 ( .A(n_1562), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1569), .Y(n_1562) );
AND2x4_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1566), .Y(n_1564) );
OAI21xp33_ASAP7_75t_SL g1909 ( .A1(n_1565), .A2(n_1907), .B(n_1910), .Y(n_1909) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_1566), .B(n_1568), .Y(n_1567) );
BUFx2_ASAP7_75t_L g1656 ( .A(n_1567), .Y(n_1656) );
INVx2_ASAP7_75t_L g1611 ( .A(n_1570), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1576), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1571), .B(n_1598), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1571), .B(n_1608), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1571), .B(n_1603), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1571), .B(n_1613), .Y(n_1633) );
INVxp67_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
BUFx2_ASAP7_75t_L g1588 ( .A(n_1572), .Y(n_1588) );
BUFx3_ASAP7_75t_L g1632 ( .A(n_1572), .Y(n_1632) );
OR2x2_ASAP7_75t_L g1716 ( .A(n_1572), .B(n_1581), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1573), .B(n_1574), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1576), .B(n_1632), .Y(n_1631) );
NOR2xp33_ASAP7_75t_L g1714 ( .A(n_1576), .B(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1576), .Y(n_1725) );
NAND3xp33_ASAP7_75t_SL g1743 ( .A(n_1576), .B(n_1605), .C(n_1667), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1580), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1577), .B(n_1581), .Y(n_1599) );
INVx2_ASAP7_75t_L g1604 ( .A(n_1577), .Y(n_1604) );
OR2x2_ASAP7_75t_L g1609 ( .A(n_1577), .B(n_1581), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1577), .B(n_1632), .Y(n_1678) );
NOR2xp33_ASAP7_75t_L g1706 ( .A(n_1577), .B(n_1632), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1579), .Y(n_1577) );
NOR2x1_ASAP7_75t_L g1587 ( .A(n_1580), .B(n_1588), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1580), .B(n_1632), .Y(n_1729) );
INVx2_ASAP7_75t_SL g1580 ( .A(n_1581), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1581), .B(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
NOR2xp33_ASAP7_75t_L g1741 ( .A(n_1586), .B(n_1688), .Y(n_1741) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1587), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1588), .B(n_1603), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1588), .B(n_1599), .Y(n_1650) );
A2O1A1Ixp33_ASAP7_75t_L g1595 ( .A1(n_1589), .A2(n_1596), .B(n_1600), .C(n_1601), .Y(n_1595) );
OAI221xp5_ASAP7_75t_L g1635 ( .A1(n_1589), .A2(n_1590), .B1(n_1636), .B2(n_1638), .C(n_1640), .Y(n_1635) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g1745 ( .A1(n_1590), .A2(n_1624), .B1(n_1686), .B2(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1591), .B(n_1654), .Y(n_1676) );
OR2x2_ASAP7_75t_L g1688 ( .A(n_1591), .B(n_1689), .Y(n_1688) );
INVx3_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
OR2x2_ASAP7_75t_L g1712 ( .A(n_1592), .B(n_1654), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1753 ( .A(n_1592), .B(n_1653), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1594), .Y(n_1592) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1598), .Y(n_1674) );
O2A1O1Ixp33_ASAP7_75t_L g1731 ( .A1(n_1598), .A2(n_1732), .B(n_1733), .C(n_1734), .Y(n_1731) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1599), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1599), .B(n_1606), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1605 ( .A(n_1600), .B(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1600), .Y(n_1625) );
NOR2xp33_ASAP7_75t_L g1642 ( .A(n_1600), .B(n_1643), .Y(n_1642) );
NOR2xp33_ASAP7_75t_L g1702 ( .A(n_1600), .B(n_1688), .Y(n_1702) );
INVx2_ASAP7_75t_L g1710 ( .A(n_1600), .Y(n_1710) );
AOI21xp33_ASAP7_75t_SL g1601 ( .A1(n_1602), .A2(n_1605), .B(n_1607), .Y(n_1601) );
OAI211xp5_ASAP7_75t_L g1699 ( .A1(n_1602), .A2(n_1680), .B(n_1686), .C(n_1700), .Y(n_1699) );
A2O1A1Ixp33_ASAP7_75t_SL g1744 ( .A1(n_1602), .A2(n_1718), .B(n_1745), .C(n_1750), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1603), .B(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1603), .Y(n_1694) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1604), .B(n_1632), .Y(n_1672) );
OAI321xp33_ASAP7_75t_L g1734 ( .A1(n_1604), .A2(n_1723), .A3(n_1735), .B1(n_1737), .B2(n_1738), .C(n_1740), .Y(n_1734) );
NOR2xp33_ASAP7_75t_L g1608 ( .A(n_1606), .B(n_1609), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1606), .B(n_1613), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1606), .B(n_1678), .Y(n_1739) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1607), .Y(n_1749) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1609), .Y(n_1613) );
OR2x2_ASAP7_75t_L g1643 ( .A(n_1609), .B(n_1644), .Y(n_1643) );
NOR2xp33_ASAP7_75t_L g1684 ( .A(n_1609), .B(n_1685), .Y(n_1684) );
O2A1O1Ixp33_ASAP7_75t_L g1610 ( .A1(n_1611), .A2(n_1612), .B(n_1614), .C(n_1615), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1612), .B(n_1632), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1613), .B(n_1663), .Y(n_1711) );
CKINVDCx5p33_ASAP7_75t_R g1668 ( .A(n_1614), .Y(n_1668) );
AOI211xp5_ASAP7_75t_SL g1681 ( .A1(n_1614), .A2(n_1682), .B(n_1684), .C(n_1687), .Y(n_1681) );
NAND4xp25_ASAP7_75t_L g1761 ( .A(n_1614), .B(n_1663), .C(n_1700), .D(n_1762), .Y(n_1761) );
INVx3_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx3_ASAP7_75t_L g1640 ( .A(n_1616), .Y(n_1640) );
A2O1A1Ixp33_ASAP7_75t_SL g1658 ( .A1(n_1616), .A2(n_1659), .B(n_1681), .C(n_1697), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1616), .B(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1621), .Y(n_1765) );
NAND4xp25_ASAP7_75t_L g1623 ( .A(n_1624), .B(n_1628), .C(n_1641), .D(n_1645), .Y(n_1623) );
OR2x2_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1626), .Y(n_1624) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1626), .Y(n_1752) );
AOI21xp33_ASAP7_75t_L g1628 ( .A1(n_1629), .A2(n_1634), .B(n_1635), .Y(n_1628) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
NOR2xp33_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1633), .Y(n_1630) );
OR2x2_ASAP7_75t_L g1636 ( .A(n_1632), .B(n_1637), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1632), .B(n_1639), .Y(n_1691) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1633), .Y(n_1722) );
AOI221xp5_ASAP7_75t_L g1659 ( .A1(n_1634), .A2(n_1660), .B1(n_1664), .B2(n_1669), .C(n_1671), .Y(n_1659) );
AOI21xp5_ASAP7_75t_L g1750 ( .A1(n_1634), .A2(n_1648), .B(n_1690), .Y(n_1750) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1636), .Y(n_1707) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1640), .B(n_1652), .Y(n_1651) );
O2A1O1Ixp33_ASAP7_75t_L g1708 ( .A1(n_1640), .A2(n_1670), .B(n_1709), .C(n_1712), .Y(n_1708) );
OAI211xp5_ASAP7_75t_L g1730 ( .A1(n_1640), .A2(n_1731), .B(n_1744), .C(n_1751), .Y(n_1730) );
INVxp67_ASAP7_75t_SL g1641 ( .A(n_1642), .Y(n_1641) );
O2A1O1Ixp33_ASAP7_75t_L g1751 ( .A1(n_1642), .A2(n_1752), .B(n_1753), .C(n_1754), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1643), .B(n_1661), .Y(n_1660) );
NOR2xp33_ASAP7_75t_L g1760 ( .A(n_1643), .B(n_1748), .Y(n_1760) );
OR2x2_ASAP7_75t_L g1724 ( .A(n_1644), .B(n_1725), .Y(n_1724) );
INVxp67_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
NOR2xp33_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1649), .Y(n_1646) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1648), .B(n_1652), .Y(n_1696) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
OAI332xp33_ASAP7_75t_L g1713 ( .A1(n_1651), .A2(n_1710), .A3(n_1714), .B1(n_1717), .B2(n_1720), .B3(n_1722), .C1(n_1723), .C2(n_1724), .Y(n_1713) );
INVx2_ASAP7_75t_L g1700 ( .A(n_1652), .Y(n_1700) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1653), .Y(n_1667) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1654), .Y(n_1689) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1654), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1657), .Y(n_1654) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1662), .B(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
OR2x2_ASAP7_75t_L g1665 ( .A(n_1666), .B(n_1668), .Y(n_1665) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1667), .Y(n_1719) );
AOI211xp5_ASAP7_75t_L g1726 ( .A1(n_1667), .A2(n_1685), .B(n_1727), .C(n_1728), .Y(n_1726) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1673), .Y(n_1733) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1676), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1679), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_1680), .B(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
OAI21xp33_ASAP7_75t_L g1687 ( .A1(n_1688), .A2(n_1690), .B(n_1692), .Y(n_1687) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVxp33_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
NOR2xp33_ASAP7_75t_L g1693 ( .A(n_1694), .B(n_1695), .Y(n_1693) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1694), .B(n_1725), .Y(n_1763) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
OAI21xp5_ASAP7_75t_L g1703 ( .A1(n_1696), .A2(n_1704), .B(n_1707), .Y(n_1703) );
NOR4xp25_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1708), .C(n_1713), .D(n_1726), .Y(n_1697) );
NAND3xp33_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1701), .C(n_1703), .Y(n_1698) );
A2O1A1Ixp33_ASAP7_75t_L g1754 ( .A1(n_1700), .A2(n_1755), .B(n_1759), .C(n_1761), .Y(n_1754) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1711), .Y(n_1709) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
INVxp67_ASAP7_75t_L g1758 ( .A(n_1724), .Y(n_1758) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
NOR2xp33_ASAP7_75t_L g1740 ( .A(n_1741), .B(n_1742), .Y(n_1740) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVxp33_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
NOR2xp33_ASAP7_75t_L g1747 ( .A(n_1748), .B(n_1749), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_1756), .B(n_1758), .Y(n_1755) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx2_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
NAND2xp5_ASAP7_75t_L g1768 ( .A(n_1769), .B(n_1804), .Y(n_1768) );
AND4x1_ASAP7_75t_L g1769 ( .A(n_1770), .B(n_1780), .C(n_1788), .D(n_1795), .Y(n_1769) );
AOI221xp5_ASAP7_75t_L g1770 ( .A1(n_1771), .A2(n_1776), .B1(n_1777), .B2(n_1778), .C(n_1779), .Y(n_1770) );
AND2x4_ASAP7_75t_L g1771 ( .A(n_1772), .B(n_1773), .Y(n_1771) );
INVx3_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
AOI22xp33_ASAP7_75t_L g1780 ( .A1(n_1781), .A2(n_1782), .B1(n_1785), .B2(n_1786), .Y(n_1780) );
BUFx2_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
AOI22xp33_ASAP7_75t_L g1788 ( .A1(n_1789), .A2(n_1790), .B1(n_1792), .B2(n_1793), .Y(n_1788) );
BUFx2_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
BUFx2_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
AOI21xp5_ASAP7_75t_L g1804 ( .A1(n_1805), .A2(n_1814), .B(n_1815), .Y(n_1804) );
INVx2_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
AND2x4_ASAP7_75t_L g1806 ( .A(n_1807), .B(n_1808), .Y(n_1806) );
INVx2_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
AND2x4_ASAP7_75t_L g1823 ( .A(n_1811), .B(n_1824), .Y(n_1823) );
AND2x2_ASAP7_75t_L g1827 ( .A(n_1811), .B(n_1828), .Y(n_1827) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1811), .Y(n_1847) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
AOI31xp33_ASAP7_75t_L g1815 ( .A1(n_1816), .A2(n_1833), .A3(n_1848), .B(n_1855), .Y(n_1815) );
AOI211xp5_ASAP7_75t_L g1816 ( .A1(n_1817), .A2(n_1818), .B(n_1821), .C(n_1829), .Y(n_1816) );
INVx2_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
INVx2_ASAP7_75t_SL g1822 ( .A(n_1823), .Y(n_1822) );
INVx2_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx3_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
AOI221xp5_ASAP7_75t_L g1833 ( .A1(n_1834), .A2(n_1836), .B1(n_1837), .B2(n_1843), .C(n_1845), .Y(n_1833) );
HB1xp67_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_SL g1846 ( .A(n_1847), .Y(n_1846) );
AOI22xp33_ASAP7_75t_L g1848 ( .A1(n_1849), .A2(n_1850), .B1(n_1852), .B2(n_1853), .Y(n_1848) );
INVx6_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
INVx4_ASAP7_75t_L g1853 ( .A(n_1854), .Y(n_1853) );
CKINVDCx14_ASAP7_75t_R g1856 ( .A(n_1857), .Y(n_1856) );
INVx4_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1860), .Y(n_1859) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1861), .Y(n_1860) );
INVxp33_ASAP7_75t_L g1863 ( .A(n_1864), .Y(n_1863) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
HB1xp67_ASAP7_75t_L g1867 ( .A(n_1868), .Y(n_1867) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1869), .Y(n_1868) );
NAND2xp5_ASAP7_75t_L g1882 ( .A(n_1883), .B(n_1889), .Y(n_1882) );
INVx1_ASAP7_75t_L g1904 ( .A(n_1905), .Y(n_1904) );
CKINVDCx5p33_ASAP7_75t_R g1905 ( .A(n_1906), .Y(n_1905) );
HB1xp67_ASAP7_75t_L g1908 ( .A(n_1909), .Y(n_1908) );
endmodule