module fake_netlist_1_8253_n_812 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_812);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_812;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_808;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_476;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g95 ( .A(n_79), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_60), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_18), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_52), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_82), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_30), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_57), .Y(n_102) );
BUFx8_ASAP7_75t_SL g103 ( .A(n_39), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_92), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_85), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_94), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_48), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_40), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_10), .Y(n_113) );
BUFx10_ASAP7_75t_L g114 ( .A(n_58), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_65), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_44), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_66), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_56), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_44), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_68), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_70), .Y(n_121) );
BUFx10_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_14), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_91), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_31), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_86), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_0), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_74), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_32), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_64), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_53), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_69), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_29), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_24), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_18), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_59), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_51), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_5), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_28), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_106), .B(n_129), .Y(n_141) );
NOR2x1_ASAP7_75t_L g142 ( .A(n_135), .B(n_0), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_129), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_135), .Y(n_144) );
BUFx2_ASAP7_75t_L g145 ( .A(n_106), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_106), .B(n_1), .Y(n_146) );
INVx2_ASAP7_75t_SL g147 ( .A(n_114), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_135), .B(n_133), .Y(n_148) );
BUFx12f_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_95), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_97), .Y(n_153) );
CKINVDCx11_ASAP7_75t_R g154 ( .A(n_122), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_97), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_109), .B(n_1), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_108), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_135), .B(n_2), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_135), .B(n_2), .Y(n_159) );
BUFx8_ASAP7_75t_SL g160 ( .A(n_103), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_133), .B(n_3), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_133), .B(n_3), .Y(n_162) );
INVx5_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
OAI22xp33_ASAP7_75t_R g164 ( .A1(n_146), .A2(n_134), .B1(n_125), .B2(n_119), .Y(n_164) );
AO22x2_ASAP7_75t_L g165 ( .A1(n_141), .A2(n_125), .B1(n_119), .B2(n_134), .Y(n_165) );
AO22x2_ASAP7_75t_L g166 ( .A1(n_141), .A2(n_137), .B1(n_96), .B2(n_128), .Y(n_166) );
BUFx10_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_150), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_140), .A2(n_95), .B1(n_109), .B2(n_132), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_145), .B(n_122), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_140), .A2(n_132), .B1(n_138), .B2(n_98), .Y(n_174) );
OAI22xp33_ASAP7_75t_SL g175 ( .A1(n_141), .A2(n_139), .B1(n_101), .B2(n_116), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_143), .A2(n_113), .B1(n_127), .B2(n_110), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_151), .B(n_96), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
OAI22xp5_ASAP7_75t_SL g180 ( .A1(n_152), .A2(n_112), .B1(n_123), .B2(n_103), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_143), .A2(n_122), .B1(n_104), .B2(n_136), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_145), .A2(n_122), .B1(n_104), .B2(n_136), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_145), .A2(n_122), .B1(n_117), .B2(n_102), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_149), .A2(n_137), .B1(n_102), .B2(n_105), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_149), .A2(n_117), .B1(n_105), .B2(n_128), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_147), .B(n_107), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_149), .B(n_114), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_161), .A2(n_107), .B1(n_126), .B2(n_111), .Y(n_194) );
OAI22xp33_ASAP7_75t_SL g195 ( .A1(n_146), .A2(n_111), .B1(n_126), .B2(n_130), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_149), .B(n_114), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_154), .B(n_108), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_154), .A2(n_131), .B1(n_124), .B2(n_121), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_147), .A2(n_120), .B1(n_118), .B2(n_115), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_147), .A2(n_100), .B1(n_99), .B2(n_108), .Y(n_201) );
OR2x6_ASAP7_75t_L g202 ( .A(n_161), .B(n_99), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_147), .B(n_4), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_204) );
AO22x2_ASAP7_75t_L g205 ( .A1(n_161), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_151), .B(n_7), .Y(n_206) );
XNOR2xp5_ASAP7_75t_L g207 ( .A(n_160), .B(n_8), .Y(n_207) );
INVx1_ASAP7_75t_SL g208 ( .A(n_151), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_161), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_159), .A2(n_9), .B1(n_11), .B2(n_12), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_161), .A2(n_12), .B1(n_13), .B2(n_15), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_180), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_179), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_184), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_191), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_193), .B(n_151), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_198), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_209), .B(n_151), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_192), .B(n_151), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_179), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_208), .B(n_162), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_173), .B(n_148), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_167), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_187), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_167), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_171), .B(n_148), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_176), .B(n_148), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_174), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_202), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_190), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_166), .B(n_148), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_202), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_196), .B(n_156), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_208), .B(n_162), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_202), .Y(n_238) );
NAND2x1p5_ASAP7_75t_L g239 ( .A(n_203), .B(n_162), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_200), .B(n_156), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_206), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_170), .Y(n_242) );
XOR2xp5_ASAP7_75t_L g243 ( .A(n_207), .B(n_160), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_182), .B(n_162), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_177), .B(n_162), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_178), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_178), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_165), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_189), .A2(n_142), .B(n_162), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_165), .B(n_142), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_194), .B(n_155), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_165), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_194), .B(n_155), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_166), .B(n_142), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_189), .B(n_155), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_166), .B(n_155), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_205), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_205), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_183), .B(n_163), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_203), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_185), .B(n_163), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_199), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_204), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_212), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_211), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_211), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_197), .B(n_181), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_187), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_188), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_188), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_186), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_195), .B(n_163), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_169), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_169), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_201), .B(n_163), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_169), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_246), .A2(n_175), .B(n_163), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_234), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_215), .B(n_163), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_215), .B(n_163), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_216), .B(n_164), .Y(n_283) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_239), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_216), .B(n_163), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_218), .B(n_163), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_214), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_232), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_217), .Y(n_291) );
AND2x6_ASAP7_75t_L g292 ( .A(n_234), .B(n_150), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_232), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_245), .B(n_13), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_245), .B(n_15), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_246), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_247), .B(n_163), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_217), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_264), .B(n_16), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_234), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_219), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_247), .B(n_150), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_222), .B(n_169), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_219), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_256), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_250), .B(n_150), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_256), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_224), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_223), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_250), .B(n_150), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_278), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_224), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_235), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_254), .B(n_150), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_248), .B(n_153), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_248), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_254), .B(n_153), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_239), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_239), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_264), .B(n_16), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_214), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_221), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_223), .B(n_153), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_231), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_244), .B(n_153), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_231), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_267), .B(n_153), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_278), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_265), .B(n_153), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_297), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_297), .Y(n_335) );
AND2x6_ASAP7_75t_L g336 ( .A(n_294), .B(n_235), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_283), .B(n_265), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_292), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
INVx6_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_302), .B(n_266), .Y(n_341) );
OR2x6_ASAP7_75t_L g342 ( .A(n_313), .B(n_238), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_283), .B(n_242), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_302), .B(n_266), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_313), .B(n_284), .Y(n_347) );
OR2x6_ASAP7_75t_L g348 ( .A(n_313), .B(n_238), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_287), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_297), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_292), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_283), .B(n_269), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_301), .B(n_269), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_297), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_313), .B(n_228), .Y(n_356) );
NOR2xp33_ASAP7_75t_SL g357 ( .A(n_313), .B(n_222), .Y(n_357) );
INVx5_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_284), .B(n_228), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_287), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_297), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_279), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_302), .B(n_267), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_305), .B(n_268), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_301), .B(n_273), .Y(n_365) );
INVx6_ASAP7_75t_L g366 ( .A(n_297), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_285), .Y(n_367) );
INVx5_ASAP7_75t_L g368 ( .A(n_347), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_347), .B(n_321), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_347), .B(n_321), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_340), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
BUFx2_ASAP7_75t_SL g378 ( .A(n_358), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_363), .B(n_305), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_340), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_340), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_357), .A2(n_323), .B1(n_300), .B2(n_295), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_367), .Y(n_383) );
NOR2xp33_ASAP7_75t_SL g384 ( .A(n_357), .B(n_358), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_359), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_337), .A2(n_296), .B1(n_295), .B2(n_268), .Y(n_386) );
INVx4_ASAP7_75t_L g387 ( .A(n_358), .Y(n_387) );
BUFx12f_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
BUFx4_ASAP7_75t_R g389 ( .A(n_338), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_344), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_367), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_358), .B(n_321), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_358), .Y(n_395) );
INVx5_ASAP7_75t_L g396 ( .A(n_336), .Y(n_396) );
BUFx8_ASAP7_75t_L g397 ( .A(n_338), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_383), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_383), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_373), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_385), .A2(n_362), .B1(n_300), .B2(n_323), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_373), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_382), .A2(n_337), .B1(n_359), .B2(n_296), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_390), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_379), .B(n_363), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_388), .Y(n_406) );
INVx3_ASAP7_75t_SL g407 ( .A(n_396), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_386), .A2(n_359), .B1(n_343), .B2(n_365), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_382), .A2(n_359), .B1(n_323), .B2(n_300), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_385), .A2(n_356), .B1(n_338), .B2(n_258), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_368), .Y(n_413) );
OAI22xp33_ASAP7_75t_SL g414 ( .A1(n_369), .A2(n_258), .B1(n_257), .B2(n_259), .Y(n_414) );
CKINVDCx6p67_ASAP7_75t_R g415 ( .A(n_368), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_388), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_389), .Y(n_418) );
INVx6_ASAP7_75t_L g419 ( .A(n_368), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_394), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_370), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_368), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_368), .Y(n_423) );
BUFx12f_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_385), .A2(n_356), .B1(n_257), .B2(n_259), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_370), .Y(n_426) );
INVx6_ASAP7_75t_L g427 ( .A(n_368), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_391), .B(n_367), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_386), .A2(n_356), .B1(n_352), .B2(n_363), .Y(n_432) );
INVx4_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_368), .A2(n_356), .B1(n_352), .B2(n_308), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_391), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_374), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_368), .B(n_349), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_370), .A2(n_308), .B1(n_346), .B2(n_341), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_369), .Y(n_440) );
BUFx10_ASAP7_75t_L g441 ( .A(n_371), .Y(n_441) );
CKINVDCx11_ASAP7_75t_R g442 ( .A(n_371), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_403), .A2(n_371), .B1(n_292), .B2(n_308), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_398), .Y(n_444) );
OAI22xp33_ASAP7_75t_SL g445 ( .A1(n_417), .A2(n_369), .B1(n_384), .B2(n_379), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_401), .A2(n_369), .B1(n_396), .B2(n_371), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_410), .A2(n_432), .B1(n_409), .B2(n_418), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
AOI222xp33_ASAP7_75t_L g449 ( .A1(n_410), .A2(n_279), .B1(n_341), .B2(n_346), .C1(n_240), .C2(n_274), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_399), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_424), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_432), .A2(n_292), .B1(n_308), .B2(n_397), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_399), .B(n_369), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_399), .B(n_307), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_409), .A2(n_292), .B1(n_397), .B2(n_301), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_424), .A2(n_292), .B1(n_397), .B2(n_301), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_424), .A2(n_292), .B1(n_397), .B2(n_301), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_437), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_417), .B(n_213), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_436), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_442), .A2(n_292), .B1(n_397), .B2(n_301), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_402), .B(n_360), .Y(n_462) );
INVx5_ASAP7_75t_L g463 ( .A(n_406), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_439), .A2(n_249), .B1(n_230), .B2(n_280), .C1(n_291), .C2(n_299), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_436), .B(n_307), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_404), .B(n_360), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_404), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_415), .A2(n_292), .B1(n_397), .B2(n_353), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_436), .Y(n_469) );
OAI21xp5_ASAP7_75t_SL g470 ( .A1(n_406), .A2(n_243), .B(n_351), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_415), .A2(n_353), .B1(n_381), .B2(n_376), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_415), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_434), .A2(n_381), .B1(n_376), .B2(n_342), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_434), .A2(n_381), .B1(n_376), .B2(n_342), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_439), .A2(n_376), .B1(n_342), .B2(n_348), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_431), .B(n_307), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_412), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_440), .B(n_396), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_416), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_440), .Y(n_481) );
OAI222xp33_ASAP7_75t_L g482 ( .A1(n_413), .A2(n_396), .B1(n_372), .B2(n_380), .C1(n_342), .C2(n_348), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_408), .A2(n_342), .B1(n_348), .B2(n_375), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_429), .Y(n_484) );
INVx5_ASAP7_75t_L g485 ( .A(n_406), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_411), .A2(n_396), .B1(n_306), .B2(n_348), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_420), .B(n_364), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_440), .A2(n_396), .B1(n_378), .B2(n_384), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_431), .B(n_307), .Y(n_489) );
INVx4_ASAP7_75t_R g490 ( .A(n_413), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_420), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_416), .A2(n_304), .B(n_355), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_422), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_408), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_428), .B(n_364), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_429), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_431), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_437), .Y(n_499) );
OAI21xp5_ASAP7_75t_SL g500 ( .A1(n_406), .A2(n_243), .B(n_351), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_421), .Y(n_501) );
AOI222xp33_ASAP7_75t_L g502 ( .A1(n_405), .A2(n_249), .B1(n_299), .B2(n_291), .C1(n_316), .C2(n_236), .Y(n_502) );
INVx4_ASAP7_75t_L g503 ( .A(n_430), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
BUFx12f_ASAP7_75t_L g505 ( .A(n_441), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_411), .A2(n_425), .B1(n_423), .B2(n_430), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_426), .A2(n_375), .B1(n_393), .B2(n_321), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_419), .A2(n_378), .B1(n_392), .B2(n_393), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_447), .A2(n_426), .B1(n_438), .B2(n_419), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_506), .A2(n_438), .B1(n_419), .B2(n_427), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_464), .A2(n_438), .B1(n_419), .B2(n_427), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_505), .A2(n_419), .B1(n_427), .B2(n_422), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_449), .A2(n_446), .B1(n_455), .B2(n_502), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_453), .B(n_437), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_486), .A2(n_427), .B1(n_419), .B2(n_422), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_443), .A2(n_427), .B1(n_441), .B2(n_425), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_448), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_452), .A2(n_441), .B1(n_435), .B2(n_430), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_468), .A2(n_435), .B1(n_407), .B2(n_433), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_476), .A2(n_441), .B1(n_435), .B2(n_375), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_470), .A2(n_414), .B1(n_299), .B2(n_291), .C(n_263), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_505), .A2(n_433), .B1(n_378), .B2(n_392), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_463), .B(n_485), .C(n_503), .Y(n_524) );
OAI222xp33_ASAP7_75t_L g525 ( .A1(n_494), .A2(n_433), .B1(n_372), .B2(n_387), .C1(n_395), .C2(n_393), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_473), .A2(n_375), .B1(n_393), .B2(n_407), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_448), .B(n_414), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_445), .B(n_407), .Y(n_528) );
AOI222xp33_ASAP7_75t_L g529 ( .A1(n_500), .A2(n_316), .B1(n_333), .B2(n_328), .C1(n_320), .C2(n_311), .Y(n_529) );
OAI222xp33_ASAP7_75t_L g530 ( .A1(n_494), .A2(n_387), .B1(n_395), .B2(n_225), .C1(n_227), .C2(n_389), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_503), .A2(n_387), .B1(n_395), .B2(n_437), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_475), .A2(n_310), .B1(n_311), .B2(n_320), .C(n_328), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_467), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_477), .A2(n_333), .B1(n_336), .B2(n_314), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_480), .A2(n_260), .B1(n_229), .B2(n_310), .C(n_153), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_477), .A2(n_336), .B1(n_309), .B2(n_314), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_489), .A2(n_336), .B1(n_309), .B2(n_327), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_483), .A2(n_322), .B1(n_309), .B2(n_329), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_463), .A2(n_437), .B1(n_336), .B2(n_374), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_474), .B(n_318), .Y(n_540) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_499), .A2(n_331), .B(n_304), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_489), .A2(n_336), .B1(n_329), .B2(n_330), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_450), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_461), .A2(n_336), .B1(n_318), .B2(n_330), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_463), .A2(n_377), .B1(n_374), .B2(n_366), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_478), .B(n_319), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_485), .A2(n_377), .B1(n_374), .B2(n_366), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_481), .A2(n_471), .B1(n_495), .B2(n_501), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_456), .A2(n_366), .B1(n_361), .B2(n_350), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_481), .A2(n_319), .B1(n_366), .B2(n_326), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_485), .A2(n_339), .B1(n_334), .B2(n_317), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_495), .A2(n_366), .B1(n_326), .B2(n_354), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g553 ( .A(n_459), .B(n_331), .C(n_253), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_457), .A2(n_361), .B1(n_354), .B2(n_350), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_501), .A2(n_326), .B1(n_335), .B2(n_354), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_485), .A2(n_361), .B1(n_354), .B2(n_350), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_485), .A2(n_345), .B1(n_335), .B2(n_354), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_485), .A2(n_345), .B1(n_335), .B2(n_354), .Y(n_558) );
OAI222xp33_ASAP7_75t_L g559 ( .A1(n_472), .A2(n_317), .B1(n_251), .B2(n_253), .C1(n_339), .C2(n_334), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_478), .B(n_17), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_453), .B(n_153), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_451), .A2(n_326), .B1(n_335), .B2(n_350), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_451), .A2(n_350), .B1(n_345), .B2(n_281), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_444), .A2(n_345), .B1(n_281), .B2(n_315), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g565 ( .A1(n_491), .A2(n_229), .B1(n_260), .B2(n_261), .C1(n_303), .C2(n_281), .Y(n_565) );
OAI222xp33_ASAP7_75t_L g566 ( .A1(n_508), .A2(n_317), .B1(n_334), .B2(n_339), .C1(n_286), .C2(n_282), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_454), .A2(n_298), .B1(n_281), .B2(n_261), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_484), .B(n_374), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_479), .A2(n_377), .B1(n_374), .B2(n_298), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_507), .A2(n_262), .B1(n_277), .B2(n_241), .C(n_282), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_454), .A2(n_315), .B1(n_241), .B2(n_374), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_479), .A2(n_377), .B1(n_298), .B2(n_317), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_465), .A2(n_315), .B1(n_377), .B2(n_294), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_488), .A2(n_377), .B1(n_290), .B2(n_293), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_487), .A2(n_377), .B1(n_290), .B2(n_294), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_465), .A2(n_315), .B1(n_294), .B2(n_303), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_491), .B(n_17), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_479), .A2(n_315), .B1(n_303), .B2(n_298), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_479), .A2(n_153), .B1(n_157), .B2(n_286), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_492), .B(n_19), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_498), .A2(n_157), .B1(n_288), .B2(n_233), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_498), .A2(n_157), .B1(n_288), .B2(n_233), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_497), .A2(n_157), .B1(n_277), .B2(n_262), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_497), .A2(n_157), .B1(n_220), .B2(n_324), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_492), .B(n_20), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_484), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_482), .B(n_21), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_496), .A2(n_462), .B1(n_466), .B2(n_460), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_460), .A2(n_157), .B1(n_325), .B2(n_324), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_469), .A2(n_157), .B1(n_325), .B2(n_324), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_469), .B(n_21), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_493), .A2(n_325), .B1(n_324), .B2(n_289), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_499), .A2(n_157), .B1(n_325), .B2(n_289), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_588), .B(n_504), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_513), .A2(n_504), .B1(n_458), .B2(n_490), .C(n_237), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_522), .A2(n_458), .B1(n_490), .B2(n_289), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_587), .B(n_458), .C(n_285), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_510), .A2(n_458), .B(n_289), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_527), .B(n_22), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g601 ( .A1(n_524), .A2(n_237), .B(n_23), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_524), .B(n_285), .C(n_275), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_514), .B(n_22), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_518), .B(n_23), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_509), .A2(n_285), .B1(n_25), .B2(n_26), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_533), .B(n_24), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_533), .B(n_25), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_586), .B(n_26), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_548), .B(n_276), .C(n_275), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_517), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_610) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_511), .B(n_27), .C(n_30), .D(n_31), .Y(n_611) );
OAI221xp5_ASAP7_75t_SL g612 ( .A1(n_521), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_560), .B(n_33), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_577), .B(n_35), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_553), .A2(n_36), .B1(n_37), .B2(n_38), .C(n_39), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_561), .B(n_37), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_561), .B(n_38), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_586), .B(n_41), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_580), .B(n_276), .C(n_255), .Y(n_619) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_516), .B(n_41), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_585), .B(n_255), .C(n_271), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_543), .B(n_42), .Y(n_622) );
OAI221xp5_ASAP7_75t_SL g623 ( .A1(n_519), .A2(n_42), .B1(n_43), .B2(n_45), .C(n_46), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_574), .B(n_270), .C(n_332), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_591), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_568), .B(n_47), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_516), .B(n_332), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_568), .B(n_49), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g629 ( .A(n_529), .B(n_272), .C(n_226), .D(n_221), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_516), .B(n_50), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_529), .A2(n_332), .B1(n_312), .B2(n_55), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_540), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g633 ( .A1(n_530), .A2(n_54), .B(n_61), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_546), .B(n_63), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_526), .A2(n_332), .B1(n_312), .B2(n_72), .C(n_75), .Y(n_635) );
AOI21xp5_ASAP7_75t_SL g636 ( .A1(n_528), .A2(n_67), .B(n_71), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_525), .A2(n_76), .B(n_77), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_515), .B(n_78), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_512), .A2(n_80), .B(n_81), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_538), .B(n_83), .Y(n_640) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_523), .A2(n_84), .B(n_87), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_538), .B(n_89), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_532), .A2(n_565), .B1(n_535), .B2(n_570), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_531), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_541), .B(n_90), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_569), .B(n_93), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_565), .A2(n_312), .B1(n_332), .B2(n_536), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_537), .A2(n_312), .B1(n_332), .B2(n_542), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_555), .B(n_312), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_539), .A2(n_312), .B1(n_332), .B2(n_544), .C(n_572), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_545), .B(n_332), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_552), .B(n_550), .Y(n_652) );
NAND3xp33_ASAP7_75t_SL g653 ( .A(n_547), .B(n_520), .C(n_534), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_564), .B(n_575), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_592), .B(n_567), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_567), .B(n_571), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_563), .B(n_562), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_566), .B(n_559), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_551), .B(n_554), .Y(n_659) );
NOR3xp33_ASAP7_75t_SL g660 ( .A(n_549), .B(n_558), .C(n_551), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_579), .B(n_584), .C(n_582), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_593), .B(n_590), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g663 ( .A1(n_573), .A2(n_578), .B(n_576), .Y(n_663) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_556), .A2(n_581), .B(n_557), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_583), .B(n_587), .C(n_513), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_589), .B(n_588), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_587), .B(n_513), .C(n_524), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_587), .B(n_513), .C(n_524), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_667), .B(n_668), .C(n_644), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_601), .B(n_660), .C(n_658), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_620), .B(n_658), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_665), .A2(n_620), .B1(n_653), .B2(n_629), .Y(n_672) );
NAND4xp75_ASAP7_75t_L g673 ( .A(n_603), .B(n_659), .C(n_594), .D(n_666), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_600), .B(n_595), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_637), .B(n_598), .C(n_633), .Y(n_675) );
NAND4xp75_ASAP7_75t_L g676 ( .A(n_604), .B(n_654), .C(n_638), .D(n_608), .Y(n_676) );
NAND2x1_ASAP7_75t_L g677 ( .A(n_636), .B(n_602), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_613), .B(n_614), .C(n_641), .Y(n_678) );
XOR2xp5_ASAP7_75t_L g679 ( .A(n_652), .B(n_611), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_627), .B(n_626), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_606), .B(n_607), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_622), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_663), .B(n_657), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_627), .B(n_599), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_613), .A2(n_614), .B1(n_612), .B2(n_610), .C(n_615), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_643), .A2(n_656), .B1(n_631), .B2(n_655), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_618), .B(n_617), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_643), .A2(n_605), .B1(n_616), .B2(n_623), .C(n_650), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_630), .B(n_628), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_664), .B(n_639), .C(n_609), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_645), .B(n_624), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_647), .A2(n_596), .B1(n_661), .B2(n_662), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_621), .A2(n_648), .B1(n_619), .B2(n_642), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_635), .B(n_634), .C(n_640), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_651), .B(n_646), .Y(n_695) );
NAND4xp75_ASAP7_75t_L g696 ( .A(n_649), .B(n_620), .C(n_658), .D(n_644), .Y(n_696) );
OAI211xp5_ASAP7_75t_SL g697 ( .A1(n_667), .A2(n_668), .B(n_601), .C(n_644), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_620), .B(n_524), .Y(n_698) );
NAND2x1_ASAP7_75t_L g699 ( .A(n_660), .B(n_516), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_668), .B(n_667), .Y(n_700) );
CKINVDCx14_ASAP7_75t_R g701 ( .A(n_603), .Y(n_701) );
NAND4xp75_ASAP7_75t_L g702 ( .A(n_620), .B(n_658), .C(n_644), .D(n_660), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_667), .B(n_668), .C(n_644), .Y(n_703) );
NAND3xp33_ASAP7_75t_SL g704 ( .A(n_633), .B(n_601), .C(n_637), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_620), .B(n_524), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_667), .B(n_668), .C(n_644), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_597), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_632), .B(n_625), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_632), .B(n_625), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_667), .B(n_668), .C(n_644), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_601), .B(n_611), .C(n_612), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_601), .B(n_611), .C(n_612), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_667), .A2(n_668), .B1(n_665), .B2(n_620), .Y(n_713) );
NOR2x1_ASAP7_75t_L g714 ( .A(n_601), .B(n_524), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_601), .A2(n_633), .B(n_637), .C(n_667), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_601), .A2(n_633), .B(n_637), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g717 ( .A(n_601), .B(n_611), .C(n_612), .Y(n_717) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_673), .B(n_702), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_714), .A2(n_690), .B(n_670), .Y(n_719) );
BUFx2_ASAP7_75t_L g720 ( .A(n_701), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_707), .Y(n_721) );
INVx5_ASAP7_75t_L g722 ( .A(n_680), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_701), .Y(n_723) );
BUFx2_ASAP7_75t_L g724 ( .A(n_680), .Y(n_724) );
XNOR2xp5_ASAP7_75t_L g725 ( .A(n_713), .B(n_679), .Y(n_725) );
XNOR2x2_ASAP7_75t_L g726 ( .A(n_698), .B(n_705), .Y(n_726) );
XOR2x2_ASAP7_75t_L g727 ( .A(n_671), .B(n_696), .Y(n_727) );
XOR2x2_ASAP7_75t_L g728 ( .A(n_671), .B(n_676), .Y(n_728) );
NAND4xp75_ASAP7_75t_L g729 ( .A(n_672), .B(n_716), .C(n_705), .D(n_698), .Y(n_729) );
NAND4xp75_ASAP7_75t_L g730 ( .A(n_700), .B(n_683), .C(n_688), .D(n_685), .Y(n_730) );
XNOR2x2_ASAP7_75t_L g731 ( .A(n_704), .B(n_678), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_708), .B(n_709), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_683), .B(n_700), .Y(n_733) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_682), .Y(n_734) );
INVx3_ASAP7_75t_L g735 ( .A(n_699), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_689), .Y(n_736) );
NAND4xp75_ASAP7_75t_L g737 ( .A(n_674), .B(n_693), .C(n_684), .D(n_681), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_674), .Y(n_738) );
AND4x1_ASAP7_75t_L g739 ( .A(n_675), .B(n_717), .C(n_712), .D(n_711), .Y(n_739) );
NAND4xp75_ASAP7_75t_L g740 ( .A(n_684), .B(n_691), .C(n_697), .D(n_695), .Y(n_740) );
NAND4xp75_ASAP7_75t_L g741 ( .A(n_715), .B(n_669), .C(n_710), .D(n_706), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_703), .Y(n_742) );
XNOR2xp5_ASAP7_75t_L g743 ( .A(n_686), .B(n_692), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_677), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_720), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_734), .Y(n_746) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_729), .B(n_720), .Y(n_747) );
XOR2x2_ASAP7_75t_L g748 ( .A(n_730), .B(n_717), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_723), .Y(n_749) );
XNOR2x1_ASAP7_75t_L g750 ( .A(n_730), .B(n_743), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_721), .Y(n_751) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_718), .B(n_686), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_731), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_739), .B(n_692), .Y(n_754) );
INVxp67_ASAP7_75t_L g755 ( .A(n_731), .Y(n_755) );
XOR2x2_ASAP7_75t_L g756 ( .A(n_739), .B(n_712), .Y(n_756) );
OAI22x1_ASAP7_75t_L g757 ( .A1(n_725), .A2(n_743), .B1(n_742), .B2(n_744), .Y(n_757) );
INVxp67_ASAP7_75t_L g758 ( .A(n_733), .Y(n_758) );
INVx1_ASAP7_75t_SL g759 ( .A(n_732), .Y(n_759) );
XOR2x2_ASAP7_75t_L g760 ( .A(n_725), .B(n_711), .Y(n_760) );
XNOR2xp5_ASAP7_75t_L g761 ( .A(n_718), .B(n_687), .Y(n_761) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_726), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_735), .B(n_694), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_722), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_738), .Y(n_765) );
INVx2_ASAP7_75t_SL g766 ( .A(n_749), .Y(n_766) );
AO22x2_ASAP7_75t_L g767 ( .A1(n_750), .A2(n_729), .B1(n_741), .B2(n_737), .Y(n_767) );
OA22x2_ASAP7_75t_L g768 ( .A1(n_757), .A2(n_719), .B1(n_744), .B2(n_726), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_749), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_754), .A2(n_727), .B1(n_718), .B2(n_728), .Y(n_770) );
XNOR2x1_ASAP7_75t_L g771 ( .A(n_756), .B(n_727), .Y(n_771) );
AOI22x1_ASAP7_75t_L g772 ( .A1(n_762), .A2(n_719), .B1(n_735), .B2(n_727), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_745), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_747), .A2(n_741), .B1(n_740), .B2(n_724), .Y(n_774) );
INVx3_ASAP7_75t_L g775 ( .A(n_764), .Y(n_775) );
INVxp67_ASAP7_75t_L g776 ( .A(n_754), .Y(n_776) );
OA22x2_ASAP7_75t_L g777 ( .A1(n_753), .A2(n_735), .B1(n_736), .B2(n_728), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_751), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_773), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_778), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_769), .Y(n_781) );
CKINVDCx16_ASAP7_75t_R g782 ( .A(n_770), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_766), .Y(n_783) );
OAI322xp33_ASAP7_75t_L g784 ( .A1(n_768), .A2(n_755), .A3(n_750), .B1(n_752), .B2(n_758), .C1(n_761), .C2(n_759), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_766), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_775), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_776), .Y(n_787) );
AO22x1_ASAP7_75t_L g788 ( .A1(n_787), .A2(n_774), .B1(n_763), .B2(n_768), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_782), .A2(n_767), .B1(n_771), .B2(n_777), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_779), .Y(n_790) );
NAND4xp75_ASAP7_75t_SL g791 ( .A(n_784), .B(n_767), .C(n_777), .D(n_772), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_783), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_792), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_790), .Y(n_794) );
OAI31xp33_ASAP7_75t_L g795 ( .A1(n_791), .A2(n_771), .A3(n_767), .B(n_785), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g796 ( .A(n_795), .B(n_787), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_793), .B(n_760), .Y(n_797) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_793), .B(n_781), .Y(n_798) );
NOR2x1_ASAP7_75t_L g799 ( .A(n_796), .B(n_794), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_798), .Y(n_800) );
AND4x1_ASAP7_75t_L g801 ( .A(n_799), .B(n_789), .C(n_797), .D(n_756), .Y(n_801) );
AND4x1_ASAP7_75t_L g802 ( .A(n_800), .B(n_794), .C(n_748), .D(n_767), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_802), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_801), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_804), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_805), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_806), .A2(n_803), .B1(n_748), .B2(n_760), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_807), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_808), .A2(n_765), .B1(n_788), .B2(n_786), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_809), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_810), .A2(n_765), .B1(n_780), .B2(n_775), .C(n_763), .Y(n_811) );
AOI211xp5_ASAP7_75t_L g812 ( .A1(n_811), .A2(n_780), .B(n_746), .C(n_763), .Y(n_812) );
endmodule