module real_aes_8221_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_0), .Y(n_770) );
INVx1_ASAP7_75t_L g112 ( .A(n_1), .Y(n_112) );
INVx1_ASAP7_75t_L g465 ( .A(n_2), .Y(n_465) );
INVx1_ASAP7_75t_L g193 ( .A(n_3), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_4), .A2(n_38), .B1(n_154), .B2(n_495), .Y(n_510) );
AOI21xp33_ASAP7_75t_L g161 ( .A1(n_5), .A2(n_135), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_6), .B(n_128), .Y(n_478) );
AND2x6_ASAP7_75t_L g140 ( .A(n_7), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_8), .A2(n_243), .B(n_244), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_9), .B(n_39), .Y(n_113) );
INVx1_ASAP7_75t_L g168 ( .A(n_10), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_11), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
INVx1_ASAP7_75t_L g459 ( .A(n_13), .Y(n_459) );
INVx1_ASAP7_75t_L g249 ( .A(n_14), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_15), .B(n_176), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_16), .B(n_129), .Y(n_536) );
AO32x2_ASAP7_75t_L g508 ( .A1(n_17), .A2(n_128), .A3(n_173), .B1(n_487), .B2(n_509), .Y(n_508) );
OAI22xp5_ASAP7_75t_SL g761 ( .A1(n_18), .A2(n_62), .B1(n_762), .B2(n_763), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_18), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_19), .B(n_154), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_20), .B(n_149), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_21), .B(n_129), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_22), .A2(n_50), .B1(n_154), .B2(n_495), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_23), .B(n_135), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_24), .A2(n_76), .B1(n_154), .B2(n_176), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_25), .B(n_154), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_26), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_27), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_29), .B(n_170), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_30), .B(n_166), .Y(n_195) );
INVx1_ASAP7_75t_L g182 ( .A(n_31), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_32), .B(n_170), .Y(n_525) );
INVx2_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_34), .B(n_154), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_35), .B(n_170), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_36), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_37), .A2(n_140), .B(n_144), .C(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g180 ( .A(n_40), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_41), .B(n_166), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_42), .B(n_154), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_43), .A2(n_86), .B1(n_212), .B2(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_44), .B(n_154), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_45), .B(n_154), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_46), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_47), .A2(n_69), .B1(n_739), .B2(n_740), .Y(n_738) );
CKINVDCx16_ASAP7_75t_R g740 ( .A(n_47), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_48), .B(n_464), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_49), .B(n_135), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_51), .A2(n_60), .B1(n_154), .B2(n_176), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_52), .A2(n_144), .B1(n_176), .B2(n_178), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_53), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_54), .B(n_154), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_55), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_56), .B(n_154), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_57), .A2(n_153), .B(n_165), .C(n_167), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_58), .Y(n_225) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_62), .A2(n_101), .B1(n_114), .B2(n_752), .C1(n_757), .C2(n_771), .Y(n_100) );
INVx1_ASAP7_75t_L g762 ( .A(n_62), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_63), .B(n_154), .Y(n_466) );
INVx1_ASAP7_75t_L g132 ( .A(n_64), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_65), .Y(n_106) );
AO32x2_ASAP7_75t_L g492 ( .A1(n_66), .A2(n_128), .A3(n_229), .B1(n_487), .B2(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g485 ( .A(n_67), .Y(n_485) );
INVx1_ASAP7_75t_L g520 ( .A(n_68), .Y(n_520) );
INVx1_ASAP7_75t_L g739 ( .A(n_69), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_SL g148 ( .A1(n_70), .A2(n_149), .B(n_150), .C(n_153), .Y(n_148) );
INVxp67_ASAP7_75t_L g151 ( .A(n_71), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_72), .B(n_176), .Y(n_521) );
INVx1_ASAP7_75t_L g105 ( .A(n_73), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_74), .Y(n_186) );
INVx1_ASAP7_75t_L g218 ( .A(n_75), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_77), .A2(n_140), .B(n_144), .C(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_78), .B(n_495), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_79), .B(n_176), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_80), .B(n_194), .Y(n_208) );
INVx2_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_82), .B(n_149), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_83), .B(n_176), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_84), .A2(n_140), .B(n_144), .C(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g109 ( .A(n_85), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g117 ( .A(n_85), .B(n_111), .Y(n_117) );
INVx2_ASAP7_75t_L g446 ( .A(n_85), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_87), .A2(n_99), .B1(n_176), .B2(n_177), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_88), .B(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_89), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_90), .A2(n_140), .B(n_144), .C(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_91), .Y(n_239) );
INVx1_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_93), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_94), .B(n_194), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_95), .B(n_176), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_96), .B(n_128), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_97), .B(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_98), .A2(n_135), .B(n_142), .Y(n_134) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_SL g756 ( .A(n_104), .Y(n_756) );
INVx1_ASAP7_75t_L g755 ( .A(n_106), .Y(n_755) );
OA21x2_ASAP7_75t_L g772 ( .A1(n_106), .A2(n_756), .B(n_769), .Y(n_772) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_109), .Y(n_767) );
BUFx2_ASAP7_75t_L g769 ( .A(n_109), .Y(n_769) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_110), .B(n_446), .Y(n_750) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g445 ( .A(n_111), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI222xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_738), .B1(n_741), .B2(n_746), .C1(n_747), .C2(n_751), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_118), .B1(n_444), .B2(n_447), .Y(n_115) );
INVx2_ASAP7_75t_L g743 ( .A(n_116), .Y(n_743) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_119), .A2(n_742), .B1(n_744), .B2(n_745), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_119), .A2(n_760), .B1(n_761), .B2(n_764), .Y(n_759) );
INVx2_ASAP7_75t_L g764 ( .A(n_119), .Y(n_764) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND4x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_362), .C(n_409), .D(n_429), .Y(n_120) );
NOR3xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_292), .C(n_317), .Y(n_121) );
OAI211xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_200), .B(n_252), .C(n_282), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_171), .Y(n_124) );
INVx3_ASAP7_75t_SL g334 ( .A(n_125), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_125), .B(n_265), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_125), .B(n_187), .Y(n_415) );
AND2x2_ASAP7_75t_L g438 ( .A(n_125), .B(n_304), .Y(n_438) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_159), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g256 ( .A(n_127), .B(n_160), .Y(n_256) );
INVx3_ASAP7_75t_L g269 ( .A(n_127), .Y(n_269) );
AND2x2_ASAP7_75t_L g274 ( .A(n_127), .B(n_159), .Y(n_274) );
OR2x2_ASAP7_75t_L g325 ( .A(n_127), .B(n_266), .Y(n_325) );
BUFx2_ASAP7_75t_L g345 ( .A(n_127), .Y(n_345) );
AND2x2_ASAP7_75t_L g355 ( .A(n_127), .B(n_266), .Y(n_355) );
AND2x2_ASAP7_75t_L g361 ( .A(n_127), .B(n_172), .Y(n_361) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B(n_156), .Y(n_127) );
INVx4_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_128), .A2(n_471), .B(n_478), .Y(n_470) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_130), .B(n_131), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx2_ASAP7_75t_L g243 ( .A(n_135), .Y(n_243) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_136), .B(n_140), .Y(n_184) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g464 ( .A(n_137), .Y(n_464) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx1_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
INVx1_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
INVx1_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
INVx4_ASAP7_75t_SL g155 ( .A(n_140), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_140), .A2(n_458), .B(n_462), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_140), .A2(n_472), .B(n_475), .Y(n_471) );
BUFx3_ASAP7_75t_L g487 ( .A(n_140), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_140), .A2(n_500), .B(n_504), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_140), .A2(n_519), .B(n_522), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_147), .B(n_148), .C(n_155), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_155), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_143), .A2(n_155), .B(n_245), .C(n_246), .Y(n_244) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_145), .Y(n_154) );
BUFx3_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
INVx1_ASAP7_75t_L g495 ( .A(n_145), .Y(n_495) );
INVx1_ASAP7_75t_L g503 ( .A(n_149), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_152), .B(n_168), .Y(n_167) );
INVx5_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_152), .A2(n_166), .B1(n_494), .B2(n_496), .Y(n_493) );
O2A1O1Ixp5_ASAP7_75t_SL g519 ( .A1(n_153), .A2(n_194), .B(n_520), .C(n_521), .Y(n_519) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_154), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_155), .A2(n_175), .B1(n_183), .B2(n_184), .Y(n_174) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_157), .A2(n_161), .B(n_169), .Y(n_160) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_158), .B(n_215), .Y(n_214) );
AO21x1_ASAP7_75t_L g531 ( .A1(n_158), .A2(n_532), .B(n_535), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_158), .B(n_487), .C(n_532), .Y(n_550) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_160), .B(n_266), .Y(n_280) );
INVx2_ASAP7_75t_L g290 ( .A(n_160), .Y(n_290) );
AND2x2_ASAP7_75t_L g303 ( .A(n_160), .B(n_269), .Y(n_303) );
OR2x2_ASAP7_75t_L g314 ( .A(n_160), .B(n_266), .Y(n_314) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_160), .B(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g372 ( .A(n_160), .Y(n_372) );
AND2x2_ASAP7_75t_L g418 ( .A(n_160), .B(n_172), .Y(n_418) );
O2A1O1Ixp5_ASAP7_75t_L g484 ( .A1(n_165), .A2(n_463), .B(n_485), .C(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_165), .A2(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g235 ( .A(n_166), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_166), .A2(n_467), .B1(n_510), .B2(n_511), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_166), .A2(n_467), .B1(n_533), .B2(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
INVx2_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_170), .A2(n_242), .B(n_251), .Y(n_241) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_170), .A2(n_499), .B(n_507), .Y(n_498) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_170), .A2(n_518), .B(n_525), .Y(n_517) );
INVx3_ASAP7_75t_SL g291 ( .A(n_171), .Y(n_291) );
OR2x2_ASAP7_75t_L g344 ( .A(n_171), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_187), .Y(n_171) );
INVx3_ASAP7_75t_L g266 ( .A(n_172), .Y(n_266) );
AND2x2_ASAP7_75t_L g333 ( .A(n_172), .B(n_188), .Y(n_333) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_172), .Y(n_401) );
AOI33xp33_ASAP7_75t_L g405 ( .A1(n_172), .A2(n_334), .A3(n_341), .B1(n_350), .B2(n_406), .B3(n_407), .Y(n_405) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_185), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_173), .B(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_173), .A2(n_189), .B(n_197), .Y(n_188) );
INVx2_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
INVx2_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_178) );
INVx2_ASAP7_75t_L g181 ( .A(n_179), .Y(n_181) );
INVx4_ASAP7_75t_L g247 ( .A(n_179), .Y(n_247) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_184), .A2(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_184), .A2(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_L g254 ( .A(n_187), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_187), .B(n_269), .Y(n_268) );
NOR3xp33_ASAP7_75t_L g328 ( .A(n_187), .B(n_329), .C(n_331), .Y(n_328) );
AND2x2_ASAP7_75t_L g354 ( .A(n_187), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_187), .B(n_361), .Y(n_364) );
AND2x2_ASAP7_75t_L g417 ( .A(n_187), .B(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
OR2x2_ASAP7_75t_L g367 ( .A(n_188), .B(n_266), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .C(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g467 ( .A(n_194), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_194), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_194), .A2(n_482), .B(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_196), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_199), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_199), .B(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_226), .Y(n_200) );
AOI32xp33_ASAP7_75t_L g318 ( .A1(n_201), .A2(n_319), .A3(n_321), .B1(n_323), .B2(n_326), .Y(n_318) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_201), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g421 ( .A(n_201), .Y(n_421) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g353 ( .A(n_202), .B(n_337), .Y(n_353) );
AND2x2_ASAP7_75t_L g373 ( .A(n_202), .B(n_299), .Y(n_373) );
AND2x2_ASAP7_75t_L g441 ( .A(n_202), .B(n_359), .Y(n_441) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_216), .Y(n_202) );
INVx3_ASAP7_75t_L g262 ( .A(n_203), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_203), .B(n_260), .Y(n_276) );
OR2x2_ASAP7_75t_L g281 ( .A(n_203), .B(n_259), .Y(n_281) );
INVx1_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_270), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_203), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_203), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g351 ( .A(n_203), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_203), .B(n_436), .Y(n_435) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B(n_213), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_210), .A2(n_221), .B(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g250 ( .A(n_212), .Y(n_250) );
INVx1_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_213), .A2(n_457), .B(n_468), .Y(n_456) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_213), .A2(n_480), .B(n_488), .Y(n_479) );
INVx2_ASAP7_75t_L g260 ( .A(n_216), .Y(n_260) );
AND2x2_ASAP7_75t_L g306 ( .A(n_216), .B(n_227), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_216), .B(n_241), .Y(n_316) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_223), .B(n_224), .Y(n_216) );
INVx2_ASAP7_75t_L g436 ( .A(n_226), .Y(n_436) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_240), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_227), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
AND2x2_ASAP7_75t_L g321 ( .A(n_227), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g337 ( .A(n_227), .B(n_300), .Y(n_337) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
AND2x2_ASAP7_75t_L g299 ( .A(n_228), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g350 ( .A(n_228), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_228), .B(n_260), .Y(n_382) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_238), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_236), .Y(n_232) );
AND2x2_ASAP7_75t_L g261 ( .A(n_240), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g322 ( .A(n_240), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_240), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g359 ( .A(n_240), .Y(n_359) );
INVx1_ASAP7_75t_L g392 ( .A(n_240), .Y(n_392) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g270 ( .A(n_241), .B(n_260), .Y(n_270) );
INVx1_ASAP7_75t_L g300 ( .A(n_241), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_247), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g461 ( .A(n_247), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_247), .A2(n_523), .B(n_524), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B1(n_263), .B2(n_270), .C(n_271), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_254), .B(n_274), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_254), .B(n_337), .Y(n_414) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_256), .B(n_304), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_256), .B(n_265), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_256), .B(n_279), .Y(n_408) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
AND2x2_ASAP7_75t_L g305 ( .A(n_261), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g383 ( .A(n_261), .Y(n_383) );
AND2x2_ASAP7_75t_L g315 ( .A(n_262), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_262), .B(n_285), .Y(n_331) );
AND2x2_ASAP7_75t_L g395 ( .A(n_262), .B(n_321), .Y(n_395) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g304 ( .A(n_266), .B(n_273), .Y(n_304) );
AND2x2_ASAP7_75t_L g400 ( .A(n_267), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_269), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_270), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_270), .B(n_277), .Y(n_365) );
AND2x2_ASAP7_75t_L g385 ( .A(n_270), .B(n_285), .Y(n_385) );
AND2x2_ASAP7_75t_L g406 ( .A(n_270), .B(n_350), .Y(n_406) );
OAI32xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_275), .A3(n_277), .B1(n_278), .B2(n_281), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_SL g279 ( .A(n_273), .Y(n_279) );
NAND2x1_ASAP7_75t_L g320 ( .A(n_273), .B(n_303), .Y(n_320) );
OR2x2_ASAP7_75t_L g324 ( .A(n_273), .B(n_325), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_273), .B(n_372), .Y(n_425) );
INVx1_ASAP7_75t_L g293 ( .A(n_274), .Y(n_293) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_275), .A2(n_366), .B1(n_412), .B2(n_415), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g283 ( .A(n_276), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g326 ( .A(n_276), .B(n_299), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_276), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g404 ( .A(n_276), .B(n_337), .Y(n_404) );
INVxp67_ASAP7_75t_L g340 ( .A(n_277), .Y(n_340) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g410 ( .A(n_279), .B(n_397), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_279), .B(n_360), .Y(n_433) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_281), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g426 ( .A(n_281), .B(n_427), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_286), .B(n_289), .Y(n_282) );
AND2x2_ASAP7_75t_L g295 ( .A(n_284), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g379 ( .A(n_288), .B(n_299), .Y(n_379) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g397 ( .A(n_290), .B(n_355), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_290), .B(n_354), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_291), .B(n_303), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_297), .C(n_307), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_293), .A2(n_328), .B1(n_332), .B2(n_335), .C(n_338), .Y(n_327) );
AOI31xp33_ASAP7_75t_L g422 ( .A1(n_293), .A2(n_423), .A3(n_424), .B(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_303), .B2(n_305), .Y(n_297) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g423 ( .A(n_303), .Y(n_423) );
INVx1_ASAP7_75t_L g386 ( .A(n_304), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g429 ( .A1(n_306), .A2(n_430), .B(n_432), .C(n_434), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B1(n_311), .B2(n_315), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_312), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_314), .A2(n_348), .B1(n_367), .B2(n_403), .C(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g398 ( .A(n_315), .Y(n_398) );
INVx1_ASAP7_75t_L g352 ( .A(n_316), .Y(n_352) );
NAND3xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_327), .C(n_342), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_319), .A2(n_369), .B(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_321), .B(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g428 ( .A(n_322), .Y(n_428) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_349), .Y(n_366) );
INVx1_ASAP7_75t_L g341 ( .A(n_330), .Y(n_341) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g339 ( .A(n_333), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_333), .B(n_371), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g338 ( .A(n_334), .B(n_339), .C(n_340), .D(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .B1(n_353), .B2(n_354), .C1(n_356), .C2(n_360), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g440 ( .A(n_344), .Y(n_440) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_356), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_SL g416 ( .A1(n_361), .A2(n_417), .B(n_419), .Y(n_416) );
NOR4xp25_ASAP7_75t_L g362 ( .A(n_363), .B(n_374), .C(n_387), .D(n_402), .Y(n_362) );
OAI221xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_365), .B1(n_366), .B2(n_367), .C(n_368), .Y(n_363) );
INVx1_ASAP7_75t_L g443 ( .A(n_364), .Y(n_443) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_371), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OAI222xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_380), .B2(n_381), .C1(n_384), .C2(n_386), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI211xp5_ASAP7_75t_L g409 ( .A1(n_379), .A2(n_410), .B(n_411), .C(n_422), .Y(n_409) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OAI222xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .B1(n_394), .B2(n_396), .C1(n_398), .C2(n_399), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_404), .A2(n_407), .B1(n_440), .B2(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_437), .B(n_439), .C(n_442), .Y(n_434) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx6_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g744 ( .A(n_445), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_447), .Y(n_745) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_448), .B(n_704), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_608), .C(n_692), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_551), .C(n_573), .D(n_589), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_489), .B1(n_512), .B2(n_530), .C(n_537), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_469), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_453), .B(n_530), .Y(n_563) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_453), .B(n_591), .C(n_604), .D(n_606), .Y(n_603) );
INVxp67_ASAP7_75t_L g720 ( .A(n_453), .Y(n_720) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g602 ( .A(n_454), .B(n_540), .Y(n_602) );
AND2x2_ASAP7_75t_L g626 ( .A(n_454), .B(n_469), .Y(n_626) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g593 ( .A(n_455), .B(n_529), .Y(n_593) );
AND2x2_ASAP7_75t_L g633 ( .A(n_455), .B(n_614), .Y(n_633) );
AND2x2_ASAP7_75t_L g650 ( .A(n_455), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_455), .B(n_470), .Y(n_674) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g528 ( .A(n_456), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g545 ( .A(n_456), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g557 ( .A(n_456), .B(n_470), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_456), .B(n_479), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B(n_466), .C(n_467), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_467), .A2(n_476), .B(n_477), .Y(n_475) );
AND2x2_ASAP7_75t_L g560 ( .A(n_469), .B(n_561), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_469), .A2(n_610), .B1(n_613), .B2(n_615), .C(n_619), .Y(n_609) );
AND2x2_ASAP7_75t_L g668 ( .A(n_469), .B(n_633), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_469), .B(n_650), .Y(n_702) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
INVx3_ASAP7_75t_L g529 ( .A(n_470), .Y(n_529) );
AND2x2_ASAP7_75t_L g577 ( .A(n_470), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g631 ( .A(n_470), .B(n_546), .Y(n_631) );
AND2x2_ASAP7_75t_L g689 ( .A(n_470), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g530 ( .A(n_479), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g546 ( .A(n_479), .Y(n_546) );
INVx1_ASAP7_75t_L g601 ( .A(n_479), .Y(n_601) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_479), .Y(n_607) );
AND2x2_ASAP7_75t_L g652 ( .A(n_479), .B(n_529), .Y(n_652) );
OR2x2_ASAP7_75t_L g691 ( .A(n_479), .B(n_531), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_484), .B(n_487), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_489), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_497), .Y(n_489) );
AND2x2_ASAP7_75t_L g687 ( .A(n_490), .B(n_684), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_490), .B(n_669), .Y(n_719) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g618 ( .A(n_491), .B(n_542), .Y(n_618) );
AND2x2_ASAP7_75t_L g667 ( .A(n_491), .B(n_515), .Y(n_667) );
INVx1_ASAP7_75t_L g713 ( .A(n_491), .Y(n_713) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_492), .Y(n_527) );
AND2x2_ASAP7_75t_L g568 ( .A(n_492), .B(n_542), .Y(n_568) );
INVx1_ASAP7_75t_L g585 ( .A(n_492), .Y(n_585) );
AND2x2_ASAP7_75t_L g591 ( .A(n_492), .B(n_508), .Y(n_591) );
AND2x2_ASAP7_75t_L g659 ( .A(n_497), .B(n_567), .Y(n_659) );
INVx2_ASAP7_75t_L g724 ( .A(n_497), .Y(n_724) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
AND2x2_ASAP7_75t_L g541 ( .A(n_498), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g554 ( .A(n_498), .B(n_516), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_498), .B(n_515), .Y(n_582) );
INVx1_ASAP7_75t_L g588 ( .A(n_498), .Y(n_588) );
INVx1_ASAP7_75t_L g605 ( .A(n_498), .Y(n_605) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_498), .Y(n_617) );
INVx2_ASAP7_75t_L g685 ( .A(n_498), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_503), .Y(n_500) );
INVx2_ASAP7_75t_L g542 ( .A(n_508), .Y(n_542) );
BUFx2_ASAP7_75t_L g639 ( .A(n_508), .Y(n_639) );
AND2x2_ASAP7_75t_L g684 ( .A(n_508), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_526), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_514), .B(n_621), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_514), .A2(n_683), .B(n_697), .Y(n_707) );
AND2x2_ASAP7_75t_L g732 ( .A(n_514), .B(n_618), .Y(n_732) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g654 ( .A(n_516), .Y(n_654) );
AND2x2_ASAP7_75t_L g683 ( .A(n_516), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_517), .Y(n_567) );
INVx2_ASAP7_75t_L g586 ( .A(n_517), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_517), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g540 ( .A(n_527), .Y(n_540) );
OR2x2_ASAP7_75t_L g553 ( .A(n_527), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g621 ( .A(n_527), .B(n_617), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_527), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g722 ( .A(n_527), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_527), .B(n_659), .Y(n_734) );
AND2x2_ASAP7_75t_L g613 ( .A(n_528), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g636 ( .A(n_528), .B(n_530), .Y(n_636) );
INVx2_ASAP7_75t_L g548 ( .A(n_529), .Y(n_548) );
AND2x2_ASAP7_75t_L g576 ( .A(n_529), .B(n_549), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_529), .B(n_601), .Y(n_657) );
AND2x2_ASAP7_75t_L g571 ( .A(n_530), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g718 ( .A(n_530), .Y(n_718) );
AND2x2_ASAP7_75t_L g730 ( .A(n_530), .B(n_593), .Y(n_730) );
AND2x2_ASAP7_75t_L g556 ( .A(n_531), .B(n_546), .Y(n_556) );
INVx1_ASAP7_75t_L g651 ( .A(n_531), .Y(n_651) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g549 ( .A(n_536), .B(n_550), .Y(n_549) );
INVxp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_540), .B(n_587), .Y(n_596) );
OR2x2_ASAP7_75t_L g728 ( .A(n_540), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g645 ( .A(n_541), .B(n_586), .Y(n_645) );
AND2x2_ASAP7_75t_L g653 ( .A(n_541), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g712 ( .A(n_541), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g736 ( .A(n_541), .B(n_583), .Y(n_736) );
NOR2xp67_ASAP7_75t_L g694 ( .A(n_542), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g723 ( .A(n_542), .B(n_586), .Y(n_723) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
AND2x2_ASAP7_75t_L g575 ( .A(n_545), .B(n_576), .Y(n_575) );
INVxp67_ASAP7_75t_L g737 ( .A(n_545), .Y(n_737) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g572 ( .A(n_548), .Y(n_572) );
AND2x2_ASAP7_75t_L g623 ( .A(n_548), .B(n_556), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_548), .B(n_691), .Y(n_717) );
INVx2_ASAP7_75t_L g562 ( .A(n_549), .Y(n_562) );
INVx3_ASAP7_75t_L g614 ( .A(n_549), .Y(n_614) );
OR2x2_ASAP7_75t_L g642 ( .A(n_549), .B(n_643), .Y(n_642) );
AOI311xp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .A3(n_557), .B(n_558), .C(n_569), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_552), .A2(n_590), .B(n_592), .C(n_594), .Y(n_589) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g574 ( .A(n_554), .Y(n_574) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g592 ( .A(n_556), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_556), .B(n_572), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_556), .B(n_557), .Y(n_725) );
AND2x2_ASAP7_75t_L g647 ( .A(n_557), .B(n_561), .Y(n_647) );
AOI21xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_563), .B(n_564), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g705 ( .A(n_561), .B(n_593), .Y(n_705) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_562), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g599 ( .A(n_562), .Y(n_599) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
AND2x2_ASAP7_75t_L g590 ( .A(n_566), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g635 ( .A(n_568), .Y(n_635) );
AND2x4_ASAP7_75t_L g697 ( .A(n_568), .B(n_666), .Y(n_697) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g648 ( .A1(n_571), .A2(n_637), .B1(n_649), .B2(n_653), .C1(n_655), .C2(n_659), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B(n_577), .C(n_580), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_574), .B(n_618), .Y(n_641) );
INVx1_ASAP7_75t_L g663 ( .A(n_576), .Y(n_663) );
INVx1_ASAP7_75t_L g597 ( .A(n_578), .Y(n_597) );
OR2x2_ASAP7_75t_L g662 ( .A(n_579), .B(n_663), .Y(n_662) );
OAI21xp33_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_583), .B(n_587), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_581), .B(n_599), .C(n_600), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_581), .A2(n_618), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_585), .Y(n_638) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_586), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g695 ( .A(n_586), .Y(n_695) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_586), .Y(n_711) );
INVx2_ASAP7_75t_L g669 ( .A(n_587), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_591), .B(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g643 ( .A(n_593), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B1(n_598), .B2(n_602), .C(n_603), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_597), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g731 ( .A(n_597), .Y(n_731) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g612 ( .A(n_604), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_604), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g670 ( .A(n_604), .B(n_618), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_604), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g703 ( .A(n_604), .B(n_638), .Y(n_703) );
BUFx3_ASAP7_75t_L g666 ( .A(n_605), .Y(n_666) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND5xp2_ASAP7_75t_L g608 ( .A(n_609), .B(n_627), .C(n_648), .D(n_660), .E(n_675), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI32xp33_ASAP7_75t_L g700 ( .A1(n_612), .A2(n_639), .A3(n_655), .B1(n_701), .B2(n_703), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_614), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g624 ( .A(n_618), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B1(n_624), .B2(n_625), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_634), .B1(n_636), .B2(n_637), .C(n_640), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g699 ( .A(n_631), .B(n_650), .Y(n_699) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_636), .A2(n_697), .B1(n_715), .B2(n_720), .C(n_721), .Y(n_714) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx2_ASAP7_75t_L g680 ( .A(n_639), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_644), .B2(n_646), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g658 ( .A(n_650), .Y(n_658) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AOI222xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B1(n_668), .B2(n_669), .C1(n_670), .C2(n_671), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_669), .A2(n_716), .B1(n_718), .B2(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_686), .B(n_688), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g729 ( .A(n_684), .Y(n_729) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_696), .B(n_698), .C(n_700), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B(n_708), .C(n_733), .Y(n_704) );
CKINVDCx16_ASAP7_75t_R g709 ( .A(n_705), .Y(n_709) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI211xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B(n_714), .C(n_726), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B(n_725), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g746 ( .A(n_738), .Y(n_746) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVxp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_765), .B(n_768), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_SL g768 ( .A(n_769), .B(n_770), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
endmodule