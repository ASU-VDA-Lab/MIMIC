module fake_jpeg_23174_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_23),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_1),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_20),
.B(n_17),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_14),
.B1(n_19),
.B2(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_13),
.B1(n_21),
.B2(n_18),
.Y(n_53)
);

OA21x2_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_16),
.B(n_19),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_26),
.B1(n_13),
.B2(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_15),
.B1(n_27),
.B2(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_46),
.Y(n_68)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_28),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_62),
.C(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_64),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_50),
.Y(n_71)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx12f_ASAP7_75t_SL g83 ( 
.A(n_66),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_44),
.B(n_39),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_55),
.B(n_62),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_77),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_75),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_43),
.C(n_31),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_76),
.C(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_37),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_87),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_88),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_72),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_47),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_99),
.Y(n_107)
);

AOI22x1_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_66),
.B1(n_76),
.B2(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_90),
.B1(n_83),
.B2(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_6),
.A3(n_9),
.B1(n_12),
.B2(n_20),
.C1(n_3),
.C2(n_4),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_87),
.C(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_108),
.C(n_95),
.Y(n_111)
);

AO221x1_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_70),
.B1(n_60),
.B2(n_64),
.C(n_47),
.Y(n_105)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_98),
.C(n_96),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_31),
.C(n_33),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_115),
.B(n_116),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_99),
.B1(n_84),
.B2(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_106),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_85),
.A3(n_86),
.B1(n_88),
.B2(n_33),
.C(n_32),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_2),
.B(n_3),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_121),
.B(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_32),
.B1(n_23),
.B2(n_20),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_104),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_116),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_124),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_2),
.B(n_32),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_17),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_125),
.Y(n_129)
);


endmodule