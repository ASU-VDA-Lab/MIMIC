module fake_jpeg_17482_n_386 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_40),
.B(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g80 ( 
.A(n_47),
.Y(n_80)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_61),
.Y(n_93)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_66),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_19),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_68),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_14),
.B(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_3),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_70),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_38),
.B1(n_26),
.B2(n_24),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_83),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_38),
.B1(n_24),
.B2(n_26),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_73),
.B(n_90),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_23),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_89),
.C(n_5),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_18),
.B1(n_26),
.B2(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_18),
.B1(n_37),
.B2(n_19),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_15),
.C(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_29),
.Y(n_90)
);

AND2x4_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_36),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_109),
.B(n_5),
.C(n_6),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_43),
.B(n_17),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_98),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_47),
.B(n_17),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_39),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_101),
.A2(n_111),
.B1(n_112),
.B2(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_35),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_42),
.B(n_34),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_44),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_113),
.B(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_49),
.B(n_27),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_53),
.A2(n_22),
.B1(n_34),
.B2(n_36),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_46),
.B(n_22),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_48),
.A2(n_20),
.B1(n_36),
.B2(n_34),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_140),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_3),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_126),
.A2(n_131),
.B(n_139),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_36),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_154),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_133),
.A2(n_172),
.B1(n_75),
.B2(n_82),
.Y(n_207)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_4),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_93),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_146),
.Y(n_182)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_156),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_5),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_80),
.B(n_91),
.Y(n_197)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_12),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_108),
.Y(n_185)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_7),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_7),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_7),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_164),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_74),
.B(n_8),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_166),
.C(n_170),
.Y(n_187)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g186 ( 
.A(n_159),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_77),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g162 ( 
.A1(n_71),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_112),
.B1(n_111),
.B2(n_170),
.Y(n_177)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_9),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_114),
.B(n_12),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g168 ( 
.A(n_80),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_169),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_76),
.B(n_9),
.C(n_10),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_81),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_188),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_177),
.B(n_191),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_161),
.A2(n_81),
.B1(n_122),
.B2(n_87),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_99),
.B1(n_108),
.B2(n_117),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_163),
.B1(n_169),
.B2(n_148),
.Y(n_228)
);

NOR2x1_ASAP7_75t_R g250 ( 
.A(n_185),
.B(n_197),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_153),
.B(n_78),
.Y(n_191)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_91),
.C(n_102),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_212),
.C(n_128),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_121),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_102),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_132),
.B(n_107),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_208),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_139),
.B1(n_166),
.B2(n_147),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_107),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_152),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_129),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_75),
.C(n_155),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_143),
.B(n_131),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_194),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_124),
.A2(n_149),
.B1(n_134),
.B2(n_167),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_166),
.B1(n_147),
.B2(n_127),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_149),
.A2(n_125),
.A3(n_126),
.B1(n_162),
.B2(n_131),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_139),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_149),
.B(n_126),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_218),
.A2(n_220),
.B1(n_231),
.B2(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_136),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_222),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_138),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_229),
.Y(n_262)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_227),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_232),
.B1(n_247),
.B2(n_255),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_138),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_230),
.B(n_233),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_158),
.B(n_142),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_162),
.B1(n_144),
.B2(n_150),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_130),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_238),
.C(n_242),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_130),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_253),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_153),
.C(n_159),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_168),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_239),
.Y(n_275)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_142),
.Y(n_240)
);

AOI21x1_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_186),
.B(n_174),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_SL g246 ( 
.A1(n_182),
.A2(n_185),
.B(n_187),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_248),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_208),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_200),
.C(n_187),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_193),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_182),
.A2(n_213),
.B1(n_177),
.B2(n_179),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_209),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_188),
.A2(n_183),
.B(n_176),
.C(n_210),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_254),
.A2(n_175),
.B1(n_174),
.B2(n_195),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_179),
.A2(n_197),
.B1(n_193),
.B2(n_186),
.Y(n_255)
);

INVx4_ASAP7_75t_SL g256 ( 
.A(n_240),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_256),
.A2(n_209),
.B1(n_205),
.B2(n_195),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_259),
.B(n_266),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_278),
.B(n_239),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_264),
.B(n_270),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_180),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_252),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_272),
.B(n_284),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_219),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_274),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_224),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_225),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_245),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_230),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_255),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_204),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_227),
.C(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_263),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_300),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_256),
.A2(n_240),
.B1(n_250),
.B2(n_217),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_290),
.A2(n_292),
.B1(n_309),
.B2(n_276),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_260),
.A2(n_250),
.B1(n_217),
.B2(n_235),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_293),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_232),
.B1(n_247),
.B2(n_228),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_294),
.A2(n_301),
.B1(n_306),
.B2(n_308),
.Y(n_317)
);

AOI22x1_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_254),
.B1(n_239),
.B2(n_231),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_295),
.A2(n_258),
.B1(n_257),
.B2(n_262),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_312),
.C(n_267),
.Y(n_318)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_297),
.Y(n_323)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_299),
.Y(n_331)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_247),
.B1(n_234),
.B2(n_251),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_302),
.A2(n_282),
.B(n_277),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_251),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_305),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_283),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_220),
.B1(n_218),
.B2(n_238),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_241),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_293),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_268),
.A2(n_234),
.B1(n_287),
.B2(n_277),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_311),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_270),
.B(n_226),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_268),
.A2(n_238),
.B1(n_190),
.B2(n_199),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_294),
.B1(n_312),
.B2(n_272),
.Y(n_320)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_267),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_318),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_291),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_320),
.A2(n_295),
.B1(n_292),
.B2(n_298),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_261),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_309),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_276),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_330),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_326),
.B(n_334),
.Y(n_346)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_301),
.B(n_261),
.CI(n_284),
.CON(n_327),
.SN(n_327)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_327),
.B(n_295),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_285),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_264),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_290),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_335),
.A2(n_289),
.B(n_314),
.C(n_300),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_334),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_340),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_302),
.B(n_288),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_342),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_343),
.A2(n_325),
.B1(n_323),
.B2(n_328),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_258),
.Y(n_344)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_314),
.Y(n_345)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_321),
.B(n_199),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_348),
.C(n_318),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_181),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_181),
.Y(n_351)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_335),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_352),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_349),
.Y(n_366)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_350),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_359),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_356),
.B(n_339),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_343),
.A2(n_328),
.B1(n_315),
.B2(n_317),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_357),
.A2(n_343),
.B1(n_346),
.B2(n_327),
.Y(n_369)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_336),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_365),
.B(n_369),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_349),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_363),
.A2(n_343),
.B1(n_346),
.B2(n_327),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_368),
.A2(n_371),
.B1(n_370),
.B2(n_369),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_347),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_370),
.A2(n_354),
.B(n_358),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_373),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_358),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_376),
.B(n_359),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_374),
.A2(n_361),
.B1(n_364),
.B2(n_355),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_356),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_379),
.B(n_380),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_L g382 ( 
.A1(n_381),
.A2(n_367),
.B(n_362),
.Y(n_382)
);

OAI321xp33_ASAP7_75t_L g383 ( 
.A1(n_382),
.A2(n_357),
.A3(n_371),
.B1(n_378),
.B2(n_353),
.C(n_366),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_378),
.B(n_322),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g385 ( 
.A(n_384),
.B(n_339),
.CI(n_319),
.CON(n_385),
.SN(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_316),
.Y(n_386)
);


endmodule