module real_jpeg_7915_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_327, n_1, n_328, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_327;
input n_1;
input n_328;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_63),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_3),
.A2(n_32),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_32),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_3),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_28),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_3),
.B(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_54),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_29),
.B(n_49),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_127),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_4),
.A2(n_38),
.B1(n_69),
.B2(n_70),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_10),
.A2(n_69),
.B1(n_70),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_10),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_107),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_107),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_107),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_11),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_143),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_143),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_143),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_12),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_69),
.B1(n_70),
.B2(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_114),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_13),
.A2(n_53),
.B1(n_69),
.B2(n_70),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_45),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_14),
.A2(n_45),
.B1(n_69),
.B2(n_70),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_16),
.A2(n_69),
.B1(n_70),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_16),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_102),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_102),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_102),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_17),
.A2(n_43),
.B1(n_44),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_17),
.A2(n_69),
.B1(n_70),
.B2(n_82),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_82),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_17),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_88),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_74),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_55),
.B1(n_56),
.B2(n_73),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_22),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_35),
.B(n_36),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_25),
.A2(n_35),
.B1(n_87),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_26),
.A2(n_31),
.B1(n_37),
.B2(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_26),
.A2(n_31),
.B1(n_59),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_26),
.A2(n_31),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_26),
.A2(n_31),
.B1(n_153),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_26),
.A2(n_31),
.B1(n_169),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_26),
.A2(n_31),
.B1(n_209),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_26),
.A2(n_31),
.B1(n_220),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_26),
.A2(n_31),
.B1(n_246),
.B2(n_264),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_51)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_30),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_31),
.B(n_127),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_32),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_32),
.B(n_34),
.Y(n_157)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_33),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_47),
.B1(n_51),
.B2(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_48),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_44),
.A2(n_48),
.B(n_127),
.C(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_46),
.A2(n_54),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_51),
.B1(n_62),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_47),
.A2(n_51),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_47),
.A2(n_51),
.B1(n_224),
.B2(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_47),
.A2(n_51),
.B1(n_249),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_47),
.A2(n_51),
.B1(n_81),
.B2(n_267),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.C(n_64),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_58),
.B1(n_64),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_61),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_64),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_68),
.B(n_72),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_68),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_65),
.A2(n_68),
.B1(n_113),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_65),
.A2(n_68),
.B1(n_140),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_65),
.A2(n_68),
.B1(n_149),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_65),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_65),
.A2(n_68),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_65),
.A2(n_68),
.B1(n_232),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_65),
.A2(n_68),
.B1(n_241),
.B2(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_68),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_68),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_69),
.B(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_69),
.B(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_72),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.C(n_83),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_312),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.C(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_80),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_80),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_83),
.B(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI321xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_309),
.A3(n_319),
.B1(n_324),
.B2(n_325),
.C(n_327),
.Y(n_90)
);

AOI321xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_257),
.A3(n_297),
.B1(n_303),
.B2(n_308),
.C(n_328),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_214),
.C(n_253),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_184),
.B(n_213),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_163),
.B(n_183),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_145),
.B(n_162),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_134),
.B(n_144),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_120),
.B(n_133),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_108),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_103),
.A2(n_104),
.B1(n_161),
.B2(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_124),
.B1(n_125),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_115),
.B2(n_119),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_119),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_115),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_128),
.B(n_132),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_126),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_125),
.B1(n_142),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_124),
.A2(n_125),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_124),
.A2(n_125),
.B1(n_195),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_124),
.A2(n_125),
.B1(n_229),
.B2(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_124),
.A2(n_125),
.B(n_239),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_136),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_139),
.C(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_147),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.CI(n_154),
.CON(n_147),
.SN(n_147)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_159),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_165),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_176),
.B2(n_177),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_179),
.C(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_175),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_168),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_173),
.C(n_175),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_186),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_199),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_198),
.C(n_199),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_193),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_207),
.B2(n_208),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_207),
.C(n_210),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_204),
.A2(n_206),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_205),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_215),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_234),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_216),
.B(n_234),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.C(n_233),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_225),
.C(n_226),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_233),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_230),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_251),
.B2(n_252),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_242),
.C(n_252),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_240),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_247),
.C(n_250),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_255),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_276),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_258),
.B(n_276),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_269),
.C(n_275),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_260),
.B1(n_269),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_265),
.C(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_263),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_264),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_269),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_271),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_291),
.B(n_293),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_272),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_272),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_295),
.B2(n_296),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_287),
.B2(n_288),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_288),
.C(n_296),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_284),
.B(n_286),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_284),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_286),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_286),
.A2(n_311),
.B1(n_315),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_294),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_304),
.B(n_307),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_317),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_317),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.C(n_316),
.Y(n_310)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);


endmodule