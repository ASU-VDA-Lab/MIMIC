module real_jpeg_16815_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_572;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_581),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_0),
.B(n_582),
.Y(n_581)
);

AOI22x1_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_102),
.B1(n_184),
.B2(n_188),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_1),
.A2(n_45),
.B1(n_102),
.B2(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_102),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_2),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_2),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

OAI22x1_ASAP7_75t_SL g141 ( 
.A1(n_3),
.A2(n_54),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_3),
.A2(n_54),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_3),
.A2(n_54),
.B1(n_261),
.B2(n_264),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_4),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_5),
.A2(n_56),
.B1(n_223),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_5),
.A2(n_296),
.B1(n_393),
.B2(n_395),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_5),
.A2(n_296),
.B1(n_449),
.B2(n_453),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_5),
.A2(n_296),
.B1(n_496),
.B2(n_498),
.Y(n_495)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_6),
.A2(n_312),
.A3(n_314),
.B1(n_317),
.B2(n_321),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_6),
.A2(n_220),
.B1(n_320),
.B2(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_6),
.B(n_27),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_6),
.B(n_121),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_6),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_6),
.B(n_67),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_6),
.A2(n_320),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

OAI32xp33_ASAP7_75t_L g533 ( 
.A1(n_6),
.A2(n_534),
.A3(n_539),
.B1(n_540),
.B2(n_543),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_7),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_7),
.A2(n_279),
.B1(n_304),
.B2(n_307),
.Y(n_303)
);

OAI22x1_ASAP7_75t_L g457 ( 
.A1(n_7),
.A2(n_279),
.B1(n_458),
.B2(n_462),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_7),
.A2(n_279),
.B1(n_519),
.B2(n_522),
.Y(n_518)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_8),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_8),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_8),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_9),
.A2(n_45),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_9),
.A2(n_300),
.B1(n_357),
.B2(n_361),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_9),
.A2(n_300),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_9),
.A2(n_300),
.B1(n_477),
.B2(n_480),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g582 ( 
.A(n_10),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_11),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_11),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_11),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_11),
.Y(n_452)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_13),
.A2(n_39),
.B1(n_44),
.B2(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_13),
.A2(n_47),
.B1(n_164),
.B2(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_13),
.A2(n_47),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_13),
.A2(n_47),
.B1(n_329),
.B2(n_335),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_15),
.A2(n_110),
.B1(n_115),
.B2(n_116),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_15),
.A2(n_115),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_15),
.A2(n_115),
.B1(n_217),
.B2(n_222),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_15),
.A2(n_115),
.B1(n_344),
.B2(n_348),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_16),
.Y(n_334)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_240),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_238),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_212),
.Y(n_21)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_22),
.B(n_212),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_149),
.C(n_171),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_24),
.A2(n_149),
.B1(n_150),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_24),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_65),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_25),
.B(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_25),
.B(n_66),
.C(n_108),
.Y(n_237)
);

OAI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_38),
.B(n_48),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_26),
.A2(n_38),
.B1(n_59),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_26),
.A2(n_59),
.B1(n_295),
.B2(n_353),
.Y(n_352)
);

OAI22x1_ASAP7_75t_SL g381 ( 
.A1(n_26),
.A2(n_59),
.B1(n_276),
.B2(n_298),
.Y(n_381)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_27),
.B(n_49),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_27),
.B(n_207),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_27),
.A2(n_58),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_29),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_30),
.Y(n_144)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_30),
.Y(n_167)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_35),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_35),
.Y(n_538)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_42),
.Y(n_210)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_42),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_60)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_53),
.Y(n_224)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_57),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_57),
.Y(n_323)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_59),
.A2(n_206),
.B(n_211),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_59),
.A2(n_276),
.B(n_281),
.Y(n_275)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_62),
.Y(n_354)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_63),
.Y(n_278)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_64),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_108),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_66),
.A2(n_226),
.B1(n_227),
.B2(n_236),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_66),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_82),
.B(n_96),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_67),
.B(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_67),
.B(n_268),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_67),
.A2(n_82),
.B1(n_444),
.B2(n_448),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_67),
.A2(n_82),
.B1(n_448),
.B2(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_68),
.B(n_97),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_68),
.A2(n_194),
.B1(n_202),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_68),
.A2(n_202),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_76),
.B2(n_78),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_70),
.Y(n_336)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_70),
.Y(n_461)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_76),
.Y(n_349)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_77),
.Y(n_265)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_77),
.Y(n_484)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_77),
.Y(n_497)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_82),
.B(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_82),
.A2(n_160),
.B(n_561),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_86),
.Y(n_454)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_90),
.Y(n_441)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_94),
.Y(n_539)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_97),
.A2(n_202),
.B(n_203),
.Y(n_351)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_100),
.Y(n_468)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_106),
.Y(n_271)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_107),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_119),
.B(n_139),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_109),
.A2(n_119),
.B1(n_121),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_114),
.Y(n_363)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_118),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_119),
.B(n_141),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_119),
.A2(n_229),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_120),
.A2(n_163),
.B1(n_230),
.B2(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_120),
.A2(n_230),
.B1(n_303),
.B2(n_356),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_120),
.A2(n_140),
.B(n_231),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_120),
.A2(n_230),
.B1(n_356),
.B2(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_120),
.A2(n_230),
.B1(n_392),
.B2(n_527),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_129),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_123),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_125),
.Y(n_470)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_137),
.Y(n_129)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_141),
.Y(n_283)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_144),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_144),
.Y(n_547)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

INVxp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_150),
.A2(n_151),
.B(n_161),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_161),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_160),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_153),
.B(n_372),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_156),
.Y(n_521)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_166),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_166),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_171),
.A2(n_172),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_191),
.B(n_204),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_173),
.A2(n_174),
.B1(n_204),
.B2(n_205),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_173),
.A2(n_174),
.B1(n_193),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2x1_ASAP7_75t_R g192 ( 
.A(n_174),
.B(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_178),
.B(n_183),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_177),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_178),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_178),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_178),
.A2(n_457),
.B(n_464),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_178),
.A2(n_320),
.B1(n_492),
.B2(n_495),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_178),
.A2(n_476),
.B1(n_495),
.B2(n_507),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g494 ( 
.A(n_182),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_183),
.Y(n_552)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_187),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_190),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_193),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_202),
.B(n_203),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g427 ( 
.A1(n_195),
.A2(n_428),
.A3(n_432),
.B1(n_437),
.B2(n_439),
.Y(n_427)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_237),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_225),
.Y(n_214)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_235),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_232),
.Y(n_531)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_284),
.B(n_580),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_242),
.B(n_246),
.Y(n_580)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_252),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_248),
.A2(n_250),
.B1(n_251),
.B2(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_248),
.Y(n_420)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_252),
.B(n_419),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_275),
.C(n_282),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g411 ( 
.A(n_253),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_266),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_254),
.B(n_266),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_255),
.Y(n_464)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_258),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_259),
.A2(n_328),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_260),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_274),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_275),
.B(n_282),
.Y(n_412)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_574),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_421),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_404),
.C(n_416),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_384),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_373),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_290),
.B(n_373),
.C(n_576),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_350),
.C(n_364),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_291),
.B(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_310),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_293),
.B(n_301),
.C(n_310),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_326),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_311),
.B(n_326),
.Y(n_389)
);

INVx8_ASAP7_75t_L g528 ( 
.A(n_312),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_320),
.B(n_438),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_SL g444 ( 
.A1(n_320),
.A2(n_437),
.B(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_320),
.B(n_541),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_337),
.B2(n_343),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_343),
.B(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_327),
.A2(n_475),
.B1(n_485),
.B2(n_486),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_327),
.A2(n_366),
.B(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_333),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_336),
.Y(n_504)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_347),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_364),
.Y(n_403)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.C(n_355),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_355),
.Y(n_387)
);

XOR2x2_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_371),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_371),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_368),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_SL g486 ( 
.A(n_369),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_377),
.C(n_383),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_383),
.Y(n_375)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_376),
.Y(n_383)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_381),
.C(n_382),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_402),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_385),
.B(n_402),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.C(n_390),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_386),
.B(n_571),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_390),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_396),
.C(n_398),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_391),
.B(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_396),
.A2(n_397),
.B1(n_399),
.B2(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_399),
.Y(n_565)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g574 ( 
.A1(n_405),
.A2(n_575),
.B(n_577),
.C(n_578),
.D(n_579),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_406),
.B(n_407),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_413),
.B1(n_414),
.B2(n_415),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_408),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_411),
.C(n_413),
.Y(n_417)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_416),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_417),
.B(n_418),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_568),
.B(n_573),
.Y(n_421)
);

AOI21x1_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_555),
.B(n_567),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_513),
.B(n_554),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_472),
.B(n_512),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_455),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_426),
.B(n_455),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_442),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_427),
.A2(n_442),
.B1(n_443),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_427),
.Y(n_488)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx8_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_465),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_456),
.B(n_466),
.C(n_471),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_457),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_471),
.Y(n_465)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_467),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_470),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_473),
.A2(n_489),
.B(n_511),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_487),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_487),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_505),
.B(n_510),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_500),
.Y(n_490)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_509),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_509),
.Y(n_510)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_553),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_514),
.B(n_553),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_532),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_526),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_516),
.B(n_526),
.C(n_532),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_518),
.Y(n_561)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

XOR2x2_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_551),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_533),
.B(n_551),
.Y(n_559)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_548),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_556),
.B(n_557),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_556),
.B(n_557),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_558),
.A2(n_562),
.B1(n_563),
.B2(n_566),
.Y(n_557)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_558),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_560),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_560),
.C(n_562),
.Y(n_569)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_570),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_569),
.B(n_570),
.Y(n_573)
);


endmodule