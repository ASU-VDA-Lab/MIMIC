module fake_jpeg_13169_n_399 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_399);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_399;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_6),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_6),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_1),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_62),
.Y(n_100)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_48),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_49),
.Y(n_137)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_63),
.Y(n_92)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_70),
.B1(n_31),
.B2(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_84),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_20),
.A2(n_1),
.B(n_2),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_80),
.Y(n_89)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_87),
.B1(n_27),
.B2(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_6),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_41),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_7),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_86),
.Y(n_128)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_98),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_93),
.A2(n_37),
.B1(n_36),
.B2(n_16),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_69),
.B1(n_54),
.B2(n_46),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_94),
.A2(n_129),
.B1(n_130),
.B2(n_138),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_42),
.B1(n_29),
.B2(n_28),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_95),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_99),
.B(n_106),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_27),
.B1(n_23),
.B2(n_87),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_68),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_32),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_32),
.Y(n_120)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_31),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_38),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_74),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_58),
.B(n_42),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_55),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_139),
.A2(n_178),
.B1(n_182),
.B2(n_185),
.Y(n_186)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_140),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_141),
.A2(n_177),
.B1(n_104),
.B2(n_119),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_93),
.A2(n_75),
.B1(n_51),
.B2(n_57),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_153),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_95),
.A2(n_56),
.B1(n_82),
.B2(n_81),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_89),
.A2(n_41),
.B(n_16),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_150),
.A2(n_92),
.B(n_88),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_86),
.B1(n_85),
.B2(n_72),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_151),
.A2(n_157),
.B1(n_168),
.B2(n_134),
.Y(n_215)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_27),
.B1(n_38),
.B2(n_37),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_110),
.A2(n_16),
.B1(n_37),
.B2(n_36),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_23),
.B1(n_36),
.B2(n_41),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_100),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_150),
.Y(n_212)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_34),
.B1(n_21),
.B2(n_11),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_21),
.B1(n_34),
.B2(n_12),
.Y(n_170)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_88),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_99),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_180),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_109),
.A2(n_21),
.B1(n_34),
.B2(n_12),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_183),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_126),
.A2(n_34),
.B1(n_21),
.B2(n_12),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_34),
.C(n_9),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_102),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_216),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_143),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_204),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_195),
.B(n_212),
.Y(n_244)
);

OR2x6_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_170),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_168),
.B1(n_161),
.B2(n_155),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_104),
.B(n_119),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_207),
.B1(n_211),
.B2(n_221),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_155),
.B(n_127),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_205),
.B(n_189),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_148),
.A2(n_125),
.B1(n_121),
.B2(n_134),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_147),
.B(n_127),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_170),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_217),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_139),
.B1(n_124),
.B2(n_149),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_159),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_140),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_122),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_170),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_141),
.A2(n_124),
.B1(n_123),
.B2(n_133),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_139),
.B1(n_177),
.B2(n_132),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_248),
.B1(n_197),
.B2(n_203),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_197),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_191),
.B(n_181),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_251),
.B(n_197),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_139),
.B(n_185),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_232),
.A2(n_250),
.B(n_190),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_152),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_172),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_158),
.B1(n_115),
.B2(n_112),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_249),
.B1(n_190),
.B2(n_202),
.Y(n_275)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_194),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_203),
.C(n_200),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_162),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_222),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_154),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_169),
.B1(n_132),
.B2(n_133),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_208),
.A2(n_180),
.B(n_165),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_213),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_115),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_254),
.C(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_160),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_171),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_257),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_210),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_128),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_259),
.B(n_286),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_229),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_233),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_262),
.B(n_268),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_253),
.A2(n_212),
.B1(n_197),
.B2(n_187),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_274),
.B(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_264),
.A2(n_272),
.B1(n_243),
.B2(n_232),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_278),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_225),
.A2(n_186),
.B1(n_202),
.B2(n_198),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_200),
.B(n_193),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_234),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_193),
.B(n_220),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_239),
.B(n_238),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_222),
.C(n_209),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_285),
.C(n_258),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_253),
.A2(n_220),
.B(n_201),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_226),
.B(n_228),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_261),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_SL g285 ( 
.A(n_251),
.B(n_231),
.C(n_227),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_267),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_231),
.B1(n_251),
.B2(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_296),
.Y(n_315)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_239),
.B1(n_243),
.B2(n_246),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_297),
.B(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_254),
.C(n_257),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_303),
.C(n_304),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_309),
.B1(n_312),
.B2(n_277),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_272),
.A2(n_239),
.B1(n_249),
.B2(n_250),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_274),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_256),
.C(n_242),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_281),
.C(n_285),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_306),
.A2(n_271),
.B(n_260),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_236),
.C(n_230),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_286),
.C(n_259),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_265),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_239),
.B1(n_196),
.B2(n_198),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_273),
.B(n_223),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_269),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_263),
.A2(n_196),
.B1(n_167),
.B2(n_178),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_290),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_320),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_316),
.A2(n_301),
.B1(n_306),
.B2(n_305),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_333),
.C(n_300),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_328),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_289),
.B(n_270),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_292),
.A2(n_276),
.B1(n_269),
.B2(n_268),
.Y(n_321)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_324),
.B(n_331),
.Y(n_339)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_323),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_295),
.A2(n_260),
.B(n_282),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_289),
.B(n_303),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_294),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_265),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_223),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_311),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_267),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_328),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_260),
.B(n_280),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_317),
.B(n_298),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_349),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_308),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_293),
.C(n_308),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_340),
.B(n_341),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_307),
.C(n_297),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_348),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_344),
.A2(n_332),
.B1(n_316),
.B2(n_302),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_292),
.B1(n_312),
.B2(n_309),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_346),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_291),
.C(n_299),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_299),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_350),
.B(n_319),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_314),
.C(n_287),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_347),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_355),
.B(n_363),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_364),
.Y(n_372)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_351),
.Y(n_359)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_359),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_315),
.B1(n_296),
.B2(n_325),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_360),
.A2(n_315),
.B1(n_345),
.B2(n_323),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_349),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_334),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_339),
.A2(n_331),
.B(n_324),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_365),
.A2(n_322),
.B(n_348),
.Y(n_370)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_362),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_338),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_367),
.A2(n_357),
.B1(n_353),
.B2(n_360),
.Y(n_380)
);

AO221x1_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_325),
.B1(n_314),
.B2(n_310),
.C(n_341),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_370),
.B(n_365),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_343),
.C(n_340),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_373),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_356),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_287),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_374),
.B(n_358),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_376),
.B(n_378),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_379),
.B(n_381),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_382),
.C(n_383),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_369),
.A2(n_364),
.B(n_361),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_371),
.A2(n_338),
.B(n_354),
.Y(n_383)
);

AOI322xp5_ASAP7_75t_L g386 ( 
.A1(n_376),
.A2(n_372),
.A3(n_283),
.B1(n_336),
.B2(n_373),
.C1(n_354),
.C2(n_218),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_387),
.Y(n_391)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_372),
.A3(n_283),
.B1(n_218),
.B2(n_201),
.C1(n_145),
.C2(n_176),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_166),
.C(n_90),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_388),
.A2(n_90),
.B(n_118),
.Y(n_392)
);

AOI21x1_ASAP7_75t_L g390 ( 
.A1(n_389),
.A2(n_128),
.B(n_108),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_390),
.A2(n_393),
.B(n_384),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_118),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_395),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_396),
.A2(n_391),
.B(n_12),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_L g398 ( 
.A(n_397),
.B(n_7),
.C(n_13),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_398),
.A2(n_13),
.B1(n_14),
.B2(n_214),
.Y(n_399)
);


endmodule