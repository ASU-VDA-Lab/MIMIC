module fake_jpeg_8818_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx2_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_26),
.B1(n_20),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_23),
.B1(n_16),
.B2(n_25),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_24),
.B1(n_17),
.B2(n_21),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_32),
.B1(n_36),
.B2(n_30),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_22),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_70),
.B1(n_75),
.B2(n_49),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_22),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_68),
.B(n_72),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_54),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_59),
.Y(n_94)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_14),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_61),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_12),
.C(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_15),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_16),
.B1(n_23),
.B2(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_18),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_17),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_59),
.C(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_27),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_91),
.C(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_50),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_96),
.B1(n_58),
.B2(n_52),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_35),
.C(n_33),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_105),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_51),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_108),
.C(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_106),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_107),
.B(n_113),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_73),
.B(n_70),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_109),
.B(n_111),
.Y(n_119)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_68),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_27),
.B(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_56),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_112),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_21),
.B(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_27),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_21),
.B(n_27),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_115),
.B(n_21),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_27),
.B(n_21),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_118),
.C(n_125),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_80),
.C(n_81),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_126),
.Y(n_139)
);

AO22x2_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_90),
.B1(n_89),
.B2(n_81),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_128),
.B(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_80),
.C(n_82),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_93),
.B1(n_88),
.B2(n_92),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_24),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_92),
.B(n_90),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_24),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_98),
.C(n_104),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_1),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_140),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_102),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_124),
.Y(n_149)
);

OAI322xp33_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_100),
.A3(n_107),
.B1(n_101),
.B2(n_115),
.C1(n_114),
.C2(n_113),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_143),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_103),
.B1(n_97),
.B2(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_12),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_123),
.B(n_128),
.Y(n_143)
);

NAND5xp2_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_124),
.C(n_129),
.D(n_125),
.E(n_131),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_133),
.B(n_3),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_124),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.C(n_152),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_1),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_158),
.B(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_144),
.A2(n_132),
.B1(n_133),
.B2(n_5),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_152),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_159),
.B(n_5),
.Y(n_164)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_149),
.C(n_146),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_6),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_5),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_157),
.B1(n_155),
.B2(n_7),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_7),
.A3(n_8),
.B1(n_122),
.B2(n_148),
.C1(n_135),
.C2(n_126),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_166),
.C(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_167),
.Y(n_176)
);


endmodule