module fake_jpeg_23632_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_16),
.B1(n_19),
.B2(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_21),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_13),
.B(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_26),
.B1(n_19),
.B2(n_17),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_30),
.C(n_32),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_30),
.C(n_16),
.Y(n_72)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_53),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_57)
);

NOR2x1p5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_31),
.B1(n_34),
.B2(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_28),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_77),
.C(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_76),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_28),
.C(n_22),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_29),
.C(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_63),
.B1(n_61),
.B2(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_93),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_96),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_83),
.B(n_71),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_52),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_95),
.B1(n_86),
.B2(n_85),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_48),
.B1(n_69),
.B2(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_62),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_64),
.B(n_68),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_75),
.C(n_80),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_15),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_86),
.B(n_72),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_97),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_107),
.B1(n_110),
.B2(n_93),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_27),
.B1(n_15),
.B2(n_23),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_25),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_114),
.C(n_117),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_116),
.B1(n_104),
.B2(n_100),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_88),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_104),
.C(n_107),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_108),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_121),
.B(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_14),
.Y(n_128)
);

AOI211xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_118),
.B(n_113),
.C(n_24),
.Y(n_126)
);

AOI31xp33_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_129),
.A3(n_125),
.B(n_9),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_119),
.C(n_18),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_0),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_23),
.B1(n_18),
.B2(n_8),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_132),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_133),
.A3(n_126),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_4),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.C(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_10),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_2),
.Y(n_138)
);


endmodule