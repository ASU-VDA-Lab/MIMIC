module real_jpeg_26591_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_0),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_0),
.A2(n_54),
.B1(n_56),
.B2(n_172),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_172),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_172),
.Y(n_312)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_2),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_31),
.B1(n_54),
.B2(n_56),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_54),
.B1(n_56),
.B2(n_83),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_83),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_83),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_5),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_54),
.B1(n_56),
.B2(n_155),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_155),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_155),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_6),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_6),
.A2(n_35),
.B1(n_54),
.B2(n_56),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_8),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_8),
.A2(n_54),
.B1(n_56),
.B2(n_135),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_135),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_135),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_10),
.A2(n_55),
.B(n_56),
.C(n_59),
.D(n_63),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_10),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_80),
.B(n_84),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_25),
.B(n_120),
.C(n_121),
.D(n_125),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_10),
.B(n_25),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_10),
.B(n_21),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_10),
.A2(n_23),
.B(n_29),
.C(n_174),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_102),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_11),
.A2(n_54),
.B1(n_56),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_65),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_65),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_12),
.A2(n_54),
.B1(n_56),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_12),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_76),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_76),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_76),
.Y(n_205)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_13),
.B(n_51),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_13),
.A2(n_56),
.B(n_60),
.C(n_62),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_54),
.B1(n_56),
.B2(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_16),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_30),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_21),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_21),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_21),
.A2(n_26),
.B1(n_205),
.B2(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_21),
.A2(n_26),
.B1(n_34),
.B2(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_22),
.A2(n_25),
.B(n_102),
.Y(n_174)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_24),
.A2(n_25),
.B1(n_72),
.B2(n_123),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_24),
.A2(n_56),
.A3(n_120),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_26),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_26),
.B(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_26),
.Y(n_247)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_33),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_33),
.B(n_339),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_338),
.B(n_340),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_326),
.B(n_337),
.Y(n_39)
);

OAI321xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_290),
.A3(n_319),
.B1(n_324),
.B2(n_325),
.C(n_342),
.Y(n_40)
);

AOI321xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_240),
.A3(n_279),
.B1(n_284),
.B2(n_289),
.C(n_343),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_192),
.C(n_236),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_163),
.B(n_191),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_141),
.B(n_162),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_115),
.B(n_140),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_89),
.B(n_114),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_67),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_48),
.B(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_58),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.A3(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_50),
.B(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_54),
.B(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_59),
.A2(n_62),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_59),
.A2(n_62),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_59),
.A2(n_62),
.B1(n_256),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_63),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_66),
.A2(n_77),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_66),
.A2(n_159),
.B1(n_190),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_66),
.A2(n_159),
.B1(n_214),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_66),
.A2(n_159),
.B(n_265),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_74),
.C(n_79),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_71),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_71),
.A2(n_121),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_71),
.A2(n_121),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_71),
.A2(n_121),
.B1(n_268),
.B2(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_71),
.A2(n_121),
.B(n_331),
.Y(n_330)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_75),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_84),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_80),
.A2(n_88),
.B1(n_134),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_80),
.A2(n_88),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_80),
.A2(n_212),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_80),
.A2(n_97),
.B(n_230),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_105),
.B(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_87),
.A2(n_94),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx5_ASAP7_75t_SL g229 ( 
.A(n_87),
.Y(n_229)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_113),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_98),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_98),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_97),
.B(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_106),
.B(n_112),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_117),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_131),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_128),
.C(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_127),
.A2(n_147),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_127),
.A2(n_200),
.B1(n_226),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_127),
.A2(n_200),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_143),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_156),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_157),
.C(n_158),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_150),
.C(n_153),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_165),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_167),
.B(n_168),
.C(n_177),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_175),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_185),
.C(n_188),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_181),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_187),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_193),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_216),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_194),
.B(n_216),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_209),
.C(n_215),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_198),
.C(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_203),
.B2(n_208),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B(n_202),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_203),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_206),
.B(n_207),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_206),
.A2(n_207),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_206),
.A2(n_247),
.B1(n_275),
.B2(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_206),
.A2(n_247),
.B1(n_302),
.B2(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_215),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_227),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_218),
.B(n_227),
.C(n_235),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_222),
.C(n_224),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_231),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_238),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_260),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_260),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_252),
.C(n_259),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_252),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_251),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_243),
.Y(n_251)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_249),
.C(n_251),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_258),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_258),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g306 ( 
.A1(n_258),
.A2(n_273),
.B(n_276),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_278),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_270),
.B1(n_271),
.B2(n_277),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_266),
.B(n_269),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_266),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_269),
.A2(n_292),
.B1(n_293),
.B2(n_304),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_277),
.C(n_278),
.Y(n_320)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_280),
.A2(n_285),
.B(n_288),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_307),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_307),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_304),
.C(n_305),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_301),
.B2(n_303),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_296),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_300),
.C(n_301),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_297),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_298),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_300),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_311),
.C(n_315),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_301),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_303),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_310),
.C(n_318),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_305),
.A2(n_306),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_318),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_312),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_328),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_336),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_330),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_335),
.C(n_336),
.Y(n_339)
);


endmodule