module fake_jpeg_2254_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_50),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_40),
.B1(n_36),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_49),
.B1(n_51),
.B2(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

BUFx2_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_1),
.Y(n_73)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_72),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_52),
.B1(n_59),
.B2(n_49),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_37),
.B1(n_43),
.B2(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_40),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_41),
.A3(n_37),
.B1(n_43),
.B2(n_4),
.Y(n_76)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AO21x2_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_16),
.B(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_84),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_67),
.B1(n_61),
.B2(n_5),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_1),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_71),
.B(n_2),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_92),
.B1(n_96),
.B2(n_79),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_93),
.B(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_3),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_17),
.C(n_29),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.C(n_22),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_7),
.B(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_9),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_77),
.B(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_103),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_78),
.B(n_80),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_101),
.B(n_9),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_21),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_10),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_25),
.C(n_32),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_108),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_103),
.C(n_11),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_102),
.B(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_114),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

OAI31xp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_106),
.A3(n_11),
.B(n_12),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_12),
.Y(n_120)
);


endmodule