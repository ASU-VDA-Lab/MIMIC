module fake_jpeg_7596_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_149;
wire n_48;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_24),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_8),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_58),
.B1(n_25),
.B2(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_59),
.B1(n_60),
.B2(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_22),
.B1(n_18),
.B2(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_70),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_39),
.B(n_32),
.C(n_17),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_42),
.B(n_17),
.C(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_41),
.B1(n_18),
.B2(n_22),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_58),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_41),
.B1(n_25),
.B2(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_39),
.B1(n_25),
.B2(n_40),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_88),
.B1(n_59),
.B2(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_27),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.C(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_27),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_40),
.B1(n_26),
.B2(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_91),
.B(n_67),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_114),
.B1(n_68),
.B2(n_47),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_106),
.B1(n_110),
.B2(n_79),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_42),
.B(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_0),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_78),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_51),
.B1(n_47),
.B2(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_46),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_46),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_80),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_38),
.B(n_16),
.C(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_116),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_29),
.B1(n_26),
.B2(n_38),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_128),
.Y(n_161)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_121),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_78),
.B1(n_71),
.B2(n_63),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_132),
.B1(n_137),
.B2(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_131),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_78),
.B1(n_63),
.B2(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_111),
.B1(n_108),
.B2(n_107),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_143),
.C(n_23),
.Y(n_171)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_141),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_67),
.B1(n_84),
.B2(n_89),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_84),
.B1(n_70),
.B2(n_85),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_91),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_99),
.B(n_109),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_144),
.B(n_147),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_146),
.B1(n_166),
.B2(n_119),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_106),
.B1(n_90),
.B2(n_99),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_109),
.B(n_103),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_148),
.A2(n_156),
.B(n_159),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_105),
.C(n_15),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_92),
.B1(n_80),
.B2(n_105),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_154),
.B1(n_160),
.B2(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_92),
.B1(n_80),
.B2(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_87),
.B1(n_46),
.B2(n_64),
.Y(n_160)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_171),
.B(n_57),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_103),
.B1(n_38),
.B2(n_48),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_103),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_23),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_153),
.A3(n_151),
.B1(n_171),
.B2(n_162),
.C1(n_135),
.C2(n_159),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_11),
.C(n_13),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_181),
.B1(n_182),
.B2(n_184),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_125),
.B1(n_116),
.B2(n_120),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_178),
.B1(n_185),
.B2(n_192),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_133),
.B1(n_141),
.B2(n_117),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_135),
.B1(n_122),
.B2(n_48),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_48),
.B1(n_127),
.B2(n_57),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_127),
.B1(n_57),
.B2(n_29),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_152),
.B1(n_156),
.B2(n_169),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_160),
.B(n_172),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_26),
.B1(n_29),
.B2(n_16),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_19),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_187),
.C(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_205),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_207),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_189),
.B1(n_186),
.B2(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_166),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_216),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_215),
.C(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_165),
.C(n_144),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_174),
.B(n_16),
.CI(n_19),
.CON(n_218),
.SN(n_218)
);

XNOR2x1_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_202),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_175),
.A2(n_164),
.B1(n_19),
.B2(n_23),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_219),
.A2(n_191),
.B1(n_195),
.B2(n_183),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_223),
.C(n_235),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_174),
.C(n_190),
.Y(n_223)
);

NAND2x1p5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_190),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_232),
.B(n_218),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_179),
.C(n_193),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_226),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_184),
.B1(n_191),
.B2(n_192),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_204),
.B1(n_219),
.B2(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_211),
.B1(n_204),
.B2(n_1),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_30),
.C(n_2),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_201),
.B(n_30),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_213),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_231),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_210),
.C(n_199),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_247),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_199),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_242),
.B(n_245),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_248),
.B1(n_233),
.B2(n_227),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_246),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_202),
.B1(n_3),
.B2(n_1),
.Y(n_248)
);

OAI221xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_224),
.B1(n_232),
.B2(n_225),
.C(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

AO221x1_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_230),
.B1(n_234),
.B2(n_235),
.C(n_231),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_248),
.B1(n_237),
.B2(n_238),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_242),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_14),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_240),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_249),
.B(n_245),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_261),
.Y(n_270)
);

OAI33xp33_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_263),
.A3(n_266),
.B1(n_259),
.B2(n_9),
.B3(n_10),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_237),
.B1(n_6),
.B2(n_7),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_254),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_255),
.C(n_260),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_268),
.C(n_11),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_273),
.B(n_274),
.Y(n_275)
);

OAI221xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_258),
.B1(n_252),
.B2(n_11),
.C(n_12),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_30),
.B(n_10),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.C(n_271),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_7),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_275),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_280),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_13),
.B(n_30),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_13),
.Y(n_284)
);


endmodule