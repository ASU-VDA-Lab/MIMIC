module real_jpeg_31680_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_648;
wire n_95;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_578;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_634;
wire n_153;
wire n_104;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_469;
wire n_98;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_650;
wire n_250;
wire n_254;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_602;
wire n_293;
wire n_56;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_597;
wire n_42;
wire n_313;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_641;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_0),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_1),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_341)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_1),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_1),
.A2(n_345),
.B1(n_470),
.B2(n_472),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_1),
.A2(n_345),
.B1(n_524),
.B2(n_526),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_SL g601 ( 
.A1(n_1),
.A2(n_345),
.B1(n_602),
.B2(n_604),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_2),
.B(n_655),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_3),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_3),
.A2(n_158),
.B1(n_264),
.B2(n_268),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_3),
.A2(n_158),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_3),
.A2(n_158),
.B1(n_333),
.B2(n_499),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_4),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_5),
.A2(n_197),
.B1(n_202),
.B2(n_203),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_5),
.A2(n_202),
.B1(n_379),
.B2(n_381),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_5),
.A2(n_202),
.B1(n_454),
.B2(n_457),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_5),
.A2(n_202),
.B1(n_445),
.B2(n_542),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_64),
.B1(n_69),
.B2(n_71),
.Y(n_63)
);

INVx2_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_71),
.B1(n_166),
.B2(n_169),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_6),
.A2(n_71),
.B1(n_276),
.B2(n_280),
.Y(n_275)
);

AO22x1_ASAP7_75t_L g424 ( 
.A1(n_6),
.A2(n_71),
.B1(n_425),
.B2(n_427),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_6),
.A2(n_71),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_7),
.A2(n_32),
.B1(n_36),
.B2(n_40),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_7),
.A2(n_40),
.B1(n_117),
.B2(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_7),
.A2(n_40),
.B1(n_247),
.B2(n_251),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_7),
.A2(n_40),
.B1(n_371),
.B2(n_373),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_8),
.A2(n_100),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_8),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_8),
.A2(n_142),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_8),
.A2(n_142),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_8),
.A2(n_142),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_9),
.A2(n_409),
.B1(n_411),
.B2(n_414),
.Y(n_408)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_9),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_9),
.A2(n_381),
.B1(n_414),
.B2(n_491),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_9),
.A2(n_414),
.B1(n_576),
.B2(n_578),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_9),
.A2(n_414),
.B1(n_623),
.B2(n_626),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_10),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_10),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_10),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_11),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_13),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_13),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_13),
.A2(n_288),
.B1(n_403),
.B2(n_405),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_13),
.A2(n_288),
.B1(n_506),
.B2(n_507),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_13),
.A2(n_288),
.B1(n_542),
.B2(n_566),
.Y(n_565)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_14),
.Y(n_93)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g463 ( 
.A1(n_15),
.A2(n_411),
.B1(n_464),
.B2(n_467),
.Y(n_463)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_15),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_15),
.A2(n_214),
.B1(n_467),
.B2(n_532),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g593 ( 
.A1(n_15),
.A2(n_467),
.B1(n_594),
.B2(n_597),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_15),
.A2(n_467),
.B1(n_634),
.B2(n_637),
.Y(n_633)
);

OAI221xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_21),
.B1(n_648),
.B2(n_656),
.C(n_657),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_16),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_17),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_17),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_17),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_18),
.Y(n_212)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_18),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_18),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_18),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_19),
.A2(n_31),
.B1(n_41),
.B2(n_46),
.Y(n_30)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_19),
.B(n_173),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_19),
.A2(n_206),
.A3(n_208),
.B1(n_213),
.B2(n_218),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_19),
.A2(n_54),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_19),
.B(n_333),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_19),
.A2(n_332),
.B(n_356),
.Y(n_355)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_21),
.B(n_650),
.C(n_654),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_555),
.B(n_641),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_394),
.B(n_550),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_307),
.B(n_393),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_256),
.B(n_306),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_185),
.B(n_255),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_148),
.Y(n_26)
);

AOI21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_84),
.B(n_145),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_61),
.B(n_83),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_52),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_31),
.A2(n_46),
.B1(n_63),
.B2(n_72),
.Y(n_62)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_35),
.Y(n_344)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_35),
.Y(n_413)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_35),
.Y(n_466)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_41),
.A2(n_46),
.B1(n_408),
.B2(n_462),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_45),
.Y(n_152)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_45),
.Y(n_418)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_46),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_46),
.A2(n_140),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_46),
.A2(n_341),
.B1(n_408),
.B2(n_415),
.Y(n_407)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_46),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_49),
.Y(n_195)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_49),
.Y(n_339)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g60 ( 
.A(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_51),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_96),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_SL g128 ( 
.A1(n_54),
.A2(n_95),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_54),
.B(n_214),
.Y(n_213)
);

NOR2xp67_ASAP7_75t_R g292 ( 
.A(n_54),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_56),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_57),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_74),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_67),
.Y(n_290)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_75),
.A2(n_133),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_75),
.A2(n_133),
.B1(n_263),
.B2(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_75),
.A2(n_133),
.B1(n_378),
.B2(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_75),
.A2(n_133),
.B1(n_402),
.B2(n_469),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_75),
.A2(n_133),
.B1(n_469),
.B2(n_490),
.Y(n_489)
);

AO21x2_ASAP7_75t_L g571 ( 
.A1(n_75),
.A2(n_133),
.B(n_531),
.Y(n_571)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AO21x2_ASAP7_75t_L g133 ( 
.A1(n_76),
.A2(n_105),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_76)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_138),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_113),
.B1(n_114),
.B2(n_137),
.Y(n_85)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_86),
.B(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_94),
.B1(n_99),
.B2(n_104),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_98),
.Y(n_217)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_109),
.Y(n_385)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_137),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_128),
.B2(n_132),
.Y(n_114)
);

NAND2x1_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_165),
.Y(n_164)
);

AOI22x1_ASAP7_75t_L g227 ( 
.A1(n_115),
.A2(n_132),
.B1(n_165),
.B2(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_115),
.A2(n_132),
.B1(n_530),
.B2(n_535),
.Y(n_529)
);

NAND2x1_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_154),
.B1(n_193),
.B2(n_196),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_143),
.A2(n_196),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_143),
.A2(n_287),
.B1(n_337),
.B2(n_340),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_162),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_172),
.C(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B(n_172),
.C(n_184),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_164),
.C(n_172),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_R g189 ( 
.A(n_163),
.B(n_164),
.Y(n_189)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_168),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_171),
.Y(n_406)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

AOI22x1_ASAP7_75t_L g502 ( 
.A1(n_173),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_173),
.A2(n_503),
.B1(n_505),
.B2(n_523),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_SL g618 ( 
.A1(n_173),
.A2(n_503),
.B(n_619),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AO21x2_ASAP7_75t_L g233 ( 
.A1(n_174),
.A2(n_218),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_181),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_175),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_175),
.Y(n_492)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2x1_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_188),
.B(n_190),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_225),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_191),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_205),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_205),
.Y(n_260)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_210),
.Y(n_244)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_211),
.Y(n_433)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_212),
.Y(n_599)
);

INVx3_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_220),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_227),
.B(n_231),
.C(n_305),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_233),
.A2(n_245),
.B1(n_246),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_233),
.A2(n_245),
.B1(n_275),
.B2(n_387),
.Y(n_386)
);

OA22x2_ASAP7_75t_L g431 ( 
.A1(n_233),
.A2(n_245),
.B1(n_387),
.B2(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_233),
.A2(n_245),
.B1(n_432),
.B2(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_233),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_233),
.A2(n_245),
.B1(n_574),
.B2(n_575),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_233),
.A2(n_245),
.B1(n_575),
.B2(n_593),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_235),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_247),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_249),
.Y(n_316)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_249),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_254),
.Y(n_510)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_254),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_304),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_304),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_272),
.B2(n_273),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_270),
.B2(n_271),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_261),
.B(n_271),
.C(n_272),
.Y(n_392)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_267),
.Y(n_474)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_267),
.Y(n_534)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_274),
.B(n_292),
.C(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_279),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_282),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_292),
.Y(n_283)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

BUFx4f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_293),
.A2(n_355),
.B1(n_359),
.B2(n_370),
.Y(n_354)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_293),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_293),
.A2(n_359),
.B1(n_442),
.B2(n_449),
.Y(n_441)
);

OAI22x1_ASAP7_75t_SL g496 ( 
.A1(n_293),
.A2(n_359),
.B1(n_442),
.B2(n_497),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_293),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_294),
.B(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_298),
.B1(n_302),
.B2(n_303),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_299),
.Y(n_525)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_300),
.Y(n_577)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_300),
.Y(n_579)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_300),
.Y(n_596)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_392),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_308),
.B(n_392),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_352),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_350),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_310),
.B(n_350),
.C(n_352),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_336),
.B1(n_348),
.B2(n_349),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_311),
.B(n_349),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_311),
.B(n_349),
.Y(n_459)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_314),
.A3(n_317),
.B1(n_324),
.B2(n_331),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_322),
.Y(n_426)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_322),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_323),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_335),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_335),
.Y(n_636)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_344),
.Y(n_347)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

BUFx2_ASAP7_75t_SL g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_376),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_SL g399 ( 
.A(n_354),
.B(n_377),
.C(n_386),
.Y(n_399)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_359),
.A2(n_601),
.B1(n_607),
.B2(n_608),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_359),
.A2(n_601),
.B1(n_621),
.B2(n_622),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_359),
.Y(n_632)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_360),
.A2(n_423),
.B1(n_424),
.B2(n_430),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_360),
.A2(n_423),
.B1(n_498),
.B2(n_541),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_360),
.A2(n_423),
.B1(n_541),
.B2(n_565),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_365),
.B2(n_367),
.Y(n_361)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_362),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_362),
.Y(n_451)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_368),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_368),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_369),
.Y(n_372)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_369),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_369),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_369),
.Y(n_628)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_375),
.Y(n_448)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_375),
.Y(n_501)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_375),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_386),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND4xp25_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_435),
.C(n_513),
.D(n_545),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_396),
.B(n_397),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_419),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_399),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_400),
.B(n_419),
.C(n_547),
.Y(n_546)
);

XOR2x2_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_407),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_407),
.Y(n_439)
);

BUFx6f_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2x1_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_431),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_431),
.C(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_423),
.Y(n_607)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

A2O1A1O1Ixp25_ASAP7_75t_L g550 ( 
.A1(n_435),
.A2(n_513),
.B(n_551),
.C(n_553),
.D(n_554),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_475),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_436),
.B(n_475),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_458),
.C(n_460),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_438),
.B(n_460),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_477),
.C(n_479),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_452),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_441),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_447),
.Y(n_639)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_452),
.Y(n_479)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_453),
.Y(n_504)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_458),
.B(n_549),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_468),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_468),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_463),
.A2(n_484),
.B(n_486),
.Y(n_483)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx4f_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_476),
.B(n_481),
.C(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_493),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_483),
.B1(n_487),
.B2(n_488),
.Y(n_481)
);

XNOR2x1_ASAP7_75t_L g539 ( 
.A(n_482),
.B(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_489),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_483),
.A2(n_540),
.B(n_582),
.Y(n_581)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_493),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_494),
.A2(n_495),
.B1(n_511),
.B2(n_512),
.Y(n_493)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_495),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_502),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_496),
.Y(n_519)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_502),
.Y(n_518)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_518),
.C(n_519),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_516),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_516),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_517),
.B(n_559),
.C(n_560),
.Y(n_558)
);

XOR2x1_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_537),
.Y(n_520)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_521),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_529),
.B(n_536),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_529),
.Y(n_536)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_527),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_534),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_536),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_537),
.Y(n_559)
);

XNOR2x1_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_539),
.Y(n_537)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_548),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_546),
.B(n_548),
.C(n_552),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_556),
.B(n_609),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_584),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_561),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_558),
.B(n_561),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_580),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_581),
.C(n_583),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_569),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_570),
.C(n_573),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_564),
.B(n_590),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_564),
.B(n_588),
.C(n_590),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_565),
.Y(n_608)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_570),
.A2(n_571),
.B1(n_572),
.B2(n_573),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

XNOR2x1_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_592),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_571),
.B(n_600),
.C(n_615),
.Y(n_614)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_583),
.Y(n_580)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_585),
.A2(n_644),
.B(n_645),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_587),
.Y(n_585)
);

NOR2x1_ASAP7_75t_L g645 ( 
.A(n_586),
.B(n_587),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_589),
.Y(n_587)
);

XOR2x1_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_600),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_592),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_593),
.Y(n_619)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx8_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_610),
.B(n_630),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_611),
.A2(n_643),
.B(n_646),
.Y(n_642)
);

NOR2x1_ASAP7_75t_R g611 ( 
.A(n_612),
.B(n_629),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_612),
.B(n_629),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_613),
.A2(n_614),
.B1(n_616),
.B2(n_617),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_613),
.B(n_618),
.C(n_620),
.Y(n_640)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_620),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_621),
.A2(n_622),
.B1(n_632),
.B2(n_633),
.Y(n_631)
);

AO21x1_ASAP7_75t_L g652 ( 
.A1(n_621),
.A2(n_632),
.B(n_633),
.Y(n_652)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_628),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_630),
.A2(n_642),
.B(n_647),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_631),
.B(n_640),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_631),
.B(n_640),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_631),
.B(n_652),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_631),
.B(n_652),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_635),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_649),
.B(n_654),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_651),
.B(n_653),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_654),
.Y(n_656)
);


endmodule