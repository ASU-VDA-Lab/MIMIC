module fake_aes_1975_n_646 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_646);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_646;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_420;
wire n_446;
wire n_165;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g75 ( .A(n_15), .Y(n_75) );
INVxp67_ASAP7_75t_L g76 ( .A(n_45), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_42), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_23), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_0), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_53), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_37), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_6), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_40), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_27), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_12), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_33), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_47), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_61), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_32), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_17), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_49), .Y(n_93) );
CKINVDCx14_ASAP7_75t_R g94 ( .A(n_10), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_69), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_50), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g97 ( .A(n_51), .B(n_14), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_36), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_0), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_74), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_57), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_13), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_10), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_21), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_56), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_34), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_16), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_66), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_43), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_16), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_13), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_6), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_62), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_25), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_94), .B(n_1), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_81), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_94), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_105), .B(n_1), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_110), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_106), .B(n_2), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
AND2x6_ASAP7_75t_L g137 ( .A(n_108), .B(n_30), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_99), .B(n_3), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
INVxp33_ASAP7_75t_SL g140 ( .A(n_96), .Y(n_140) );
INVx6_ASAP7_75t_L g141 ( .A(n_108), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_81), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_75), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_86), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_75), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_79), .B(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_82), .B(n_5), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_119), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_84), .B(n_5), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_88), .B(n_38), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_100), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_84), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_87), .B(n_7), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_75), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_125), .B(n_120), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_125), .B(n_96), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
INVx1_ASAP7_75t_SL g166 ( .A(n_140), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
INVx1_ASAP7_75t_SL g168 ( .A(n_134), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
AOI21x1_ASAP7_75t_L g170 ( .A1(n_123), .A2(n_118), .B(n_100), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_160), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_121), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_147), .B(n_87), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_123), .B(n_76), .Y(n_181) );
AO22x2_ASAP7_75t_L g182 ( .A1(n_147), .A2(n_117), .B1(n_116), .B2(n_115), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_132), .B(n_109), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_157), .B(n_114), .Y(n_185) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_157), .B(n_97), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_128), .B(n_113), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_128), .B(n_112), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_129), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_124), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_126), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_156), .B(n_104), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_130), .B(n_103), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_130), .A2(n_110), .B1(n_111), .B2(n_102), .Y(n_201) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_149), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_135), .B(n_107), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_150), .Y(n_206) );
NOR2xp33_ASAP7_75t_SL g207 ( .A(n_153), .B(n_101), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_136), .B(n_98), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_136), .B(n_95), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_124), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_139), .B(n_92), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_149), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_139), .B(n_93), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_202), .B(n_144), .Y(n_215) );
OR2x6_ASAP7_75t_L g216 ( .A(n_182), .B(n_151), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_175), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_205), .B(n_144), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_205), .B(n_159), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_196), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_198), .B(n_133), .C(n_148), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_169), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_183), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_162), .Y(n_226) );
INVx5_ASAP7_75t_L g227 ( .A(n_175), .Y(n_227) );
BUFx12f_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_182), .Y(n_229) );
OR2x2_ASAP7_75t_SL g230 ( .A(n_166), .B(n_133), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_182), .Y(n_231) );
INVx5_ASAP7_75t_L g232 ( .A(n_175), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_169), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_167), .B(n_158), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_168), .B(n_151), .Y(n_236) );
AND2x6_ASAP7_75t_L g237 ( .A(n_190), .B(n_152), .Y(n_237) );
AND3x1_ASAP7_75t_SL g238 ( .A(n_196), .B(n_152), .C(n_158), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_161), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_162), .B(n_159), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_205), .B(n_150), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g243 ( .A1(n_167), .A2(n_138), .B1(n_78), .B2(n_77), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_190), .A2(n_89), .B(n_90), .C(n_91), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_181), .B(n_150), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_179), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_186), .B(n_149), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_199), .B(n_149), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_171), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_172), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_201), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_176), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_176), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_177), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_199), .B(n_7), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_177), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_193), .A2(n_153), .B1(n_137), .B2(n_141), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_162), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_189), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_186), .B(n_153), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_179), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_191), .B(n_129), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_164), .Y(n_269) );
INVx5_ASAP7_75t_L g270 ( .A(n_213), .Y(n_270) );
INVx5_ASAP7_75t_L g271 ( .A(n_213), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_163), .B(n_141), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_237), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_218), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g275 ( .A(n_225), .B(n_180), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_216), .A2(n_193), .B1(n_184), .B2(n_180), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_269), .B(n_185), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_216), .A2(n_185), .B1(n_208), .B2(n_153), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_215), .B(n_185), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_268), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_239), .Y(n_281) );
AOI21x1_ASAP7_75t_L g282 ( .A1(n_266), .A2(n_203), .B(n_212), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_239), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_215), .B(n_208), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_226), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_236), .B(n_200), .Y(n_286) );
NAND2x2_ASAP7_75t_L g287 ( .A(n_259), .B(n_214), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_228), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_216), .A2(n_207), .B1(n_200), .B2(n_209), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_253), .Y(n_290) );
BUFx12f_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_235), .B(n_188), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
CKINVDCx8_ASAP7_75t_R g294 ( .A(n_248), .Y(n_294) );
BUFx12f_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_235), .B(n_187), .Y(n_296) );
AND2x6_ASAP7_75t_L g297 ( .A(n_220), .B(n_191), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_223), .A2(n_192), .B1(n_191), .B2(n_204), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_222), .Y(n_299) );
OAI22x1_ASAP7_75t_L g300 ( .A1(n_255), .A2(n_192), .B1(n_204), .B2(n_11), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_229), .A2(n_192), .B1(n_204), .B2(n_137), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_272), .B(n_206), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_243), .B(n_203), .Y(n_304) );
CKINVDCx12_ASAP7_75t_R g305 ( .A(n_272), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_254), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_257), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_243), .B(n_141), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_226), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_257), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_237), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_222), .B(n_251), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_217), .Y(n_313) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_272), .B(n_146), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_217), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_231), .B(n_137), .Y(n_316) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_238), .A2(n_237), .B1(n_219), .B2(n_264), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_226), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_304), .A2(n_237), .B1(n_260), .B2(n_267), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_294), .B(n_249), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_291), .A2(n_237), .B1(n_227), .B2(n_232), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_273), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_274), .B(n_258), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_274), .A2(n_244), .B1(n_258), .B2(n_263), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_312), .A2(n_227), .B1(n_232), .B2(n_247), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_304), .A2(n_252), .B1(n_240), .B2(n_256), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_273), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_281), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_284), .B(n_263), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_279), .A2(n_246), .B1(n_242), .B2(n_227), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_283), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_287), .A2(n_227), .B1(n_232), .B2(n_241), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_276), .A2(n_244), .B1(n_233), .B2(n_221), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_287), .A2(n_232), .B1(n_241), .B2(n_250), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_273), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_290), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_277), .A2(n_270), .B1(n_250), .B2(n_271), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_286), .B(n_233), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_273), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_276), .A2(n_221), .B1(n_261), .B2(n_238), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_311), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g345 ( .A1(n_317), .A2(n_261), .B1(n_245), .B2(n_141), .C(n_271), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_295), .A2(n_137), .B1(n_160), .B2(n_250), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_293), .B(n_226), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_319), .A2(n_278), .B1(n_289), .B2(n_317), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_333), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_324), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_324), .B(n_293), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_324), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_330), .A2(n_311), .B1(n_299), .B2(n_295), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_329), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_330), .A2(n_278), .B(n_306), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_333), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_341), .B(n_280), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_327), .A2(n_292), .B1(n_296), .B2(n_277), .C(n_300), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_320), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_341), .B(n_306), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_327), .A2(n_302), .B1(n_275), .B2(n_314), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_322), .Y(n_364) );
BUFx12f_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_322), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_L g369 ( .A1(n_345), .A2(n_308), .B(n_303), .C(n_307), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_332), .Y(n_370) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_337), .A2(n_288), .B(n_301), .C(n_298), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_319), .A2(n_305), .B1(n_275), .B2(n_302), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_339), .B(n_310), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_354), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_354), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_361), .B(n_334), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_351), .B(n_339), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_360), .A2(n_325), .B1(n_326), .B2(n_343), .C(n_345), .Y(n_378) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_372), .A2(n_343), .B1(n_325), .B2(n_346), .C1(n_336), .C2(n_321), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_350), .B(n_333), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_336), .B1(n_331), .B2(n_340), .C(n_314), .Y(n_382) );
AOI21xp33_ASAP7_75t_SL g383 ( .A1(n_348), .A2(n_344), .B(n_9), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_365), .A2(n_322), .B1(n_342), .B2(n_338), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_335), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_335), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_364), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_331), .B1(n_335), .B2(n_346), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_356), .B(n_328), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_301), .B1(n_344), .B2(n_313), .C(n_315), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_370), .B(n_347), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_349), .Y(n_395) );
OA21x2_ASAP7_75t_L g396 ( .A1(n_369), .A2(n_282), .B(n_142), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_368), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
OR2x6_ASAP7_75t_L g400 ( .A(n_367), .B(n_344), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_371), .A2(n_315), .B1(n_313), .B2(n_338), .C(n_328), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_359), .A2(n_297), .B1(n_347), .B2(n_338), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_361), .B(n_328), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_366), .B(n_347), .Y(n_406) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_381), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_383), .A2(n_359), .B1(n_357), .B2(n_362), .C(n_373), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_383), .A2(n_362), .B(n_359), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_374), .B(n_364), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_385), .B(n_362), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_376), .A2(n_367), .B1(n_316), .B2(n_364), .Y(n_414) );
AOI33xp33_ASAP7_75t_L g415 ( .A1(n_375), .A2(n_122), .A3(n_142), .B1(n_145), .B2(n_197), .B3(n_211), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_385), .B(n_364), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_377), .B(n_364), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_389), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_377), .B(n_145), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_378), .A2(n_342), .B1(n_316), .B2(n_137), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_394), .B(n_8), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_391), .A2(n_379), .B(n_395), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_127), .B1(n_124), .B2(n_143), .C(n_146), .Y(n_427) );
OR2x2_ASAP7_75t_SL g428 ( .A(n_380), .B(n_397), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_387), .B(n_145), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_387), .B(n_398), .Y(n_431) );
AOI21xp5_ASAP7_75t_SL g432 ( .A1(n_400), .A2(n_382), .B(n_342), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_394), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_404), .B(n_8), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_389), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_390), .A2(n_309), .B(n_285), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_395), .A2(n_309), .B(n_285), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_404), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_399), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_399), .Y(n_441) );
NOR2x1_ASAP7_75t_R g442 ( .A(n_402), .B(n_318), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_392), .B(n_55), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_406), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_406), .B(n_11), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_392), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_405), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_384), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_403), .B(n_400), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_400), .B(n_142), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_400), .B(n_14), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_396), .B(n_15), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_431), .B(n_396), .Y(n_454) );
NOR3xp33_ASAP7_75t_SL g455 ( .A(n_452), .B(n_401), .C(n_393), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_433), .B(n_396), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_431), .B(n_396), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_445), .B(n_122), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_419), .B(n_421), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_445), .B(n_122), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_420), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_426), .B(n_124), .C(n_127), .D(n_143), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_412), .B(n_160), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
AND3x2_ASAP7_75t_L g469 ( .A(n_432), .B(n_18), .C(n_19), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_420), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_412), .B(n_146), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_422), .B(n_131), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_411), .B(n_146), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_417), .B(n_143), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_422), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_410), .Y(n_476) );
AO22x1_ASAP7_75t_L g477 ( .A1(n_449), .A2(n_297), .B1(n_137), .B2(n_143), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_407), .B(n_127), .Y(n_478) );
INVx4_ASAP7_75t_L g479 ( .A(n_443), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_417), .B(n_127), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_416), .B(n_131), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_428), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_451), .B(n_131), .C(n_129), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_408), .A2(n_137), .B1(n_131), .B2(n_129), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_429), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_418), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_446), .B(n_131), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_425), .B(n_131), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_441), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_409), .A2(n_137), .B1(n_297), .B2(n_318), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_444), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_409), .A2(n_297), .B1(n_318), .B2(n_309), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_416), .B(n_20), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g499 ( .A1(n_435), .A2(n_297), .B1(n_266), .B2(n_270), .C1(n_250), .C2(n_271), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_443), .B(n_318), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_440), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_446), .B(n_309), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_22), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_448), .B(n_24), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_425), .B(n_26), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_430), .B(n_28), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_423), .B(n_29), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_423), .B(n_285), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_468), .B(n_432), .C(n_450), .D(n_414), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_462), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_464), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_464), .B(n_447), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_484), .A2(n_442), .B(n_409), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_462), .B(n_487), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_488), .B(n_410), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_470), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_488), .B(n_410), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_476), .B(n_462), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_489), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_471), .B(n_447), .Y(n_520) );
NOR2x1p5_ASAP7_75t_L g521 ( .A(n_479), .B(n_443), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_456), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_457), .B(n_430), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_459), .B(n_436), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_466), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_475), .Y(n_526) );
NAND4xp75_ASAP7_75t_L g527 ( .A(n_455), .B(n_451), .C(n_436), .D(n_427), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_482), .B(n_418), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_470), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_460), .B(n_453), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_481), .B(n_453), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_505), .B(n_438), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_483), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_491), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_479), .B(n_415), .Y(n_536) );
AND4x1_ASAP7_75t_L g537 ( .A(n_455), .B(n_424), .C(n_437), .D(n_44), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g538 ( .A(n_479), .B(n_35), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_481), .B(n_39), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_476), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_501), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_474), .B(n_48), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_480), .B(n_52), .Y(n_544) );
AND3x1_ASAP7_75t_L g545 ( .A(n_504), .B(n_498), .C(n_497), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_478), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_476), .B(n_58), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_454), .B(n_60), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_473), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_493), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_477), .A2(n_285), .B(n_224), .Y(n_551) );
OAI22xp33_ASAP7_75t_L g552 ( .A1(n_500), .A2(n_271), .B1(n_270), .B2(n_234), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_454), .B(n_63), .Y(n_553) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_498), .B(n_234), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
AOI21xp33_ASAP7_75t_SL g556 ( .A1(n_500), .A2(n_64), .B(n_65), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_467), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_495), .B(n_67), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_510), .B(n_496), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_529), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_511), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_518), .B(n_496), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_514), .B(n_458), .Y(n_563) );
XOR2x2_ASAP7_75t_SL g564 ( .A(n_554), .B(n_469), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_546), .B(n_472), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_519), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_549), .B(n_472), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_511), .B(n_472), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_522), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_528), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_525), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_536), .A2(n_465), .B(n_485), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_518), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_526), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_533), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_530), .B(n_502), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_518), .B(n_497), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_515), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_536), .A2(n_490), .B(n_492), .C(n_461), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_554), .A2(n_506), .B1(n_503), .B2(n_507), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_534), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_517), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_535), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_541), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_524), .Y(n_586) );
AND2x2_ASAP7_75t_SL g587 ( .A(n_545), .B(n_494), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_523), .B(n_463), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_512), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_516), .B(n_508), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_516), .B(n_494), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_550), .Y(n_592) );
OAI211xp5_ASAP7_75t_SL g593 ( .A1(n_532), .A2(n_499), .B(n_485), .C(n_469), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_527), .B(n_503), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_531), .B(n_557), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_555), .Y(n_596) );
AOI211xp5_ASAP7_75t_SL g597 ( .A1(n_538), .A2(n_68), .B(n_70), .C(n_72), .Y(n_597) );
AOI322xp5_ASAP7_75t_L g598 ( .A1(n_520), .A2(n_173), .A3(n_174), .B1(n_210), .B2(n_194), .C1(n_211), .C2(n_197), .Y(n_598) );
XNOR2x1_ASAP7_75t_L g599 ( .A(n_521), .B(n_73), .Y(n_599) );
XNOR2xp5_ASAP7_75t_L g600 ( .A(n_537), .B(n_224), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_194), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_532), .B(n_210), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_529), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_542), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_520), .A2(n_173), .B1(n_174), .B2(n_165), .C1(n_178), .C2(n_195), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g607 ( .A1(n_513), .A2(n_270), .B(n_178), .C(n_195), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_540), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_509), .A2(n_165), .B1(n_178), .B2(n_195), .C(n_262), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_553), .B(n_165), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_548), .A2(n_165), .B(n_178), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_556), .A2(n_165), .B(n_178), .C(n_195), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_558), .B(n_195), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_543), .A2(n_262), .B1(n_539), .B2(n_544), .C(n_547), .Y(n_614) );
OAI22xp5_ASAP7_75t_SL g615 ( .A1(n_587), .A2(n_580), .B1(n_594), .B2(n_570), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_586), .A2(n_584), .B1(n_589), .B2(n_566), .C(n_574), .Y(n_616) );
AO22x2_ASAP7_75t_L g617 ( .A1(n_608), .A2(n_571), .B1(n_581), .B2(n_575), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_579), .A2(n_587), .B(n_602), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g619 ( .A1(n_564), .A2(n_573), .B1(n_572), .B2(n_561), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_569), .A2(n_583), .B1(n_585), .B2(n_561), .C(n_563), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_577), .A2(n_593), .B1(n_565), .B2(n_562), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g622 ( .A1(n_607), .A2(n_609), .B(n_612), .C(n_591), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_582), .A2(n_578), .B1(n_599), .B2(n_595), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_576), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_560), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_576), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_577), .A2(n_591), .B1(n_567), .B2(n_568), .C(n_614), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g628 ( .A(n_623), .B(n_597), .C(n_605), .Y(n_628) );
XNOR2xp5_ASAP7_75t_L g629 ( .A(n_615), .B(n_600), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_621), .A2(n_590), .B1(n_588), .B2(n_564), .C(n_562), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_620), .B(n_592), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_619), .A2(n_596), .B1(n_604), .B2(n_603), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_618), .A2(n_559), .B1(n_560), .B2(n_606), .C(n_610), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_627), .A2(n_597), .B1(n_611), .B2(n_610), .C(n_605), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_631), .B(n_616), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_630), .A2(n_617), .B1(n_626), .B2(n_624), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_628), .Y(n_637) );
OAI322xp33_ASAP7_75t_L g638 ( .A1(n_629), .A2(n_632), .A3(n_634), .B1(n_633), .B2(n_625), .C1(n_622), .C2(n_617), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_637), .Y(n_639) );
OR4x2_ASAP7_75t_L g640 ( .A(n_638), .B(n_559), .C(n_552), .D(n_598), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_639), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_640), .A2(n_636), .B1(n_635), .B2(n_613), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_641), .B(n_640), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g644 ( .A(n_643), .B(n_642), .C(n_601), .D(n_551), .Y(n_644) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_644), .A2(n_643), .B1(n_552), .B2(n_558), .Y(n_645) );
AOI21xp33_ASAP7_75t_SL g646 ( .A1(n_645), .A2(n_262), .B(n_637), .Y(n_646) );
endmodule