module fake_netlist_1_11875_n_658 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_658);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_658;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_631;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
OR2x2_ASAP7_75t_L g74 ( .A(n_44), .B(n_43), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_65), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_33), .Y(n_76) );
INVxp67_ASAP7_75t_L g77 ( .A(n_57), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_30), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_39), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_29), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_21), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_66), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_7), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_28), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
CKINVDCx14_ASAP7_75t_R g87 ( .A(n_38), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_19), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_16), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_5), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_73), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_42), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_72), .Y(n_94) );
NOR2xp67_ASAP7_75t_L g95 ( .A(n_1), .B(n_40), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_36), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_48), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_56), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_23), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_2), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_0), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_58), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_49), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_59), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_18), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_62), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_4), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_32), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_52), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_63), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_34), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_3), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_37), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_17), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_27), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_117), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_94), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_121) );
CKINVDCx11_ASAP7_75t_R g122 ( .A(n_90), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_84), .B(n_4), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_75), .B(n_5), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_83), .A2(n_41), .B(n_69), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_117), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_99), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_127) );
XOR2xp5_ASAP7_75t_L g128 ( .A(n_102), .B(n_8), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_109), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_114), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_102), .B(n_9), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_114), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_75), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_87), .B(n_10), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_109), .B(n_10), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
NAND2xp33_ASAP7_75t_L g141 ( .A(n_114), .B(n_46), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_84), .B(n_11), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_101), .B(n_11), .Y(n_146) );
XNOR2xp5_ASAP7_75t_L g147 ( .A(n_91), .B(n_12), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_112), .A2(n_47), .B(n_68), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_78), .B(n_12), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_82), .B(n_13), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_105), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_76), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_112), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g155 ( .A1(n_104), .A2(n_13), .B1(n_14), .B2(n_20), .Y(n_155) );
CKINVDCx6p67_ASAP7_75t_R g156 ( .A(n_106), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_114), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_76), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_82), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_122), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_139), .B(n_85), .Y(n_161) );
INVx4_ASAP7_75t_SL g162 ( .A(n_151), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_158), .B(n_77), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_120), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_120), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_153), .B(n_95), .Y(n_168) );
INVxp67_ASAP7_75t_SL g169 ( .A(n_135), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_158), .B(n_85), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_153), .B(n_80), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_154), .B(n_86), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_120), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_139), .B(n_86), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_140), .B(n_89), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_145), .B(n_80), .Y(n_181) );
INVx5_ASAP7_75t_L g182 ( .A(n_120), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_137), .A2(n_96), .B1(n_100), .B2(n_93), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_123), .Y(n_184) );
INVxp67_ASAP7_75t_SL g185 ( .A(n_135), .Y(n_185) );
INVx8_ASAP7_75t_L g186 ( .A(n_123), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_134), .B(n_100), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_143), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
OR2x2_ASAP7_75t_L g191 ( .A(n_152), .B(n_129), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_140), .B(n_89), .Y(n_192) );
INVxp33_ASAP7_75t_SL g193 ( .A(n_122), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_134), .Y(n_194) );
AND2x6_ASAP7_75t_L g195 ( .A(n_143), .B(n_111), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_133), .B(n_111), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_120), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_133), .B(n_113), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_136), .B(n_81), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_126), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_138), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_138), .A2(n_96), .B1(n_119), .B2(n_88), .Y(n_205) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_150), .B(n_81), .C(n_93), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_142), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_142), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_130), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_126), .Y(n_212) );
INVx6_ASAP7_75t_L g213 ( .A(n_126), .Y(n_213) );
NOR2x1p5_ASAP7_75t_L g214 ( .A(n_156), .B(n_128), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_126), .B(n_115), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_126), .B(n_115), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_125), .A2(n_103), .B1(n_92), .B2(n_113), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_210), .B(n_124), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_194), .B(n_118), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_213), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_194), .B(n_110), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_190), .A2(n_121), .B1(n_127), .B2(n_155), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_174), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_165), .A2(n_141), .B1(n_157), .B2(n_149), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_205), .A2(n_156), .B1(n_147), .B2(n_128), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_163), .B(n_97), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_179), .A2(n_141), .B1(n_157), .B2(n_125), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_201), .B(n_74), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_169), .B(n_74), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_187), .B(n_108), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_185), .B(n_147), .Y(n_231) );
NAND2xp33_ASAP7_75t_SL g232 ( .A(n_173), .B(n_157), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_163), .B(n_149), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_186), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_168), .B(n_14), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_164), .B(n_148), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_203), .B(n_149), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_164), .B(n_125), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_201), .B(n_148), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_184), .B(n_148), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_191), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_186), .B(n_148), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_186), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_213), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_204), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_171), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_205), .B(n_148), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_172), .B(n_132), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_171), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_188), .Y(n_250) );
OAI22x1_ASAP7_75t_L g251 ( .A1(n_214), .A2(n_22), .B1(n_25), .B2(n_26), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_172), .B(n_132), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_188), .B(n_132), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_195), .A2(n_132), .B1(n_130), .B2(n_45), .Y(n_254) );
INVxp67_ASAP7_75t_L g255 ( .A(n_181), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_206), .B(n_132), .Y(n_256) );
NOR2x1p5_ASAP7_75t_L g257 ( .A(n_193), .B(n_130), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_200), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_195), .B(n_130), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_195), .B(n_130), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_213), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_209), .Y(n_262) );
INVx5_ASAP7_75t_L g263 ( .A(n_195), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_195), .B(n_31), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_204), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_177), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_207), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_177), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_168), .Y(n_269) );
INVxp67_ASAP7_75t_L g270 ( .A(n_192), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_162), .B(n_35), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_207), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_162), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_162), .B(n_50), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_160), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_183), .B(n_51), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_176), .B(n_53), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_255), .A2(n_176), .B1(n_192), .B2(n_178), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_223), .B(n_255), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_241), .B(n_197), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_270), .B(n_178), .Y(n_282) );
BUFx2_ASAP7_75t_SL g283 ( .A(n_243), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_270), .B(n_180), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_237), .A2(n_199), .B(n_197), .C(n_217), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_228), .A2(n_217), .B1(n_180), .B2(n_161), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_238), .A2(n_161), .B(n_216), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_228), .A2(n_199), .B1(n_215), .B2(n_216), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_258), .B(n_215), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_246), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_247), .A2(n_212), .B(n_202), .C(n_198), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_243), .B(n_182), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_229), .A2(n_182), .B1(n_167), .B2(n_166), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_229), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_258), .B(n_182), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_249), .Y(n_297) );
AOI33xp33_ASAP7_75t_L g298 ( .A1(n_222), .A2(n_170), .A3(n_196), .B1(n_175), .B2(n_182), .B3(n_189), .Y(n_298) );
NOR2xp33_ASAP7_75t_R g299 ( .A(n_276), .B(n_54), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_234), .A2(n_170), .B1(n_196), .B2(n_175), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_234), .B(n_263), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
AO21x1_ASAP7_75t_L g303 ( .A1(n_233), .A2(n_208), .B(n_189), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_234), .A2(n_208), .B1(n_189), .B2(n_211), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_235), .A2(n_208), .B1(n_189), .B2(n_211), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_218), .B(n_221), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_273), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_250), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_SL g309 ( .A1(n_278), .A2(n_208), .B(n_60), .C(n_64), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_225), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_269), .A2(n_55), .B(n_67), .C(n_71), .Y(n_312) );
AO32x1_ASAP7_75t_L g313 ( .A1(n_262), .A2(n_211), .A3(n_267), .B1(n_265), .B2(n_272), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_235), .B(n_211), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_218), .B(n_219), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_226), .B(n_230), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_240), .A2(n_239), .B(n_253), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_263), .B(n_277), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_226), .B(n_245), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_268), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_268), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g322 ( .A1(n_251), .A2(n_257), .B1(n_232), .B2(n_273), .C1(n_263), .C2(n_256), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_263), .B(n_264), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_271), .A2(n_275), .B(n_224), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_248), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_311), .A2(n_256), .B1(n_240), .B2(n_242), .Y(n_327) );
AO31x2_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_252), .A3(n_259), .B(n_260), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_280), .B(n_236), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_285), .A2(n_224), .B(n_227), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_292), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_299), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_285), .A2(n_227), .B(n_266), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_316), .A2(n_220), .B(n_244), .C(n_261), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_299), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_306), .A2(n_254), .B(n_274), .C(n_268), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_302), .B(n_268), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_290), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_324), .A2(n_323), .B(n_287), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_294), .B(n_315), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_319), .A2(n_286), .B1(n_282), .B2(n_284), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_289), .A2(n_288), .B(n_281), .C(n_318), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_313), .A2(n_291), .B(n_318), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_292), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g345 ( .A1(n_325), .A2(n_322), .B(n_309), .C(n_295), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_283), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_296), .B(n_301), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_323), .A2(n_317), .B(n_313), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_313), .A2(n_309), .B(n_304), .Y(n_349) );
CKINVDCx6p67_ASAP7_75t_R g350 ( .A(n_314), .Y(n_350) );
AO32x2_ASAP7_75t_L g351 ( .A1(n_313), .A2(n_298), .A3(n_300), .B1(n_312), .B2(n_279), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_308), .A2(n_298), .B(n_293), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_320), .A2(n_321), .B(n_301), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_307), .B(n_310), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_330), .A2(n_314), .B(n_305), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_330), .A2(n_293), .B(n_307), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_326), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_340), .B(n_338), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_353), .Y(n_360) );
NOR2x1_ASAP7_75t_SL g361 ( .A(n_344), .B(n_341), .Y(n_361) );
INVx4_ASAP7_75t_L g362 ( .A(n_344), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_354), .B(n_346), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_342), .A2(n_333), .B(n_352), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_352), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_349), .A2(n_343), .B(n_333), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_329), .B(n_332), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_341), .A2(n_329), .B1(n_345), .B2(n_335), .C(n_327), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_334), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_337), .B(n_331), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_331), .B(n_350), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_345), .A2(n_343), .B(n_349), .C(n_336), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_344), .B(n_347), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_347), .B(n_351), .Y(n_374) );
OAI22xp5_ASAP7_75t_SL g375 ( .A1(n_348), .A2(n_311), .B1(n_128), .B2(n_225), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_328), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_328), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_351), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_358), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_375), .A2(n_351), .B1(n_368), .B2(n_363), .C(n_359), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_376), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_376), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_362), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_359), .B(n_358), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_378), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_372), .A2(n_356), .B(n_364), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_362), .B(n_361), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_370), .B(n_365), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_378), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_362), .B(n_365), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_375), .A2(n_367), .B1(n_357), .B2(n_379), .C(n_378), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_355), .A2(n_360), .B(n_379), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_355), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_377), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_374), .B(n_370), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_377), .Y(n_400) );
AO21x2_ASAP7_75t_L g401 ( .A1(n_369), .A2(n_360), .B(n_380), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_373), .B(n_379), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_374), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_371), .B(n_380), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_380), .B(n_366), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_371), .B(n_366), .Y(n_407) );
OA21x2_ASAP7_75t_L g408 ( .A1(n_360), .A2(n_369), .B(n_366), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_359), .B(n_370), .Y(n_412) );
NOR2x1_ASAP7_75t_SL g413 ( .A(n_362), .B(n_344), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_362), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_407), .B(n_399), .Y(n_415) );
INVx5_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_407), .B(n_399), .Y(n_417) );
BUFx8_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_404), .B(n_393), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_404), .B(n_393), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_385), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_405), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_383), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_412), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_385), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_381), .B(n_392), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_392), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_385), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_382), .A2(n_394), .B1(n_412), .B2(n_386), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_397), .B(n_402), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_402), .B(n_384), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_411), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_391), .B(n_414), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_391), .B(n_389), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_414), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_414), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_403), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_406), .B(n_400), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_387), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_414), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_406), .B(n_400), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_387), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_403), .B(n_409), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_408), .B(n_409), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_396), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_390), .B(n_410), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_410), .B(n_409), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_401), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_409), .B(n_408), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_415), .B(n_409), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_418), .B(n_410), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_432), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_432), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_430), .B(n_413), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_415), .B(n_408), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
NAND2xp33_ASAP7_75t_R g471 ( .A(n_421), .B(n_408), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_417), .B(n_401), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_417), .B(n_401), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_440), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_396), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_421), .B(n_395), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_419), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_423), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_423), .B(n_395), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_426), .B(n_413), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_422), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_442), .B(n_441), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g484 ( .A(n_416), .B(n_428), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_451), .B(n_441), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_426), .B(n_439), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_439), .B(n_442), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_451), .B(n_446), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_445), .B(n_446), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_420), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_456), .B(n_462), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_420), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_429), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_418), .B(n_433), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_418), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_429), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_433), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_459), .A2(n_434), .B1(n_421), .B2(n_436), .Y(n_498) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_437), .B(n_436), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_450), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_434), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_456), .B(n_462), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_459), .B(n_434), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_459), .B(n_434), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_454), .B(n_428), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_416), .B(n_431), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_416), .B(n_437), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_459), .B(n_436), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_436), .B(n_450), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_454), .B(n_422), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_422), .B(n_424), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_460), .B(n_416), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_449), .A2(n_447), .B1(n_431), .B2(n_425), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_443), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_416), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_424), .B(n_438), .Y(n_516) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_437), .B(n_447), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_485), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_486), .B(n_435), .Y(n_519) );
INVxp67_ASAP7_75t_SL g520 ( .A(n_484), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_512), .B(n_460), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_471), .B(n_461), .C(n_457), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_515), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_485), .B(n_457), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_487), .B(n_435), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_469), .B(n_460), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_464), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_478), .B(n_435), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_469), .B(n_460), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_464), .B(n_460), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_479), .B(n_427), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_515), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_491), .B(n_424), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_488), .B(n_427), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_505), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_515), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_488), .B(n_427), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_466), .B(n_438), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_491), .B(n_438), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_490), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_467), .B(n_452), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_502), .B(n_443), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_502), .B(n_444), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_470), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_473), .B(n_444), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_505), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_473), .B(n_444), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_483), .B(n_452), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_482), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_470), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_512), .B(n_416), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_492), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_483), .B(n_448), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
OAI21xp33_ASAP7_75t_L g555 ( .A1(n_489), .A2(n_461), .B(n_425), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_474), .B(n_455), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_493), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_474), .B(n_455), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_476), .B(n_455), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_480), .B(n_458), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
BUFx3_ASAP7_75t_L g563 ( .A(n_495), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_480), .B(n_458), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_482), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_497), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_524), .B(n_510), .Y(n_568) );
AOI32xp33_ASAP7_75t_L g569 ( .A1(n_544), .A2(n_494), .A3(n_465), .B1(n_503), .B2(n_504), .Y(n_569) );
CKINVDCx16_ASAP7_75t_R g570 ( .A(n_563), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_535), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_554), .A2(n_481), .B1(n_468), .B2(n_508), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_546), .B(n_510), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_524), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_518), .B(n_509), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_561), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_563), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_540), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_503), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_552), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_519), .B(n_509), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_525), .B(n_475), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_547), .B(n_472), .Y(n_583) );
AOI211xp5_ASAP7_75t_SL g584 ( .A1(n_520), .A2(n_512), .B(n_501), .C(n_463), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_549), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_557), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_547), .B(n_511), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_522), .A2(n_498), .B(n_504), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_550), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_562), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_566), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_560), .B(n_516), .Y(n_592) );
NOR2xp67_ASAP7_75t_L g593 ( .A(n_550), .B(n_465), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_567), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_560), .B(n_516), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_549), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_564), .B(n_511), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_523), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_551), .A2(n_507), .B1(n_499), .B2(n_501), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_553), .B(n_501), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_564), .B(n_508), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_548), .B(n_514), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_570), .B(n_551), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_600), .A2(n_588), .B1(n_572), .B2(n_593), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_576), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_584), .A2(n_506), .B(n_555), .Y(n_606) );
XOR2x2_ASAP7_75t_L g607 ( .A(n_576), .B(n_551), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_569), .A2(n_521), .B(n_536), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_571), .B(n_536), .C(n_532), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_574), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_578), .A2(n_529), .B1(n_526), .B2(n_586), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_577), .A2(n_536), .B(n_523), .C(n_532), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_589), .B(n_529), .Y(n_613) );
AOI31xp33_ASAP7_75t_L g614 ( .A1(n_599), .A2(n_507), .A3(n_521), .B(n_526), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_580), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_590), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_585), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_591), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_594), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_579), .B(n_543), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_568), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_587), .B(n_556), .Y(n_622) );
OAI321xp33_ASAP7_75t_L g623 ( .A1(n_598), .A2(n_541), .A3(n_530), .B1(n_537), .B2(n_534), .C(n_531), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_607), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_604), .B(n_598), .Y(n_625) );
OAI31xp33_ASAP7_75t_L g626 ( .A1(n_608), .A2(n_612), .A3(n_603), .B(n_609), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_614), .A2(n_573), .B1(n_600), .B2(n_521), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_606), .A2(n_506), .B(n_517), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_623), .A2(n_601), .B(n_575), .C(n_597), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_615), .Y(n_630) );
AOI21xp33_ASAP7_75t_SL g631 ( .A1(n_609), .A2(n_602), .B(n_534), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_606), .A2(n_582), .B(n_583), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_605), .B(n_596), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_610), .B(n_581), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_616), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_611), .A2(n_537), .B(n_595), .Y(n_636) );
NOR2xp33_ASAP7_75t_R g637 ( .A(n_624), .B(n_621), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_626), .B(n_611), .C(n_619), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g639 ( .A1(n_625), .A2(n_618), .B(n_613), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g640 ( .A(n_628), .B(n_622), .C(n_513), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_625), .A2(n_530), .B1(n_617), .B2(n_620), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_627), .A2(n_543), .B1(n_542), .B2(n_539), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_636), .A2(n_556), .B(n_545), .C(n_558), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_638), .B(n_631), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g645 ( .A1(n_642), .A2(n_629), .B(n_632), .C(n_633), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g646 ( .A(n_637), .B(n_635), .C(n_630), .Y(n_646) );
NOR3xp33_ASAP7_75t_SL g647 ( .A(n_640), .B(n_634), .C(n_528), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_647), .B(n_641), .Y(n_648) );
NAND4xp75_ASAP7_75t_L g649 ( .A(n_644), .B(n_639), .C(n_643), .D(n_542), .Y(n_649) );
NAND3xp33_ASAP7_75t_SL g650 ( .A(n_646), .B(n_592), .C(n_596), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_649), .A2(n_645), .B1(n_545), .B2(n_559), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g652 ( .A(n_648), .B(n_533), .Y(n_652) );
XNOR2xp5_ASAP7_75t_L g653 ( .A(n_652), .B(n_650), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_651), .B1(n_585), .B2(n_463), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_538), .B(n_453), .Y(n_655) );
OR2x6_ASAP7_75t_L g656 ( .A(n_655), .B(n_453), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_416), .B1(n_463), .B2(n_565), .C(n_533), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_477), .B1(n_539), .B2(n_565), .Y(n_658) );
endmodule