module fake_jpeg_11492_n_576 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_576);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_576;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_2),
.B(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_2),
.B(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_65),
.Y(n_186)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_66),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_67),
.Y(n_195)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_22),
.B(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_70),
.B(n_71),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_22),
.B(n_9),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_74),
.B(n_78),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_9),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_80),
.Y(n_150)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_32),
.B1(n_25),
.B2(n_26),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_84),
.A2(n_44),
.B1(n_54),
.B2(n_39),
.Y(n_192)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_88),
.Y(n_204)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_90),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_91),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_92),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_37),
.B(n_11),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_104),
.B(n_115),
.Y(n_181)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_107),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_111),
.Y(n_166)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_19),
.B(n_11),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_47),
.Y(n_116)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_117),
.B(n_120),
.Y(n_188)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_19),
.B(n_17),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_122),
.B(n_123),
.Y(n_199)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_49),
.B(n_31),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_124),
.B(n_45),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_59),
.B1(n_47),
.B2(n_40),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_129),
.A2(n_144),
.B1(n_202),
.B2(n_54),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_141),
.B(n_145),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_94),
.B1(n_59),
.B2(n_47),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_151),
.B(n_176),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_96),
.A2(n_40),
.B1(n_44),
.B2(n_59),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_152),
.A2(n_169),
.B1(n_192),
.B2(n_193),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_84),
.A2(n_44),
.B1(n_28),
.B2(n_53),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_27),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_65),
.Y(n_177)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_80),
.Y(n_180)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_103),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_183),
.B(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_62),
.Y(n_189)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_190),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_93),
.A2(n_56),
.B1(n_60),
.B2(n_29),
.Y(n_193)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_67),
.Y(n_197)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_198),
.B(n_38),
.Y(n_252)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_117),
.A2(n_54),
.B1(n_45),
.B2(n_60),
.Y(n_202)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_206),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_207),
.B(n_230),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_99),
.B1(n_97),
.B2(n_102),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_208),
.A2(n_215),
.B1(n_191),
.B2(n_150),
.Y(n_281)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_209),
.Y(n_305)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_210),
.Y(n_306)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_212),
.Y(n_280)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_213),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_194),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_214),
.B(n_223),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_125),
.B1(n_109),
.B2(n_101),
.Y(n_215)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_56),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_220),
.B(n_272),
.Y(n_282)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

OAI22x1_ASAP7_75t_L g313 ( 
.A1(n_222),
.A2(n_255),
.B1(n_268),
.B2(n_196),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_117),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_224),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_148),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_225),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_54),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_226),
.A2(n_239),
.B(n_265),
.Y(n_310)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_149),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_231),
.B(n_237),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_198),
.A2(n_90),
.B1(n_88),
.B2(n_77),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_233),
.A2(n_243),
.B1(n_247),
.B2(n_196),
.Y(n_312)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_181),
.A2(n_75),
.A3(n_92),
.B1(n_91),
.B2(n_30),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g292 ( 
.A1(n_234),
.A2(n_259),
.A3(n_130),
.B1(n_36),
.B2(n_203),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_20),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_235),
.B(n_236),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_20),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_194),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_136),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_132),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_240),
.B(n_246),
.Y(n_300)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_199),
.A2(n_166),
.B(n_130),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_244),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_129),
.A2(n_24),
.B1(n_53),
.B2(n_51),
.Y(n_247)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_249),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_250),
.Y(n_329)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_251),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_252),
.B(n_254),
.Y(n_302)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_171),
.B(n_168),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_164),
.A2(n_54),
.B1(n_51),
.B2(n_50),
.Y(n_255)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_170),
.B(n_50),
.CI(n_42),
.CON(n_259),
.SN(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_159),
.Y(n_260)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_139),
.B(n_36),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_269),
.C(n_273),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_144),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_262),
.B(n_264),
.Y(n_325)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_143),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_137),
.B(n_0),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_158),
.Y(n_267)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_164),
.A2(n_42),
.B1(n_38),
.B2(n_33),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_138),
.B(n_1),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_150),
.Y(n_270)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

BUFx4f_ASAP7_75t_SL g271 ( 
.A(n_155),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_157),
.B(n_27),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_161),
.B(n_1),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g274 ( 
.A(n_127),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_275),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_126),
.B(n_31),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_133),
.B(n_24),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_276),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_205),
.B1(n_204),
.B2(n_163),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_278),
.A2(n_281),
.B1(n_323),
.B2(n_326),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_232),
.A2(n_165),
.B1(n_160),
.B2(n_182),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_284),
.A2(n_286),
.B1(n_292),
.B2(n_313),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_259),
.A2(n_191),
.B1(n_153),
.B2(n_186),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_175),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_318),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_246),
.A2(n_131),
.B1(n_140),
.B2(n_135),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

NAND2x1_ASAP7_75t_SL g299 ( 
.A(n_261),
.B(n_36),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_299),
.A2(n_308),
.B(n_279),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_239),
.B(n_186),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_269),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_250),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_315),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_226),
.A2(n_3),
.B(n_5),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_308),
.A2(n_243),
.B(n_207),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_257),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_250),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_239),
.A2(n_195),
.B1(n_135),
.B2(n_128),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_317),
.A2(n_319),
.B1(n_332),
.B2(n_251),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_220),
.B(n_195),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_234),
.A2(n_128),
.B1(n_5),
.B2(n_6),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_216),
.A2(n_238),
.B1(n_266),
.B2(n_226),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_248),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_228),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_291),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_334),
.B(n_342),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_294),
.A2(n_218),
.B1(n_256),
.B2(n_245),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_336),
.A2(n_352),
.B1(n_360),
.B2(n_367),
.Y(n_380)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_309),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_339),
.B(n_355),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_340),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_288),
.B(n_273),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_341),
.B(n_347),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_265),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_343),
.B(n_351),
.Y(n_395)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_328),
.Y(n_346)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_288),
.B(n_273),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_300),
.A2(n_243),
.B(n_265),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_349),
.A2(n_368),
.B(n_365),
.Y(n_405)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_295),
.Y(n_350)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_301),
.B(n_269),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_312),
.A2(n_292),
.B1(n_278),
.B2(n_279),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_309),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_359),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_354),
.A2(n_363),
.B(n_365),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_271),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_362),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_241),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_311),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_361),
.Y(n_410)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_302),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_310),
.A2(n_218),
.B1(n_210),
.B2(n_258),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_364),
.A2(n_366),
.B1(n_330),
.B2(n_324),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_270),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_299),
.A2(n_263),
.B1(n_244),
.B2(n_260),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_267),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_368),
.A2(n_370),
.B(n_371),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_282),
.B(n_250),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_372),
.C(n_374),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_229),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_315),
.B(n_227),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_303),
.B(n_227),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_311),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_293),
.B1(n_306),
.B2(n_314),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_287),
.B(n_219),
.C(n_271),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_313),
.A2(n_219),
.B1(n_217),
.B2(n_242),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_375),
.A2(n_306),
.B1(n_296),
.B2(n_330),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_338),
.A2(n_289),
.B1(n_277),
.B2(n_305),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_377),
.A2(n_384),
.B1(n_387),
.B2(n_399),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_383),
.A2(n_396),
.B1(n_404),
.B2(n_411),
.Y(n_413)
);

OAI22x1_ASAP7_75t_SL g384 ( 
.A1(n_356),
.A2(n_360),
.B1(n_338),
.B2(n_352),
.Y(n_384)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_356),
.A2(n_305),
.B1(n_289),
.B2(n_307),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_354),
.A2(n_296),
.B(n_277),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_392),
.A2(n_393),
.B(n_349),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_307),
.B(n_331),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_360),
.A2(n_320),
.B1(n_331),
.B2(n_293),
.Y(n_396)
);

OA22x2_ASAP7_75t_L g397 ( 
.A1(n_364),
.A2(n_320),
.B1(n_314),
.B2(n_321),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_335),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_333),
.A2(n_253),
.B1(n_302),
.B2(n_327),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_280),
.C(n_316),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_372),
.C(n_374),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_333),
.A2(n_206),
.B1(n_209),
.B2(n_321),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_402),
.A2(n_408),
.B1(n_409),
.B2(n_346),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_366),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_324),
.B1(n_283),
.B2(n_285),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_405),
.A2(n_368),
.B(n_365),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_359),
.A2(n_283),
.B1(n_285),
.B2(n_329),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_342),
.A2(n_329),
.B1(n_211),
.B2(n_213),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_336),
.A2(n_221),
.B1(n_249),
.B2(n_297),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_377),
.A2(n_344),
.B1(n_339),
.B2(n_353),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_412),
.A2(n_434),
.B1(n_411),
.B2(n_396),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_415),
.B(n_416),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_423),
.C(n_424),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_430),
.B1(n_432),
.B2(n_438),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_390),
.B(n_334),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_433),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_385),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_429),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_358),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_351),
.C(n_374),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_343),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_407),
.C(n_390),
.Y(n_456)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_426),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_370),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_427),
.Y(n_444)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_428),
.Y(n_466)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_380),
.A2(n_371),
.B1(n_341),
.B2(n_347),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_392),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_431),
.B(n_435),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_380),
.A2(n_384),
.B1(n_398),
.B2(n_405),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_337),
.B1(n_361),
.B2(n_357),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_373),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_381),
.A2(n_345),
.B(n_348),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_407),
.Y(n_450)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_437),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_393),
.A2(n_350),
.B1(n_297),
.B2(n_274),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_439),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_395),
.B(n_297),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_440),
.B(n_399),
.Y(n_451)
);

CKINVDCx6p67_ASAP7_75t_R g441 ( 
.A(n_383),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_441),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_442),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_400),
.C(n_401),
.Y(n_443)
);

A2O1A1O1Ixp25_ASAP7_75t_L g475 ( 
.A1(n_443),
.A2(n_415),
.B(n_430),
.C(n_435),
.D(n_412),
.Y(n_475)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_450),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_451),
.B(n_470),
.Y(n_491)
);

HB1xp67_ASAP7_75t_SL g452 ( 
.A(n_416),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_452),
.A2(n_454),
.B1(n_432),
.B2(n_431),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_421),
.A2(n_406),
.B1(n_404),
.B2(n_410),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_453),
.A2(n_463),
.B1(n_418),
.B2(n_422),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_460),
.C(n_465),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_401),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_434),
.A2(n_387),
.B1(n_410),
.B2(n_388),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_414),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_426),
.B1(n_441),
.B2(n_382),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_402),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_382),
.C(n_391),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_467),
.B(n_442),
.C(n_436),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_418),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_468),
.B(n_389),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_440),
.B(n_388),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_482),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_473),
.A2(n_474),
.B1(n_484),
.B2(n_492),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_477),
.Y(n_497)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_457),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_421),
.C(n_429),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_481),
.Y(n_505)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_406),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_480),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_428),
.C(n_433),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_437),
.C(n_420),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_462),
.A2(n_438),
.B1(n_439),
.B2(n_420),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_485),
.Y(n_506)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_486),
.Y(n_510)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_458),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_488),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_443),
.C(n_456),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_494),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_445),
.A2(n_441),
.B1(n_413),
.B2(n_391),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_493),
.B1(n_453),
.B2(n_454),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_461),
.A2(n_441),
.B1(n_403),
.B2(n_408),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_445),
.A2(n_386),
.B1(n_397),
.B2(n_389),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_469),
.C(n_451),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_495),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_450),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_499),
.B(n_501),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_469),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_504),
.A2(n_473),
.B1(n_484),
.B2(n_459),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_479),
.Y(n_507)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_507),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_469),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_515),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_470),
.Y(n_515)
);

NOR2x1p5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_474),
.Y(n_517)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_517),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_481),
.C(n_489),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_518),
.B(n_520),
.C(n_529),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_519),
.A2(n_468),
.B1(n_448),
.B2(n_497),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_482),
.C(n_483),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_444),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_525),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_459),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_523),
.B(n_524),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_511),
.B(n_455),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_506),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_498),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_528),
.Y(n_538)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_513),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_496),
.B(n_483),
.C(n_455),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_509),
.A2(n_490),
.B1(n_463),
.B2(n_493),
.Y(n_531)
);

OAI321xp33_ASAP7_75t_L g535 ( 
.A1(n_531),
.A2(n_502),
.A3(n_503),
.B1(n_514),
.B2(n_475),
.C(n_498),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_532),
.A2(n_544),
.B1(n_397),
.B2(n_297),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_530),
.B(n_501),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_540),
.C(n_529),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_496),
.C(n_513),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_536),
.Y(n_547)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_535),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_499),
.C(n_512),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_515),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_527),
.B(n_507),
.C(n_448),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_491),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_521),
.A2(n_492),
.B1(n_447),
.B2(n_378),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g545 ( 
.A(n_543),
.B(n_516),
.C(n_520),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_545),
.B(n_549),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_539),
.A2(n_517),
.B1(n_447),
.B2(n_378),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_546),
.A2(n_551),
.B(n_554),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_552),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_541),
.Y(n_549)
);

NAND4xp25_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_517),
.C(n_397),
.D(n_491),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_544),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_534),
.A2(n_397),
.B(n_274),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_550),
.B(n_537),
.Y(n_555)
);

OAI21x1_ASAP7_75t_SL g567 ( 
.A1(n_555),
.A2(n_557),
.B(n_562),
.Y(n_567)
);

BUFx4f_ASAP7_75t_SL g557 ( 
.A(n_549),
.Y(n_557)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_558),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_538),
.C(n_536),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_560),
.B(n_548),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_SL g562 ( 
.A1(n_546),
.A2(n_533),
.B(n_540),
.C(n_13),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_563),
.A2(n_564),
.B(n_561),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_556),
.A2(n_8),
.B(n_12),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_559),
.B(n_8),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_566),
.B(n_555),
.Y(n_568)
);

AOI31xp33_ASAP7_75t_L g572 ( 
.A1(n_568),
.A2(n_13),
.A3(n_16),
.B(n_17),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_569),
.A2(n_570),
.B(n_567),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_557),
.C(n_14),
.Y(n_570)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_571),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_572),
.B(n_16),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_16),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_17),
.Y(n_576)
);


endmodule