module fake_netlist_5_2551_n_1028 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1028);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1028;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_1024;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_918;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_795;
wire n_857;
wire n_695;
wire n_832;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_86),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_100),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_159),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_22),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_181),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_111),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_157),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_164),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_177),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_73),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_76),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_119),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_172),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_14),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_112),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_28),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_77),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_89),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_54),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_1),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_116),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_195),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_90),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_148),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_96),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_142),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_198),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_211),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_104),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_162),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_7),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_205),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_45),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_126),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_179),
.Y(n_270)
);

BUFx6f_ASAP7_75t_SL g271 ( 
.A(n_27),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_138),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_117),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_82),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_83),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_32),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_135),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_169),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_184),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_66),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_93),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_128),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_113),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_204),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_161),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_178),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_194),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_95),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_64),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_136),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_15),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_67),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_40),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_68),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_170),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_152),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_133),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_109),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_108),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_7),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_188),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_118),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_53),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_18),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_102),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_92),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_140),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_201),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_39),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_151),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_51),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_223),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_253),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_237),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_221),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_240),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_249),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_293),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_0),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_226),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_227),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_292),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_232),
.B(n_1),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_232),
.B(n_2),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_228),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_225),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_244),
.B(n_2),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_229),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_244),
.B(n_3),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_300),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_220),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_222),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_3),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_233),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_237),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_234),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_241),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_230),
.B(n_4),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_235),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_238),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_243),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_248),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_236),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_254),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_256),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_297),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_309),
.B(n_4),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_239),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_225),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_258),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_304),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_246),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_225),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_269),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_272),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_274),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_275),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_242),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_247),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_342),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_318),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_328),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_329),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_334),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_278),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_317),
.B(n_246),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_316),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_279),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_319),
.B(n_282),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_354),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_361),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_360),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_342),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_R g402 ( 
.A(n_370),
.B(n_371),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_324),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_316),
.B(n_284),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_R g408 ( 
.A(n_349),
.B(n_257),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_314),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_343),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_320),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_343),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_345),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_330),
.B(n_286),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_345),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_331),
.B(n_339),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_321),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_357),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_357),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_325),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

INVx8_ASAP7_75t_L g435 ( 
.A(n_412),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_390),
.A2(n_336),
.B1(n_338),
.B2(n_359),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_412),
.B(n_241),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_341),
.B1(n_321),
.B2(n_364),
.Y(n_441)
);

NAND3x1_ASAP7_75t_L g442 ( 
.A(n_383),
.B(n_332),
.C(n_344),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_372),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_398),
.A2(n_374),
.B1(n_376),
.B2(n_373),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_386),
.Y(n_447)
);

INVx6_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_391),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_373),
.B(n_358),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_287),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_401),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

NAND3x1_ASAP7_75t_L g460 ( 
.A(n_394),
.B(n_294),
.C(n_289),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_412),
.B(n_252),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_385),
.B(n_291),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_395),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_406),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_387),
.B(n_364),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_400),
.A2(n_315),
.B1(n_363),
.B2(n_341),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_401),
.B(n_225),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_409),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_392),
.B(n_266),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_395),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_392),
.B(n_308),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_387),
.B(n_315),
.Y(n_475)
);

INVx8_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_409),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_392),
.B(n_241),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_402),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_386),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_413),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_390),
.B(n_259),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_410),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_419),
.A2(n_301),
.B(n_231),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_380),
.B(n_260),
.Y(n_490)
);

INVx8_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

INVx6_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_421),
.B(n_241),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_379),
.B(n_261),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_421),
.B(n_245),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_411),
.A2(n_245),
.B1(n_250),
.B2(n_271),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_380),
.B(n_262),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_411),
.B(n_263),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_388),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_411),
.B(n_265),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_426),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_374),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_469),
.B(n_376),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_450),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_461),
.B(n_378),
.Y(n_509)
);

AND2x6_ASAP7_75t_SL g510 ( 
.A(n_475),
.B(n_426),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_433),
.B(n_505),
.Y(n_512)
);

INVx8_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_436),
.A2(n_225),
.B1(n_231),
.B2(n_245),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_469),
.B(n_378),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_472),
.B(n_396),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_472),
.A2(n_225),
.B1(n_231),
.B2(n_245),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_396),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_476),
.B(n_375),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_459),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_505),
.B(n_403),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_464),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_397),
.Y(n_524)
);

NOR2x1_ASAP7_75t_L g525 ( 
.A(n_452),
.B(n_415),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_476),
.B(n_375),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_476),
.B(n_380),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_481),
.B(n_405),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_488),
.A2(n_231),
.B1(n_250),
.B2(n_429),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_504),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_468),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_462),
.B(n_403),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_501),
.B(n_415),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_488),
.A2(n_231),
.B1(n_250),
.B2(n_429),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_486),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_491),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_479),
.A2(n_231),
.B1(n_250),
.B2(n_422),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_486),
.B(n_268),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_432),
.B(n_416),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_448),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_504),
.B(n_416),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_434),
.B(n_418),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_442),
.A2(n_363),
.B1(n_270),
.B2(n_273),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_444),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_435),
.B(n_277),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_487),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_478),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_482),
.B(n_425),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_479),
.A2(n_418),
.B1(n_422),
.B2(n_255),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_440),
.B(n_280),
.Y(n_550)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_484),
.A2(n_303),
.B(n_281),
.C(n_299),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_435),
.B(n_388),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_448),
.A2(n_255),
.B1(n_267),
.B2(n_307),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_435),
.B(n_388),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_435),
.B(n_283),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_443),
.B(n_449),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_457),
.Y(n_558)
);

NAND2x1_ASAP7_75t_L g559 ( 
.A(n_448),
.B(n_43),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_485),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_442),
.A2(n_492),
.B1(n_482),
.B2(n_496),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_502),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_494),
.B(n_285),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_494),
.B(n_454),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_466),
.B(n_425),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g567 ( 
.A(n_446),
.B(n_441),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_494),
.B(n_288),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_457),
.B(n_410),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_454),
.A2(n_311),
.B(n_290),
.C(n_296),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_492),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_L g572 ( 
.A(n_465),
.B(n_417),
.C(n_414),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_454),
.B(n_438),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_491),
.B(n_298),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_451),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_498),
.B(n_302),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_451),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_445),
.B(n_414),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_438),
.A2(n_267),
.B1(n_312),
.B2(n_420),
.Y(n_580)
);

A2O1A1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_491),
.A2(n_428),
.B(n_427),
.C(n_420),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_490),
.B(n_44),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_500),
.B(n_47),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_460),
.B(n_417),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_460),
.A2(n_428),
.B1(n_427),
.B2(n_97),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_431),
.B(n_48),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_497),
.A2(n_471),
.B1(n_473),
.B2(n_495),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_431),
.B(n_49),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_497),
.B(n_5),
.Y(n_589)
);

NAND2x1_ASAP7_75t_L g590 ( 
.A(n_483),
.B(n_50),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_453),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_508),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_R g593 ( 
.A(n_546),
.B(n_487),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_511),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_530),
.B(n_453),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_520),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_548),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_535),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_514),
.A2(n_471),
.B1(n_480),
.B2(n_495),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_569),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_515),
.B(n_463),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_536),
.B(n_514),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_516),
.B(n_431),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_544),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_506),
.B(n_463),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_512),
.B(n_470),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_557),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_509),
.B(n_470),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_532),
.B(n_467),
.C(n_473),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_512),
.B(n_532),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_533),
.A2(n_480),
.B(n_439),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_561),
.B(n_439),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_564),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_571),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_571),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_510),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

AO22x1_ASAP7_75t_L g621 ( 
.A1(n_524),
.A2(n_499),
.B1(n_503),
.B2(n_489),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_541),
.B(n_483),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_536),
.B(n_574),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_518),
.B(n_483),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_578),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_553),
.A2(n_467),
.B1(n_499),
.B2(n_489),
.C(n_503),
.Y(n_626)
);

BUFx4f_ASAP7_75t_L g627 ( 
.A(n_536),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_558),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_517),
.A2(n_439),
.B1(n_503),
.B2(n_489),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_566),
.B(n_447),
.Y(n_630)
);

AO22x1_ASAP7_75t_L g631 ( 
.A1(n_524),
.A2(n_493),
.B1(n_477),
.B2(n_447),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_579),
.Y(n_632)
);

NOR2x1_ASAP7_75t_R g633 ( 
.A(n_507),
.B(n_456),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_522),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_525),
.B(n_477),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_591),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_531),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_518),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_547),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_560),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_SL g641 ( 
.A(n_521),
.B(n_6),
.C(n_8),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_556),
.B(n_493),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_556),
.B(n_456),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_562),
.B(n_52),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_539),
.B(n_456),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_540),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_521),
.B(n_456),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_567),
.Y(n_649)
);

BUFx12f_ASAP7_75t_L g650 ( 
.A(n_565),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_589),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_651)
);

BUFx4f_ASAP7_75t_L g652 ( 
.A(n_513),
.Y(n_652)
);

NAND2x1p5_ASAP7_75t_L g653 ( 
.A(n_573),
.B(n_590),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_587),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_559),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_539),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_513),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_542),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_653),
.A2(n_527),
.B(n_586),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_658),
.B(n_656),
.Y(n_660)
);

AO32x2_ASAP7_75t_L g661 ( 
.A1(n_629),
.A2(n_616),
.A3(n_599),
.B1(n_631),
.B2(n_604),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_594),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_598),
.B(n_528),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_612),
.A2(n_580),
.B1(n_573),
.B2(n_517),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_593),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_631),
.A2(n_554),
.B(n_552),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_592),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_604),
.A2(n_526),
.B(n_519),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_614),
.A2(n_575),
.B(n_582),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_615),
.A2(n_534),
.B(n_529),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_594),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_651),
.A2(n_585),
.B(n_580),
.C(n_553),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_597),
.B(n_545),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_612),
.A2(n_543),
.B(n_542),
.C(n_549),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_SL g675 ( 
.A1(n_615),
.A2(n_538),
.B(n_545),
.C(n_623),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_598),
.B(n_572),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_599),
.B(n_581),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_603),
.B(n_550),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_603),
.B(n_605),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_644),
.A2(n_529),
.B1(n_534),
.B2(n_568),
.Y(n_680)
);

OA21x2_ASAP7_75t_L g681 ( 
.A1(n_622),
.A2(n_588),
.B(n_583),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_596),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_653),
.A2(n_555),
.B(n_563),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_607),
.B(n_550),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_632),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_653),
.A2(n_537),
.B(n_549),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_623),
.A2(n_537),
.B(n_577),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_595),
.A2(n_570),
.B(n_458),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_610),
.B(n_551),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_608),
.A2(n_584),
.B(n_458),
.Y(n_690)
);

OAI22x1_ASAP7_75t_L g691 ( 
.A1(n_649),
.A2(n_565),
.B1(n_584),
.B2(n_11),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_632),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_637),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_634),
.Y(n_694)
);

AOI21x1_ASAP7_75t_L g695 ( 
.A1(n_621),
.A2(n_584),
.B(n_458),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_627),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_608),
.A2(n_458),
.B(n_455),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_627),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_600),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_616),
.B(n_565),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_648),
.A2(n_455),
.B1(n_105),
.B2(n_106),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_602),
.B(n_9),
.Y(n_702)
);

BUFx2_ASAP7_75t_R g703 ( 
.A(n_619),
.Y(n_703)
);

AO31x2_ASAP7_75t_L g704 ( 
.A1(n_654),
.A2(n_10),
.A3(n_12),
.B(n_13),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_642),
.A2(n_455),
.B1(n_107),
.B2(n_110),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_639),
.B(n_455),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g707 ( 
.A1(n_654),
.A2(n_99),
.B(n_217),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_597),
.B(n_55),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_640),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_655),
.A2(n_103),
.B(n_215),
.Y(n_710)
);

OAI21xp33_ASAP7_75t_L g711 ( 
.A1(n_641),
.A2(n_12),
.B(n_13),
.Y(n_711)
);

AOI21x1_ASAP7_75t_SL g712 ( 
.A1(n_646),
.A2(n_14),
.B(n_15),
.Y(n_712)
);

AOI21xp33_ASAP7_75t_L g713 ( 
.A1(n_633),
.A2(n_16),
.B(n_17),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_669),
.A2(n_627),
.B(n_597),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_663),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_677),
.B(n_657),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_684),
.B(n_645),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_674),
.A2(n_611),
.B(n_626),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_662),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_659),
.A2(n_655),
.B(n_601),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_696),
.B(n_643),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_670),
.A2(n_638),
.B(n_645),
.C(n_652),
.Y(n_722)
);

AO31x2_ASAP7_75t_L g723 ( 
.A1(n_669),
.A2(n_680),
.A3(n_668),
.B(n_664),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_672),
.A2(n_645),
.B(n_652),
.C(n_606),
.Y(n_724)
);

CKINVDCx6p67_ASAP7_75t_R g725 ( 
.A(n_691),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_683),
.A2(n_606),
.B(n_600),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_678),
.B(n_628),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_696),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_694),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_662),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_671),
.Y(n_731)
);

AO21x2_ASAP7_75t_L g732 ( 
.A1(n_668),
.A2(n_624),
.B(n_609),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_671),
.B(n_609),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_707),
.A2(n_625),
.B(n_613),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_667),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_682),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_660),
.B(n_628),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_698),
.Y(n_738)
);

INVxp67_ASAP7_75t_SL g739 ( 
.A(n_679),
.Y(n_739)
);

AO31x2_ASAP7_75t_L g740 ( 
.A1(n_674),
.A2(n_625),
.A3(n_636),
.B(n_613),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_666),
.A2(n_636),
.B(n_617),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_665),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_693),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_695),
.A2(n_617),
.B(n_618),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_681),
.A2(n_597),
.B(n_652),
.Y(n_745)
);

OAI21xp5_ASAP7_75t_L g746 ( 
.A1(n_675),
.A2(n_630),
.B(n_647),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_672),
.A2(n_689),
.B(n_688),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_710),
.A2(n_617),
.B(n_618),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_709),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_687),
.A2(n_618),
.B(n_620),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_699),
.B(n_630),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_699),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_688),
.A2(n_620),
.B(n_647),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_698),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_L g755 ( 
.A1(n_711),
.A2(n_619),
.B1(n_630),
.B2(n_620),
.C(n_643),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_676),
.A2(n_650),
.B1(n_635),
.B2(n_643),
.Y(n_756)
);

OAI21x1_ASAP7_75t_L g757 ( 
.A1(n_697),
.A2(n_686),
.B(n_690),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_702),
.A2(n_650),
.B1(n_643),
.B2(n_657),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_677),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_712),
.A2(n_635),
.B(n_597),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_SL g761 ( 
.A(n_703),
.B(n_657),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_700),
.A2(n_643),
.B1(n_635),
.B2(n_18),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_685),
.B(n_635),
.Y(n_763)
);

AOI221xp5_ASAP7_75t_L g764 ( 
.A1(n_713),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.C(n_20),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_739),
.B(n_692),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_715),
.B(n_702),
.Y(n_766)
);

AOI221xp5_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_705),
.B1(n_701),
.B2(n_708),
.C(n_706),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_716),
.B(n_708),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_719),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_737),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_717),
.B(n_673),
.Y(n_771)
);

BUFx4f_ASAP7_75t_SL g772 ( 
.A(n_725),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_742),
.Y(n_773)
);

AOI221xp5_ASAP7_75t_L g774 ( 
.A1(n_718),
.A2(n_673),
.B1(n_712),
.B2(n_704),
.C(n_661),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_729),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_SL g776 ( 
.A1(n_722),
.A2(n_661),
.B(n_704),
.C(n_635),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_725),
.A2(n_635),
.B1(n_681),
.B2(n_661),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_761),
.A2(n_681),
.B1(n_661),
.B2(n_704),
.Y(n_778)
);

NAND3xp33_ASAP7_75t_SL g779 ( 
.A(n_722),
.B(n_704),
.C(n_20),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_747),
.A2(n_121),
.B(n_214),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_721),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_717),
.B(n_19),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_727),
.B(n_21),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_724),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_755),
.B(n_735),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_719),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_721),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_724),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_721),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_736),
.Y(n_790)
);

INVx6_ASAP7_75t_L g791 ( 
.A(n_716),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_714),
.A2(n_123),
.B(n_213),
.Y(n_792)
);

OA21x2_ASAP7_75t_L g793 ( 
.A1(n_741),
.A2(n_122),
.B(n_212),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_741),
.A2(n_120),
.B(n_209),
.Y(n_794)
);

OR2x6_ASAP7_75t_L g795 ( 
.A(n_716),
.B(n_56),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_762),
.A2(n_759),
.B1(n_756),
.B2(n_758),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_721),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_751),
.B(n_57),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_743),
.B(n_24),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_749),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_742),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_751),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_728),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_754),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_SL g805 ( 
.A1(n_763),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_805)
);

INVx3_ASAP7_75t_SL g806 ( 
.A(n_721),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_728),
.Y(n_807)
);

CKINVDCx11_ASAP7_75t_R g808 ( 
.A(n_730),
.Y(n_808)
);

AOI221xp5_ASAP7_75t_L g809 ( 
.A1(n_746),
.A2(n_752),
.B1(n_733),
.B2(n_730),
.C(n_731),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_728),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_810)
);

CKINVDCx6p67_ASAP7_75t_R g811 ( 
.A(n_721),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_733),
.B(n_33),
.Y(n_812)
);

NOR2x1_ASAP7_75t_SL g813 ( 
.A(n_732),
.B(n_58),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_738),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_738),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_815)
);

NAND4xp25_ASAP7_75t_L g816 ( 
.A(n_731),
.B(n_36),
.C(n_37),
.D(n_38),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_SL g817 ( 
.A1(n_738),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_745),
.A2(n_41),
.B1(n_42),
.B2(n_59),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_740),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_L g820 ( 
.A1(n_723),
.A2(n_41),
.B1(n_42),
.B2(n_60),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_740),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_732),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_732),
.A2(n_218),
.B(n_69),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_794),
.A2(n_753),
.B(n_726),
.Y(n_824)
);

CKINVDCx10_ASAP7_75t_R g825 ( 
.A(n_772),
.Y(n_825)
);

OAI211xp5_ASAP7_75t_SL g826 ( 
.A1(n_808),
.A2(n_723),
.B(n_740),
.C(n_757),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_780),
.A2(n_757),
.B(n_760),
.C(n_720),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_770),
.B(n_765),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_819),
.B(n_723),
.Y(n_829)
);

OAI221xp5_ASAP7_75t_L g830 ( 
.A1(n_780),
.A2(n_723),
.B1(n_753),
.B2(n_760),
.C(n_748),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_790),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_SL g832 ( 
.A1(n_784),
.A2(n_65),
.B(n_70),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_816),
.A2(n_720),
.B1(n_748),
.B2(n_744),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_784),
.A2(n_750),
.B(n_726),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_768),
.B(n_750),
.Y(n_835)
);

AOI221xp5_ASAP7_75t_L g836 ( 
.A1(n_788),
.A2(n_820),
.B1(n_816),
.B2(n_804),
.C(n_814),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_800),
.Y(n_837)
);

OAI22x1_ASAP7_75t_L g838 ( 
.A1(n_777),
.A2(n_734),
.B1(n_744),
.B2(n_74),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_775),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_821),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_788),
.A2(n_734),
.B1(n_72),
.B2(n_75),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_SL g842 ( 
.A1(n_818),
.A2(n_71),
.B1(n_78),
.B2(n_79),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_796),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_804),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_767),
.A2(n_91),
.B(n_94),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_803),
.A2(n_98),
.B1(n_114),
.B2(n_115),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_776),
.A2(n_124),
.B(n_125),
.Y(n_847)
);

OAI211xp5_ASAP7_75t_L g848 ( 
.A1(n_810),
.A2(n_127),
.B(n_129),
.C(n_130),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_815),
.A2(n_782),
.B1(n_798),
.B2(n_795),
.Y(n_849)
);

OAI221xp5_ASAP7_75t_SL g850 ( 
.A1(n_822),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.C(n_137),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_802),
.B(n_208),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_792),
.A2(n_139),
.B(n_141),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_785),
.A2(n_145),
.B(n_146),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_798),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_823),
.A2(n_155),
.B(n_156),
.Y(n_855)
);

AOI222xp33_ASAP7_75t_L g856 ( 
.A1(n_814),
.A2(n_160),
.B1(n_163),
.B2(n_165),
.C1(n_166),
.C2(n_167),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_769),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_766),
.B(n_171),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_795),
.A2(n_768),
.B1(n_779),
.B2(n_818),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_795),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_860)
);

OAI221xp5_ASAP7_75t_L g861 ( 
.A1(n_799),
.A2(n_180),
.B1(n_182),
.B2(n_185),
.C(n_186),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_786),
.Y(n_862)
);

OAI21xp33_ASAP7_75t_L g863 ( 
.A1(n_817),
.A2(n_187),
.B(n_189),
.Y(n_863)
);

OA21x2_ASAP7_75t_L g864 ( 
.A1(n_774),
.A2(n_190),
.B(n_191),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_821),
.Y(n_865)
);

AO31x2_ASAP7_75t_L g866 ( 
.A1(n_813),
.A2(n_192),
.A3(n_196),
.B(n_197),
.Y(n_866)
);

OAI22xp33_ASAP7_75t_L g867 ( 
.A1(n_801),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_789),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_812),
.B(n_206),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_783),
.A2(n_207),
.B1(n_791),
.B2(n_771),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_807),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_829),
.B(n_793),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_829),
.B(n_778),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_831),
.B(n_809),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_835),
.B(n_789),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_837),
.B(n_793),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_828),
.B(n_805),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_835),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_835),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_840),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_840),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_865),
.B(n_781),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_865),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_834),
.B(n_781),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_864),
.B(n_791),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_857),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_864),
.B(n_797),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_824),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_864),
.B(n_797),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_857),
.Y(n_890)
);

OR2x2_ASAP7_75t_SL g891 ( 
.A(n_871),
.B(n_811),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_862),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_839),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_824),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_839),
.B(n_806),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_862),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_826),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_830),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_838),
.B(n_787),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_827),
.B(n_787),
.Y(n_900)
);

AOI221xp5_ASAP7_75t_SL g901 ( 
.A1(n_836),
.A2(n_863),
.B1(n_845),
.B2(n_847),
.C(n_859),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_888),
.A2(n_855),
.B(n_868),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_901),
.A2(n_832),
.B(n_853),
.Y(n_903)
);

AND3x1_ASAP7_75t_L g904 ( 
.A(n_899),
.B(n_849),
.C(n_858),
.Y(n_904)
);

AOI33xp33_ASAP7_75t_L g905 ( 
.A1(n_897),
.A2(n_842),
.A3(n_844),
.B1(n_841),
.B2(n_843),
.B3(n_867),
.Y(n_905)
);

AOI221xp5_ASAP7_75t_L g906 ( 
.A1(n_898),
.A2(n_850),
.B1(n_861),
.B2(n_838),
.C(n_869),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_879),
.B(n_827),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_886),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_886),
.Y(n_909)
);

INVx3_ASAP7_75t_SL g910 ( 
.A(n_891),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_901),
.B(n_856),
.C(n_848),
.Y(n_911)
);

OAI221xp5_ASAP7_75t_L g912 ( 
.A1(n_898),
.A2(n_870),
.B1(n_860),
.B2(n_854),
.C(n_846),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_890),
.Y(n_913)
);

AO21x2_ASAP7_75t_L g914 ( 
.A1(n_888),
.A2(n_833),
.B(n_852),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_880),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_878),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_873),
.A2(n_851),
.B1(n_787),
.B2(n_868),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_SL g918 ( 
.A(n_877),
.B(n_773),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_898),
.A2(n_869),
.B1(n_851),
.B2(n_868),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_899),
.A2(n_825),
.B1(n_866),
.B2(n_897),
.Y(n_920)
);

AO21x2_ASAP7_75t_L g921 ( 
.A1(n_888),
.A2(n_866),
.B(n_894),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_915),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_908),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_916),
.B(n_878),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_908),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_916),
.B(n_878),
.Y(n_926)
);

AND2x4_ASAP7_75t_SL g927 ( 
.A(n_907),
.B(n_895),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_909),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_915),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_907),
.B(n_878),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_909),
.Y(n_931)
);

NOR2x1_ASAP7_75t_L g932 ( 
.A(n_913),
.B(n_893),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_915),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_913),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_910),
.B(n_879),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_921),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_927),
.B(n_910),
.Y(n_937)
);

OAI22xp33_ASAP7_75t_L g938 ( 
.A1(n_935),
.A2(n_911),
.B1(n_903),
.B2(n_873),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_930),
.B(n_878),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_932),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_923),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_925),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_924),
.B(n_885),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_934),
.B(n_874),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_929),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_938),
.B(n_944),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_SL g947 ( 
.A(n_944),
.B(n_903),
.C(n_906),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_945),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_941),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_942),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_940),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_937),
.B(n_927),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_938),
.B(n_918),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_939),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_949),
.Y(n_955)
);

OAI221xp5_ASAP7_75t_SL g956 ( 
.A1(n_946),
.A2(n_904),
.B1(n_911),
.B2(n_920),
.C(n_905),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_954),
.B(n_943),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_953),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_954),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_956),
.A2(n_953),
.B(n_947),
.Y(n_960)
);

OA21x2_ASAP7_75t_SL g961 ( 
.A1(n_958),
.A2(n_930),
.B(n_926),
.Y(n_961)
);

AOI21xp33_ASAP7_75t_L g962 ( 
.A1(n_959),
.A2(n_951),
.B(n_950),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_962),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_961),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_960),
.B(n_959),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_962),
.Y(n_966)
);

NOR4xp25_ASAP7_75t_L g967 ( 
.A(n_965),
.B(n_955),
.C(n_957),
.D(n_948),
.Y(n_967)
);

NAND3xp33_ASAP7_75t_L g968 ( 
.A(n_964),
.B(n_966),
.C(n_963),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_965),
.B(n_957),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_964),
.B(n_948),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_964),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_904),
.C(n_877),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_965),
.Y(n_973)
);

AOI211xp5_ASAP7_75t_L g974 ( 
.A1(n_968),
.A2(n_910),
.B(n_912),
.C(n_952),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_973),
.B(n_895),
.Y(n_975)
);

AOI221xp5_ASAP7_75t_L g976 ( 
.A1(n_971),
.A2(n_936),
.B1(n_934),
.B2(n_914),
.C(n_919),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_972),
.B(n_943),
.C(n_917),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_SL g978 ( 
.A1(n_969),
.A2(n_930),
.B(n_917),
.Y(n_978)
);

NAND4xp25_ASAP7_75t_L g979 ( 
.A(n_970),
.B(n_900),
.C(n_893),
.D(n_924),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_967),
.B(n_891),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_975),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_980),
.B(n_931),
.Y(n_982)
);

OAI311xp33_ASAP7_75t_L g983 ( 
.A1(n_979),
.A2(n_885),
.A3(n_928),
.B1(n_884),
.C1(n_900),
.Y(n_983)
);

OAI21xp33_ASAP7_75t_L g984 ( 
.A1(n_978),
.A2(n_974),
.B(n_977),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_976),
.Y(n_985)
);

NAND2x1_ASAP7_75t_L g986 ( 
.A(n_980),
.B(n_926),
.Y(n_986)
);

AOI221xp5_ASAP7_75t_L g987 ( 
.A1(n_980),
.A2(n_914),
.B1(n_926),
.B2(n_924),
.C(n_874),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_981),
.B(n_893),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_982),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_933),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_985),
.B(n_933),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_986),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_987),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_983),
.B(n_929),
.Y(n_994)
);

NOR2x1p5_ASAP7_75t_L g995 ( 
.A(n_981),
.B(n_878),
.Y(n_995)
);

NAND2x1_ASAP7_75t_L g996 ( 
.A(n_981),
.B(n_900),
.Y(n_996)
);

AOI221xp5_ASAP7_75t_L g997 ( 
.A1(n_985),
.A2(n_914),
.B1(n_872),
.B2(n_922),
.C(n_889),
.Y(n_997)
);

XNOR2xp5_ASAP7_75t_L g998 ( 
.A(n_992),
.B(n_995),
.Y(n_998)
);

AOI211xp5_ASAP7_75t_SL g999 ( 
.A1(n_989),
.A2(n_887),
.B(n_889),
.C(n_922),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_993),
.A2(n_878),
.B1(n_892),
.B2(n_890),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_SL g1001 ( 
.A(n_990),
.B(n_991),
.C(n_997),
.Y(n_1001)
);

XNOR2xp5_ASAP7_75t_L g1002 ( 
.A(n_988),
.B(n_875),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_996),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_994),
.B(n_872),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_SL g1005 ( 
.A(n_994),
.B(n_872),
.C(n_887),
.Y(n_1005)
);

AOI211xp5_ASAP7_75t_L g1006 ( 
.A1(n_992),
.A2(n_884),
.B(n_887),
.C(n_889),
.Y(n_1006)
);

AO22x1_ASAP7_75t_L g1007 ( 
.A1(n_992),
.A2(n_875),
.B1(n_876),
.B2(n_884),
.Y(n_1007)
);

OA22x2_ASAP7_75t_L g1008 ( 
.A1(n_992),
.A2(n_902),
.B1(n_875),
.B2(n_892),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_998),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

AOI211xp5_ASAP7_75t_L g1011 ( 
.A1(n_1000),
.A2(n_902),
.B(n_896),
.C(n_875),
.Y(n_1011)
);

CKINVDCx16_ASAP7_75t_R g1012 ( 
.A(n_1002),
.Y(n_1012)
);

OAI211xp5_ASAP7_75t_L g1013 ( 
.A1(n_1001),
.A2(n_896),
.B(n_894),
.C(n_883),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_1004),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_1012),
.B(n_1005),
.Y(n_1015)
);

XOR2xp5_ASAP7_75t_L g1016 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1014),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_1016),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1017),
.B(n_1013),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_1018),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1019),
.B(n_1015),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_SL g1022 ( 
.A1(n_1021),
.A2(n_1020),
.B(n_1007),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_SL g1023 ( 
.A1(n_1020),
.A2(n_1008),
.B(n_1006),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1022),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1023),
.Y(n_1025)
);

AOI222xp33_ASAP7_75t_L g1026 ( 
.A1(n_1025),
.A2(n_1011),
.B1(n_999),
.B2(n_876),
.C1(n_894),
.C2(n_866),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_1026),
.A2(n_1024),
.B1(n_883),
.B2(n_881),
.C(n_880),
.Y(n_1027)
);

AOI211xp5_ASAP7_75t_L g1028 ( 
.A1(n_1027),
.A2(n_866),
.B(n_882),
.C(n_880),
.Y(n_1028)
);


endmodule