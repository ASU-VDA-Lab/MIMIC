module fake_jpeg_1737_n_55 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_55);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_25),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_15),
.C(n_1),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_17),
.B(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_16),
.B1(n_18),
.B2(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_21),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_20),
.B1(n_18),
.B2(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_27),
.Y(n_36)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_40),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_28),
.C(n_2),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_34),
.C(n_2),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_9),
.B(n_11),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_45),
.C(n_9),
.Y(n_48)
);

A2O1A1O1Ixp25_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_44),
.B(n_11),
.C(n_12),
.D(n_22),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_5),
.C(n_8),
.Y(n_45)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_37),
.CI(n_10),
.CON(n_46),
.SN(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_51),
.B(n_46),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_50),
.B(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_49),
.Y(n_55)
);


endmodule