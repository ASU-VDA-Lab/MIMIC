module real_jpeg_22469_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_11, n_14, n_344, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_11;
input n_14;
input n_344;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_0),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_0),
.A2(n_65),
.B1(n_66),
.B2(n_103),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_103),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_103),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_1),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_2),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_159),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_159),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_159),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_3),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_56),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_265)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_5),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_91),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_91),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_34),
.B1(n_65),
.B2(n_66),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_22),
.B1(n_65),
.B2(n_66),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_7),
.A2(n_22),
.B1(n_48),
.B2(n_49),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_8),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_108),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_108),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_108),
.Y(n_249)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_10),
.B(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_10),
.A2(n_131),
.B(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_12),
.A2(n_49),
.B(n_61),
.C(n_88),
.D(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_12),
.B(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_12),
.B(n_47),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_12),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_12),
.A2(n_109),
.B(n_111),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_12),
.A2(n_31),
.B(n_42),
.C(n_147),
.D(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_12),
.B(n_31),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_12),
.B(n_35),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_32),
.B(n_191),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_127),
.Y(n_207)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_14),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_77),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_75),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_23),
.A2(n_28),
.B(n_127),
.C(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_26),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_26),
.B(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_27),
.A2(n_30),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_27),
.A2(n_30),
.B1(n_218),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_27),
.A2(n_209),
.B(n_249),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_27),
.A2(n_30),
.B1(n_55),
.B2(n_293),
.Y(n_313)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_28),
.Y(n_191)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_30),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_30),
.A2(n_219),
.B(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_46),
.C(n_47),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_35),
.B(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_70),
.C(n_72),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_37),
.A2(n_38),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_53),
.C(n_59),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_39),
.A2(n_40),
.B1(n_59),
.B2(n_318),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_41),
.A2(n_51),
.B1(n_168),
.B2(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_41),
.A2(n_204),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_41),
.A2(n_50),
.B1(n_51),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_47),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_42),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_42),
.A2(n_47),
.B1(n_246),
.B2(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_42),
.A2(n_47),
.B1(n_265),
.B2(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_44),
.B(n_48),
.Y(n_154)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_46),
.Y(n_155)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_62),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_49),
.A2(n_147),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_51),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_51),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_51),
.A2(n_169),
.B(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_53),
.A2(n_54),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_59),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_59),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_68),
.B(n_69),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_60),
.A2(n_68),
.B1(n_102),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_60),
.A2(n_145),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_60),
.A2(n_68),
.B1(n_201),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_60),
.A2(n_68),
.B1(n_231),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_60),
.A2(n_68),
.B1(n_240),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_61),
.A2(n_64),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_66),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_65),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_66),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_68),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_68),
.A2(n_104),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_69),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_70),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_336),
.B(n_342),
.Y(n_77)
);

OAI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_309),
.A3(n_329),
.B1(n_334),
.B2(n_335),
.C(n_344),
.Y(n_78)
);

AOI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_257),
.A3(n_297),
.B1(n_303),
.B2(n_308),
.C(n_345),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_212),
.C(n_253),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_183),
.B(n_211),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_162),
.B(n_182),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_139),
.B(n_161),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_114),
.B(n_138),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_96),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_86),
.B(n_96),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_123),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_89),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_101),
.C(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_109),
.B(n_111),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_113),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_109),
.A2(n_129),
.B1(n_158),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_109),
.A2(n_110),
.B1(n_173),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_109),
.A2(n_194),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_109),
.A2(n_110),
.B1(n_229),
.B2(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_109),
.A2(n_129),
.B(n_238),
.Y(n_270)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_124),
.B(n_137),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_122),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_132),
.B(n_136),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_129),
.Y(n_135)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_141),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_152),
.B2(n_160),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_146),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_151),
.C(n_160),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_164),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_178),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_179),
.C(n_180),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_171),
.B2(n_177),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_174),
.C(n_175),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_185),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_198),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_187),
.B(n_197),
.C(n_198),
.Y(n_254)
);

AOI22x1_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_193),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_195),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_205),
.C(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_213),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_233),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_214),
.B(n_233),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_225),
.C(n_232),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_224),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_232),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_230),
.Y(n_242)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_251),
.B2(n_252),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_241),
.C(n_252),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_239),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_247),
.C(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_255),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_275),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_258),
.B(n_275),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_268),
.C(n_274),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_259),
.A2(n_260),
.B1(n_268),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_270),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_269),
.A2(n_288),
.B(n_292),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_271),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_271),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_295),
.B2(n_296),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_286),
.B2(n_287),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_287),
.C(n_296),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_283),
.B(n_285),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_283),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_284),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_285),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_285),
.A2(n_311),
.B1(n_320),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_294),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_290),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_298),
.A2(n_304),
.B(n_307),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_322),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_322),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_320),
.C(n_321),
.Y(n_310)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_313),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_318),
.C(n_319),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_324),
.C(n_328),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_316),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_332),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_341),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_338),
.Y(n_340)
);


endmodule