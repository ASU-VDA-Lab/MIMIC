module fake_jpeg_9519_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_42),
.B1(n_37),
.B2(n_31),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_81),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_23),
.B1(n_32),
.B2(n_31),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_77),
.B1(n_98),
.B2(n_22),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_74),
.B(n_69),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_23),
.B1(n_27),
.B2(n_20),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_37),
.B(n_45),
.C(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_82),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_45),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_83),
.B(n_84),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_90),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_36),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_39),
.B1(n_38),
.B2(n_40),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_96),
.B1(n_71),
.B2(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_97),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_9),
.C(n_14),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_9),
.B(n_14),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_39),
.B1(n_48),
.B2(n_26),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_22),
.B1(n_30),
.B2(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_103),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_108),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_35),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_124),
.C(n_83),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_65),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_114),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_119),
.B1(n_85),
.B2(n_94),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_145)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_121),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_34),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_66),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_91),
.B1(n_88),
.B2(n_96),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_78),
.B1(n_77),
.B2(n_98),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_78),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_135),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_121),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_132),
.B1(n_144),
.B2(n_147),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_139),
.C(n_143),
.Y(n_185)
);

CKINVDCx12_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_88),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_150),
.B1(n_107),
.B2(n_120),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_145),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_81),
.B(n_99),
.C(n_87),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_102),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_92),
.C(n_88),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_85),
.B1(n_89),
.B2(n_86),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_76),
.B1(n_73),
.B2(n_7),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_100),
.B1(n_122),
.B2(n_84),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_106),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_156),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_106),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_161),
.B1(n_189),
.B2(n_180),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_167),
.B(n_129),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_100),
.B1(n_117),
.B2(n_122),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_173),
.B(n_189),
.Y(n_192)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_115),
.B1(n_117),
.B2(n_127),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_109),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_153),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_108),
.C(n_104),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_178),
.C(n_184),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_175),
.B1(n_181),
.B2(n_182),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_120),
.B1(n_110),
.B2(n_123),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_171),
.B1(n_149),
.B2(n_130),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_146),
.B1(n_142),
.B2(n_152),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_126),
.B1(n_76),
.B2(n_73),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_179),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_79),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_19),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_73),
.B1(n_47),
.B2(n_46),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_47),
.B1(n_46),
.B2(n_19),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_26),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_47),
.C(n_17),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_26),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_133),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_47),
.B1(n_19),
.B2(n_26),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_147),
.B1(n_144),
.B2(n_131),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_34),
.B(n_64),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_153),
.B1(n_145),
.B2(n_150),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_195),
.A2(n_204),
.B(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_169),
.B(n_141),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_196),
.B(n_215),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_198),
.A2(n_181),
.B1(n_164),
.B2(n_184),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_218),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_208),
.Y(n_238)
);

NAND4xp25_ASAP7_75t_SL g203 ( 
.A(n_166),
.B(n_130),
.C(n_131),
.D(n_47),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_168),
.A2(n_135),
.B1(n_35),
.B2(n_17),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_33),
.B1(n_24),
.B2(n_35),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_34),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_191),
.B(n_207),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_163),
.B1(n_165),
.B2(n_170),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_185),
.C(n_178),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_224),
.C(n_233),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_185),
.C(n_162),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_166),
.B1(n_95),
.B2(n_33),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_194),
.B1(n_212),
.B2(n_214),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_190),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_208),
.C(n_192),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_204),
.B(n_11),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_211),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_194),
.A2(n_25),
.B(n_17),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_199),
.A2(n_95),
.B1(n_33),
.B2(n_24),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_33),
.B1(n_24),
.B2(n_25),
.Y(n_261)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

NOR2x1_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_209),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_244),
.B(n_218),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_225),
.B(n_197),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_197),
.C(n_195),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_268),
.C(n_222),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_238),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_95),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_260),
.B(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_266),
.B1(n_220),
.B2(n_246),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_221),
.B(n_13),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_226),
.A2(n_24),
.B1(n_12),
.B2(n_11),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_267),
.B1(n_248),
.B2(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_266)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_0),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_10),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_227),
.B1(n_245),
.B2(n_236),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_283),
.B1(n_256),
.B2(n_264),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_277),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_238),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.C(n_285),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_242),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_242),
.B1(n_228),
.B2(n_223),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_252),
.B(n_268),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_0),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_239),
.C(n_230),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_288),
.B(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_251),
.C(n_228),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_281),
.C(n_282),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_264),
.B(n_267),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_294),
.B(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_296),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_258),
.B(n_243),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_279),
.C(n_2),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_265),
.B1(n_261),
.B2(n_2),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_272),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_10),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_276),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_293),
.C(n_4),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_269),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_306),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_279),
.C(n_3),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_311),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_313),
.B(n_297),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_295),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_0),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_295),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_314),
.B(n_318),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_300),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_305),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_291),
.B1(n_298),
.B2(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_322),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_326),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_312),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_328),
.B(n_329),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_303),
.Y(n_328)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_313),
.B(n_4),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_320),
.B(n_319),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_324),
.B(n_332),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_325),
.Y(n_334)
);

NAND3xp33_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_330),
.C(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_5),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_3),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_3),
.Y(n_338)
);

OAI311xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_4),
.A3(n_5),
.B1(n_329),
.C1(n_333),
.Y(n_339)
);


endmodule