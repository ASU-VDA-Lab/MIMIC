module fake_aes_5898_n_900 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_900);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_900;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_703;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_522;
wire n_883;
wire n_573;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_875;
wire n_339;
wire n_657;
wire n_583;
wire n_728;
wire n_620;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_269;
INVx1_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_218), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_44), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_223), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_219), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_114), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_243), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g274 ( .A(n_214), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_159), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_108), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_26), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_221), .Y(n_278) );
BUFx10_ASAP7_75t_L g279 ( .A(n_239), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_72), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_167), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_30), .Y(n_283) );
CKINVDCx16_ASAP7_75t_R g284 ( .A(n_237), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_46), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_251), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_220), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_196), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_143), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_38), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_235), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_62), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_83), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_232), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_88), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_236), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_193), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_180), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_156), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_226), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_33), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_29), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_231), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_70), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_248), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_99), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_6), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_247), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
INVxp33_ASAP7_75t_SL g311 ( .A(n_254), .Y(n_311) );
BUFx10_ASAP7_75t_L g312 ( .A(n_20), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_182), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_135), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_225), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_0), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_250), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_241), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_191), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_154), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_224), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_213), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_249), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_1), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_169), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_107), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_230), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_211), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_51), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_203), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_119), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_106), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_151), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_160), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_222), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_246), .Y(n_338) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_204), .Y(n_339) );
BUFx10_ASAP7_75t_L g340 ( .A(n_229), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_207), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_54), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_59), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_102), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_227), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_56), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_147), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_215), .Y(n_348) );
BUFx10_ASAP7_75t_L g349 ( .A(n_256), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_47), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_170), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_58), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_9), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_163), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_66), .Y(n_355) );
INVxp33_ASAP7_75t_L g356 ( .A(n_217), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_240), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_40), .Y(n_358) );
CKINVDCx14_ASAP7_75t_R g359 ( .A(n_149), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_148), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_140), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_194), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_260), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_49), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_233), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_263), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_134), .Y(n_367) );
INVxp33_ASAP7_75t_L g368 ( .A(n_216), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_128), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_18), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_228), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_122), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_85), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_244), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_45), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_77), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_48), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_8), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_126), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_238), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_82), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_3), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_84), .Y(n_383) );
BUFx10_ASAP7_75t_L g384 ( .A(n_130), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_113), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_370), .B(n_0), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_274), .B(n_1), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_356), .B(n_2), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_276), .A2(n_19), .B(n_17), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_289), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_284), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_279), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_316), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_290), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_368), .B(n_2), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_279), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_281), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_270), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_312), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_312), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_340), .Y(n_402) );
OA21x2_ASAP7_75t_L g403 ( .A1(n_267), .A2(n_22), .B(n_21), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_281), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_299), .A2(n_24), .B(n_23), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_340), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_391), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_391), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_395), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_395), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_387), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_392), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_389), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_398), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_393), .B(n_357), .Y(n_417) );
INVx4_ASAP7_75t_L g418 ( .A(n_399), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_399), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_396), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_400), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_329), .B1(n_361), .B2(n_378), .Y(n_422) );
CKINVDCx6p67_ASAP7_75t_R g423 ( .A(n_388), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_418), .B(n_392), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_410), .Y(n_425) );
BUFx4_ASAP7_75t_L g426 ( .A(n_411), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_410), .Y(n_427) );
NOR2xp33_ASAP7_75t_SL g428 ( .A(n_418), .B(n_286), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_415), .A2(n_401), .B1(n_406), .B2(n_402), .Y(n_429) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_413), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_420), .A2(n_405), .B(n_388), .C(n_269), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_419), .B(n_397), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_421), .B(n_359), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_414), .B(n_382), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_407), .B(n_311), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_417), .B(n_275), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_422), .B(n_280), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_417), .B(n_282), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_414), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_423), .B(n_283), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_413), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_443), .A2(n_403), .B(n_374), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_431), .A2(n_403), .B(n_379), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_435), .A2(n_403), .B(n_339), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_441), .B(n_324), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_435), .A2(n_433), .B(n_439), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_441), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_434), .B(n_291), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_429), .B(n_292), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_440), .B(n_295), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_425), .Y(n_454) );
BUFx4f_ASAP7_75t_L g455 ( .A(n_430), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_427), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_437), .B(n_358), .C(n_327), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_428), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_424), .B(n_297), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_432), .A2(n_272), .B(n_271), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_436), .A2(n_277), .B(n_273), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_438), .A2(n_288), .B(n_278), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_444), .A2(n_296), .B(n_300), .C(n_298), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_442), .B(n_301), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_428), .B(n_317), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_449), .A2(n_306), .B(n_307), .C(n_303), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_450), .A2(n_323), .B1(n_346), .B2(n_343), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_447), .A2(n_314), .B(n_310), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_456), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_445), .A2(n_319), .B(n_318), .Y(n_471) );
AO31x2_ASAP7_75t_L g472 ( .A1(n_446), .A2(n_320), .A3(n_332), .B(n_330), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_460), .B(n_369), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_462), .A2(n_335), .B(n_333), .Y(n_474) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_463), .A2(n_342), .B(n_341), .Y(n_475) );
AOI221x1_ASAP7_75t_L g476 ( .A1(n_457), .A2(n_351), .B1(n_352), .B2(n_350), .C(n_344), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_448), .B(n_308), .C(n_281), .Y(n_477) );
OAI21x1_ASAP7_75t_L g478 ( .A1(n_454), .A2(n_362), .B(n_355), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_464), .B(n_372), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_458), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_461), .A2(n_373), .B(n_366), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_452), .B(n_308), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_465), .A2(n_376), .B(n_375), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_451), .B(n_349), .Y(n_485) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_466), .A2(n_287), .B(n_380), .Y(n_486) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_459), .A2(n_285), .B1(n_294), .B2(n_293), .Y(n_487) );
OAI21x1_ASAP7_75t_L g488 ( .A1(n_459), .A2(n_381), .B(n_364), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_455), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_455), .A2(n_377), .B(n_363), .Y(n_490) );
AO31x2_ASAP7_75t_L g491 ( .A1(n_447), .A2(n_416), .A3(n_404), .B(n_398), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_449), .B(n_308), .Y(n_492) );
AO22x2_ASAP7_75t_L g493 ( .A1(n_458), .A2(n_336), .B1(n_347), .B2(n_268), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_450), .Y(n_494) );
OAI21x1_ASAP7_75t_SL g495 ( .A1(n_469), .A2(n_384), .B(n_349), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_470), .Y(n_496) );
OAI21x1_ASAP7_75t_L g497 ( .A1(n_492), .A2(n_416), .B(n_328), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_482), .B(n_3), .Y(n_498) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_471), .A2(n_304), .B(n_302), .Y(n_499) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_477), .B(n_25), .Y(n_500) );
OAI21x1_ASAP7_75t_L g501 ( .A1(n_478), .A2(n_328), .B(n_326), .Y(n_501) );
OR2x6_ASAP7_75t_L g502 ( .A(n_489), .B(n_468), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_467), .A2(n_484), .B(n_474), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_494), .Y(n_504) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_473), .B(n_326), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_488), .Y(n_506) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_483), .A2(n_404), .B(n_398), .Y(n_507) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_475), .A2(n_328), .B(n_326), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g509 ( .A1(n_493), .A2(n_309), .B(n_305), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_487), .Y(n_510) );
OAI21x1_ASAP7_75t_L g511 ( .A1(n_475), .A2(n_383), .B(n_398), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g512 ( .A1(n_493), .A2(n_315), .B(n_313), .Y(n_512) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_476), .A2(n_322), .B(n_321), .Y(n_513) );
OAI21x1_ASAP7_75t_L g514 ( .A1(n_481), .A2(n_383), .B(n_404), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_479), .B(n_485), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_480), .B(n_384), .Y(n_516) );
OAI21x1_ASAP7_75t_L g517 ( .A1(n_491), .A2(n_383), .B(n_404), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_486), .B(n_4), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_490), .B(n_4), .Y(n_519) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_472), .A2(n_491), .A3(n_7), .B(n_5), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_491), .A2(n_331), .B(n_325), .Y(n_521) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_472), .A2(n_28), .B(n_27), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_472), .B(n_5), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_482), .B(n_6), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_477), .B(n_337), .C(n_334), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_482), .B(n_7), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_469), .A2(n_345), .B(n_338), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_468), .B(n_348), .Y(n_529) );
BUFx2_ASAP7_75t_SL g530 ( .A(n_489), .Y(n_530) );
OAI21x1_ASAP7_75t_L g531 ( .A1(n_469), .A2(n_32), .B(n_31), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_482), .B(n_8), .Y(n_532) );
INVx4_ASAP7_75t_SL g533 ( .A(n_489), .Y(n_533) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_469), .A2(n_35), .B(n_34), .Y(n_534) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_469), .A2(n_37), .B(n_36), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_470), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_489), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_469), .A2(n_360), .B(n_354), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_468), .B(n_365), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_536), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_496), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_536), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_528), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_532), .B(n_9), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_502), .Y(n_545) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_517), .A2(n_10), .B(n_11), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_506), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_498), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_504), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_510), .B(n_10), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_524), .Y(n_551) );
OAI21x1_ASAP7_75t_L g552 ( .A1(n_511), .A2(n_41), .B(n_39), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_526), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_515), .B(n_11), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_520), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_520), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_533), .B(n_12), .Y(n_558) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_508), .A2(n_43), .B(n_42), .Y(n_559) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_497), .A2(n_52), .B(n_50), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_523), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_505), .B(n_12), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_513), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_518), .Y(n_565) );
NOR2x1_ASAP7_75t_R g566 ( .A(n_530), .B(n_367), .Y(n_566) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_522), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_530), .B(n_509), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_503), .A2(n_385), .B1(n_371), .B2(n_15), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_529), .B(n_13), .Y(n_570) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_521), .A2(n_13), .B(n_14), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_533), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_516), .B(n_14), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_513), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_495), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_512), .B(n_15), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_539), .B(n_16), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_499), .A2(n_500), .B1(n_535), .B2(n_534), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_537), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_499), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_507), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_527), .B(n_16), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_531), .Y(n_583) );
INVx2_ASAP7_75t_SL g584 ( .A(n_501), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_507), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_514), .Y(n_586) );
CKINVDCx9p33_ASAP7_75t_R g587 ( .A(n_500), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_525), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_538), .Y(n_589) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_517), .A2(n_53), .B(n_55), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_536), .Y(n_591) );
INVxp67_ASAP7_75t_L g592 ( .A(n_523), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_496), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_502), .Y(n_594) );
OAI222xp33_ASAP7_75t_L g595 ( .A1(n_523), .A2(n_266), .B1(n_60), .B2(n_61), .C1(n_63), .C2(n_64), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_496), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_536), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_496), .Y(n_598) );
AOI222xp33_ASAP7_75t_L g599 ( .A1(n_510), .A2(n_57), .B1(n_65), .B2(n_67), .C1(n_68), .C2(n_69), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_536), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_536), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_496), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
BUFx2_ASAP7_75t_SL g604 ( .A(n_537), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_537), .Y(n_605) );
BUFx12f_ASAP7_75t_L g606 ( .A(n_502), .Y(n_606) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_517), .A2(n_71), .B(n_73), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_536), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_537), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_536), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_536), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_503), .A2(n_74), .B(n_75), .Y(n_612) );
AO31x2_ASAP7_75t_L g613 ( .A1(n_521), .A2(n_76), .A3(n_78), .B(n_79), .Y(n_613) );
OAI21x1_ASAP7_75t_L g614 ( .A1(n_517), .A2(n_80), .B(n_81), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_541), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_592), .B(n_86), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_540), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_561), .B(n_87), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g619 ( .A(n_606), .B(n_89), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_542), .B(n_591), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_593), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_597), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_596), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_602), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_544), .B(n_90), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_550), .B(n_91), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_565), .B(n_265), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_566), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_564), .B(n_92), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_545), .B(n_264), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_594), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_600), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_543), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_573), .B(n_96), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_601), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_592), .B(n_97), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_603), .B(n_98), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_608), .B(n_100), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_610), .B(n_611), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_570), .B(n_101), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_558), .B(n_103), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_569), .A2(n_104), .B1(n_105), .B2(n_109), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_568), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_549), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_558), .B(n_110), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_575), .B(n_572), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_546), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_548), .B(n_262), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_546), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_547), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_547), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_562), .Y(n_653) );
INVx5_ASAP7_75t_L g654 ( .A(n_605), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_551), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_554), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_556), .Y(n_657) );
BUFx2_ASAP7_75t_L g658 ( .A(n_566), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_555), .B(n_111), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_557), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_579), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_563), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_574), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_563), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_576), .B(n_261), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_604), .B(n_112), .Y(n_666) );
OAI222xp33_ASAP7_75t_L g667 ( .A1(n_569), .A2(n_115), .B1(n_116), .B2(n_117), .C1(n_118), .C2(n_120), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_609), .Y(n_668) );
BUFx3_ASAP7_75t_L g669 ( .A(n_577), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_553), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_582), .B(n_121), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_580), .B(n_259), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_571), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_553), .B(n_123), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_589), .B(n_258), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_588), .B(n_124), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_599), .A2(n_125), .B1(n_127), .B2(n_129), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_571), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_590), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_599), .A2(n_131), .B1(n_132), .B2(n_133), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_612), .B(n_136), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_612), .B(n_137), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_585), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_613), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_614), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_581), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_613), .B(n_257), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_613), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_581), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_587), .Y(n_690) );
BUFx3_ASAP7_75t_L g691 ( .A(n_560), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_578), .B(n_138), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_607), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_578), .B(n_139), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_583), .B(n_141), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_567), .B(n_142), .Y(n_696) );
INVx1_ASAP7_75t_SL g697 ( .A(n_587), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_607), .B(n_144), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_584), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_552), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_567), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_559), .B(n_145), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g703 ( .A1(n_586), .A2(n_146), .B(n_150), .C(n_152), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_595), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_621), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_668), .B(n_595), .Y(n_706) );
INVx5_ASAP7_75t_L g707 ( .A(n_654), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_654), .B(n_255), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_617), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_623), .B(n_153), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_645), .B(n_155), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_644), .B(n_157), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_655), .B(n_158), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_634), .B(n_161), .Y(n_714) );
NAND2xp33_ASAP7_75t_SL g715 ( .A(n_704), .B(n_162), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_620), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_620), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_656), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_617), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_615), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_661), .B(n_164), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_651), .B(n_165), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_633), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_633), .Y(n_724) );
BUFx2_ASAP7_75t_L g725 ( .A(n_654), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_622), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_644), .B(n_166), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_636), .B(n_168), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_629), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_624), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_663), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_652), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_658), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_653), .B(n_171), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_683), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_625), .B(n_172), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_669), .B(n_173), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_666), .Y(n_738) );
AND2x4_ASAP7_75t_L g739 ( .A(n_690), .B(n_174), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_640), .B(n_175), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_686), .B(n_176), .Y(n_741) );
AND2x4_ASAP7_75t_SL g742 ( .A(n_642), .B(n_177), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_664), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_647), .B(n_178), .Y(n_744) );
AND2x4_ASAP7_75t_L g745 ( .A(n_697), .B(n_179), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_647), .B(n_181), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_627), .B(n_183), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_657), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_626), .B(n_184), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_635), .B(n_185), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_662), .Y(n_751) );
NAND2x1p5_ASAP7_75t_L g752 ( .A(n_619), .B(n_253), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_689), .Y(n_753) );
INVxp67_ASAP7_75t_L g754 ( .A(n_641), .Y(n_754) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_618), .Y(n_755) );
NOR2x1_ASAP7_75t_R g756 ( .A(n_704), .B(n_186), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_638), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_646), .B(n_188), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_671), .B(n_190), .Y(n_759) );
AND2x4_ASAP7_75t_L g760 ( .A(n_670), .B(n_192), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_638), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_676), .B(n_195), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_657), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_660), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_618), .B(n_197), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_616), .B(n_198), .Y(n_766) );
BUFx2_ASAP7_75t_L g767 ( .A(n_699), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_637), .B(n_199), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_660), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_692), .B(n_200), .Y(n_770) );
OR2x2_ASAP7_75t_L g771 ( .A(n_705), .B(n_673), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_767), .B(n_701), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_709), .B(n_678), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_732), .B(n_678), .Y(n_774) );
INVx3_ASAP7_75t_L g775 ( .A(n_707), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_751), .B(n_704), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_716), .B(n_648), .Y(n_777) );
OR2x2_ASAP7_75t_L g778 ( .A(n_717), .B(n_701), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_726), .B(n_674), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_707), .B(n_680), .C(n_677), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_718), .B(n_650), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_709), .B(n_694), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_724), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_738), .B(n_696), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_733), .B(n_631), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_724), .B(n_696), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_754), .B(n_684), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_720), .B(n_688), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_719), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_723), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_731), .B(n_693), .Y(n_791) );
AND3x2_ASAP7_75t_L g792 ( .A(n_725), .B(n_681), .C(n_682), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_731), .B(n_675), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_735), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_735), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_730), .B(n_695), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_729), .B(n_659), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_755), .B(n_685), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_757), .B(n_685), .Y(n_799) );
AND2x4_ASAP7_75t_L g800 ( .A(n_707), .B(n_700), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_748), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_748), .B(n_687), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_761), .B(n_698), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_764), .B(n_628), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_743), .B(n_691), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_769), .B(n_630), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_753), .B(n_672), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_763), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_706), .B(n_702), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_714), .B(n_639), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_722), .B(n_649), .Y(n_811) );
INVxp33_ASAP7_75t_L g812 ( .A(n_785), .Y(n_812) );
NOR2x1p5_ASAP7_75t_SL g813 ( .A(n_771), .B(n_741), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_789), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_790), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_772), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_794), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_784), .B(n_745), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_795), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_783), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_801), .Y(n_821) );
AO21x1_ASAP7_75t_L g822 ( .A1(n_772), .A2(n_745), .B(n_776), .Y(n_822) );
OAI21xp5_ASAP7_75t_SL g823 ( .A1(n_792), .A2(n_742), .B(n_708), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_778), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_808), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_774), .B(n_760), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_781), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_809), .B(n_734), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_780), .A2(n_739), .B(n_712), .Y(n_829) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_798), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_791), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_773), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_773), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_777), .Y(n_834) );
INVx3_ASAP7_75t_L g835 ( .A(n_775), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_787), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_799), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_830), .B(n_803), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_832), .Y(n_839) );
OAI311xp33_ASAP7_75t_L g840 ( .A1(n_829), .A2(n_780), .A3(n_811), .B1(n_810), .C1(n_804), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_833), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_814), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_823), .A2(n_756), .B(n_775), .Y(n_843) );
OAI21xp33_ASAP7_75t_L g844 ( .A1(n_813), .A2(n_786), .B(n_805), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_823), .A2(n_797), .B1(n_739), .B2(n_782), .Y(n_845) );
INVxp67_ASAP7_75t_L g846 ( .A(n_827), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_815), .Y(n_847) );
XNOR2x1_ASAP7_75t_L g848 ( .A(n_829), .B(n_752), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_825), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_817), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_819), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_820), .Y(n_852) );
AND2x4_ASAP7_75t_L g853 ( .A(n_835), .B(n_800), .Y(n_853) );
INVxp67_ASAP7_75t_L g854 ( .A(n_831), .Y(n_854) );
OAI21xp33_ASAP7_75t_L g855 ( .A1(n_844), .A2(n_812), .B(n_836), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_840), .A2(n_824), .B1(n_837), .B2(n_834), .C(n_828), .Y(n_856) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_848), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_852), .Y(n_858) );
NAND2xp5_ASAP7_75t_SL g859 ( .A(n_845), .B(n_822), .Y(n_859) );
OAI31xp33_ASAP7_75t_L g860 ( .A1(n_843), .A2(n_835), .A3(n_818), .B(n_816), .Y(n_860) );
NOR3xp33_ASAP7_75t_SL g861 ( .A(n_842), .B(n_715), .C(n_747), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_846), .A2(n_821), .B1(n_826), .B2(n_737), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_854), .B(n_796), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_839), .B(n_788), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_841), .B(n_802), .Y(n_865) );
INVx4_ASAP7_75t_L g866 ( .A(n_858), .Y(n_866) );
AOI211xp5_ASAP7_75t_L g867 ( .A1(n_857), .A2(n_853), .B(n_847), .C(n_838), .Y(n_867) );
NOR2x1_ASAP7_75t_L g868 ( .A(n_859), .B(n_853), .Y(n_868) );
OAI211xp5_ASAP7_75t_L g869 ( .A1(n_860), .A2(n_749), .B(n_806), .C(n_759), .Y(n_869) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_855), .A2(n_851), .B(n_850), .Y(n_870) );
HAxp5_ASAP7_75t_SL g871 ( .A(n_862), .B(n_667), .CON(n_871), .SN(n_871) );
AOI21xp5_ASAP7_75t_L g872 ( .A1(n_856), .A2(n_849), .B(n_793), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g873 ( .A1(n_865), .A2(n_802), .B(n_746), .Y(n_873) );
NOR2xp33_ASAP7_75t_SL g874 ( .A(n_866), .B(n_863), .Y(n_874) );
NOR3xp33_ASAP7_75t_SL g875 ( .A(n_869), .B(n_643), .C(n_864), .Y(n_875) );
OAI21xp33_ASAP7_75t_L g876 ( .A1(n_868), .A2(n_861), .B(n_779), .Y(n_876) );
NOR3xp33_ASAP7_75t_L g877 ( .A(n_867), .B(n_744), .C(n_665), .Y(n_877) );
AND2x2_ASAP7_75t_SL g878 ( .A(n_871), .B(n_712), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_875), .B(n_872), .Y(n_879) );
NAND3xp33_ASAP7_75t_SL g880 ( .A(n_874), .B(n_870), .C(n_873), .Y(n_880) );
O2A1O1Ixp33_ASAP7_75t_L g881 ( .A1(n_876), .A2(n_711), .B(n_713), .C(n_740), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_878), .B(n_721), .Y(n_882) );
AOI31xp33_ASAP7_75t_L g883 ( .A1(n_879), .A2(n_758), .A3(n_750), .B(n_765), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_880), .Y(n_884) );
OR2x2_ASAP7_75t_L g885 ( .A(n_882), .B(n_877), .Y(n_885) );
OA22x2_ASAP7_75t_L g886 ( .A1(n_884), .A2(n_881), .B1(n_800), .B2(n_770), .Y(n_886) );
XNOR2xp5_ASAP7_75t_L g887 ( .A(n_885), .B(n_710), .Y(n_887) );
XOR2x2_ASAP7_75t_L g888 ( .A(n_883), .B(n_762), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_886), .A2(n_632), .B1(n_807), .B2(n_728), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_887), .Y(n_890) );
OR2x6_ASAP7_75t_L g891 ( .A(n_888), .B(n_727), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g892 ( .A1(n_890), .A2(n_768), .B1(n_766), .B2(n_736), .C(n_703), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_891), .A2(n_760), .B(n_679), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_889), .A2(n_679), .B(n_202), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_892), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_894), .B(n_893), .Y(n_896) );
OA21x2_ASAP7_75t_L g897 ( .A1(n_895), .A2(n_201), .B(n_205), .Y(n_897) );
AOI21xp33_ASAP7_75t_L g898 ( .A1(n_897), .A2(n_896), .B(n_206), .Y(n_898) );
OAI21xp33_ASAP7_75t_SL g899 ( .A1(n_898), .A2(n_208), .B(n_209), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_899), .A2(n_210), .B(n_212), .Y(n_900) );
endmodule