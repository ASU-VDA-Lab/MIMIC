module real_jpeg_370_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_43;
wire n_57;
wire n_37;
wire n_21;
wire n_54;
wire n_73;
wire n_65;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_58;
wire n_31;
wire n_67;
wire n_52;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_71;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_70;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_26;
wire n_19;
wire n_48;
wire n_30;
wire n_56;
wire n_74;
wire n_16;
wire n_15;
wire n_13;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_15),
.B1(n_23),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_3),
.B(n_18),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_3),
.B(n_15),
.C(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_15),
.B1(n_23),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_6),
.A2(n_15),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_22),
.B1(n_49),
.B2(n_50),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_15),
.B1(n_23),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_8),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_58),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_37),
.B(n_57),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_27),
.B(n_36),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_20),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_17),
.Y(n_14)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_18),
.A2(n_21),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_18),
.A2(n_25),
.B1(n_42),
.B2(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_33),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_29),
.A2(n_47),
.B1(n_53),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_48),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_32),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_44),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_54),
.B2(n_56),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AO22x2_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_50),
.B1(n_68),
.B2(n_70),
.Y(n_67)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);


endmodule