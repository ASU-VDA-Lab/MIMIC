module fake_jpeg_2072_n_537 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_537);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_49),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_51),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_55),
.B(n_62),
.Y(n_161)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_57),
.Y(n_164)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g144 ( 
.A(n_59),
.Y(n_144)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_0),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_42),
.B(n_29),
.Y(n_117)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_70),
.B(n_74),
.Y(n_141)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_7),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_17),
.B(n_7),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_77),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_8),
.Y(n_77)
);

BUFx12f_ASAP7_75t_SL g78 ( 
.A(n_18),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_8),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_80),
.B(n_89),
.Y(n_160)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_37),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_44),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_44),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_117),
.B(n_27),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_44),
.B1(n_30),
.B2(n_22),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_118),
.A2(n_133),
.B1(n_147),
.B2(n_144),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_140),
.Y(n_179)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_133)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_150),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_155),
.Y(n_192)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_52),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_95),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_54),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_181),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_41),
.B1(n_45),
.B2(n_24),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_45),
.B1(n_41),
.B2(n_27),
.Y(n_217)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_171),
.Y(n_243)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_56),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_174),
.B(n_176),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_58),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_209),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_60),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_178),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_40),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_107),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_185),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_184),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_105),
.B(n_91),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_108),
.B(n_136),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_193),
.Y(n_229)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_187),
.Y(n_240)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_71),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_208),
.Y(n_228)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_64),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_198),
.Y(n_236)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_67),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_212),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_24),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_99),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_215),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_217),
.A2(n_104),
.B1(n_209),
.B2(n_26),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_126),
.B1(n_142),
.B2(n_124),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_172),
.B1(n_145),
.B2(n_210),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_129),
.C(n_164),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_223),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_133),
.Y(n_223)
);

AO22x2_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_164),
.B1(n_126),
.B2(n_142),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_209),
.B(n_191),
.C(n_197),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_178),
.A2(n_106),
.B1(n_125),
.B2(n_167),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_230),
.A2(n_233),
.B1(n_209),
.B2(n_204),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_181),
.A2(n_167),
.B1(n_134),
.B2(n_132),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_111),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_251),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_173),
.B(n_148),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_169),
.B1(n_134),
.B2(n_130),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_253),
.A2(n_277),
.B1(n_230),
.B2(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_180),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_254),
.B(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_259),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_261),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_257),
.A2(n_268),
.B1(n_272),
.B2(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_169),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_SL g306 ( 
.A(n_265),
.B(n_267),
.C(n_227),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_169),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_225),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_180),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_274),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_222),
.A2(n_204),
.B1(n_210),
.B2(n_132),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_242),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_238),
.A2(n_188),
.B1(n_26),
.B2(n_32),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_190),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_228),
.B(n_203),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_216),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_214),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_281),
.B(n_240),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_234),
.A2(n_48),
.B(n_28),
.C(n_32),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_213),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_241),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_234),
.A2(n_124),
.B1(n_128),
.B2(n_130),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_218),
.B1(n_233),
.B2(n_240),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_259),
.A2(n_248),
.B1(n_234),
.B2(n_246),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_297),
.B1(n_302),
.B2(n_309),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_280),
.Y(n_286)
);

INVx13_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_298),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_220),
.C(n_252),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_300),
.C(n_273),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_266),
.A2(n_262),
.B(n_271),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_293),
.B(n_300),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_253),
.A2(n_262),
.B1(n_268),
.B2(n_282),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_295),
.A2(n_303),
.B1(n_270),
.B2(n_274),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_252),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_265),
.A2(n_227),
.B1(n_243),
.B2(n_219),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_275),
.A2(n_227),
.B1(n_217),
.B2(n_250),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_278),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_305),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_310),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_258),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_265),
.A2(n_250),
.B1(n_131),
.B2(n_94),
.Y(n_309)
);

AO22x1_ASAP7_75t_L g310 ( 
.A1(n_255),
.A2(n_216),
.B1(n_235),
.B2(n_245),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_254),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_285),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_267),
.A2(n_237),
.B(n_245),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_321),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_261),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_317),
.B(n_337),
.Y(n_362)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_267),
.B(n_255),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_320),
.A2(n_326),
.B(n_292),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_291),
.C(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_325),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_269),
.B(n_281),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_283),
.B1(n_257),
.B2(n_263),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_327),
.A2(n_345),
.B1(n_299),
.B2(n_244),
.Y(n_371)
);

CKINVDCx12_ASAP7_75t_R g329 ( 
.A(n_304),
.Y(n_329)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_260),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_346),
.Y(n_351)
);

OR2x4_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_276),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g367 ( 
.A1(n_335),
.A2(n_342),
.B(n_314),
.Y(n_367)
);

CKINVDCx10_ASAP7_75t_R g336 ( 
.A(n_310),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_336),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_226),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_338),
.A2(n_288),
.B1(n_303),
.B2(n_298),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_305),
.B(n_226),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_341),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_235),
.Y(n_341)
);

AO21x1_ASAP7_75t_SL g342 ( 
.A1(n_306),
.A2(n_145),
.B(n_137),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_315),
.A2(n_250),
.B1(n_237),
.B2(n_131),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_244),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_296),
.Y(n_354)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_313),
.A3(n_302),
.B1(n_301),
.B2(n_310),
.Y(n_349)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_347),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_307),
.C(n_284),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_366),
.C(n_380),
.Y(n_390)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_355),
.A2(n_371),
.B1(n_374),
.B2(n_381),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_321),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_356),
.B(n_365),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_289),
.Y(n_360)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_318),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_309),
.C(n_314),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_369),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_299),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_368),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_339),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_319),
.A2(n_221),
.B1(n_231),
.B2(n_215),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_372),
.A2(n_327),
.B1(n_345),
.B2(n_346),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_319),
.A2(n_331),
.B1(n_338),
.B2(n_325),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_231),
.Y(n_375)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_221),
.Y(n_378)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_194),
.C(n_183),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_319),
.A2(n_35),
.B1(n_207),
.B2(n_201),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_355),
.A2(n_332),
.B1(n_331),
.B2(n_328),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_382),
.A2(n_386),
.B1(n_401),
.B2(n_403),
.Y(n_430)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_336),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_383),
.B(n_202),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_384),
.A2(n_394),
.B1(n_402),
.B2(n_409),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_374),
.A2(n_328),
.B1(n_326),
.B2(n_342),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_397),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_343),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_407),
.C(n_364),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_333),
.C(n_348),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_396),
.C(n_372),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_368),
.A2(n_329),
.B1(n_347),
.B2(n_324),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_356),
.C(n_361),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_183),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_192),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_399),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_192),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_350),
.A2(n_358),
.B1(n_364),
.B2(n_351),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_35),
.B1(n_85),
.B2(n_207),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_350),
.A2(n_46),
.B1(n_92),
.B2(n_72),
.Y(n_403)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_406),
.A2(n_400),
.B1(n_376),
.B2(n_397),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_359),
.B(n_195),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_362),
.A2(n_358),
.B1(n_380),
.B2(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_411),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_389),
.B(n_393),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_412),
.B(n_429),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_368),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_419),
.Y(n_446)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_401),
.Y(n_415)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_388),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_418),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_363),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_410),
.B(n_349),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_423),
.Y(n_448)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_367),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_408),
.A2(n_392),
.B(n_383),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_425),
.Y(n_454)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_405),
.A2(n_379),
.B1(n_377),
.B2(n_370),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_426),
.A2(n_434),
.B1(n_437),
.B2(n_211),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_377),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_428),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_357),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_357),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_432),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_175),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_410),
.B(n_376),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_396),
.C(n_403),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_398),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_384),
.B1(n_382),
.B2(n_386),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_438),
.A2(n_430),
.B1(n_440),
.B2(n_444),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_46),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_202),
.C(n_175),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_447),
.Y(n_464)
);

INVx13_ASAP7_75t_L g443 ( 
.A(n_424),
.Y(n_443)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_148),
.C(n_159),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_426),
.A2(n_69),
.B1(n_79),
.B2(n_139),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_449),
.A2(n_450),
.B1(n_434),
.B2(n_430),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_436),
.A2(n_154),
.B1(n_101),
.B2(n_211),
.Y(n_450)
);

INVx13_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_159),
.C(n_187),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_457),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_86),
.C(n_97),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_416),
.B(n_36),
.C(n_137),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_459),
.B(n_422),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_462),
.Y(n_495)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_413),
.C(n_433),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_463),
.A2(n_479),
.B1(n_29),
.B2(n_38),
.Y(n_483)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_466),
.B(n_471),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_452),
.A2(n_428),
.B(n_427),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_469),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_454),
.A2(n_420),
.B(n_422),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_36),
.C(n_112),
.Y(n_471)
);

OA21x2_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_28),
.B(n_48),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_48),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_165),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_473),
.B(n_0),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_442),
.C(n_439),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_474),
.B(n_475),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_455),
.A2(n_443),
.B(n_448),
.Y(n_477)
);

NAND3xp33_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_447),
.C(n_459),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_449),
.A2(n_450),
.B1(n_458),
.B2(n_448),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_478),
.A2(n_461),
.B1(n_470),
.B2(n_463),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_456),
.A2(n_46),
.B1(n_100),
.B2(n_38),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_482),
.B1(n_483),
.B2(n_59),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_474),
.B(n_446),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_485),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_468),
.A2(n_451),
.B1(n_457),
.B2(n_30),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_28),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_10),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_465),
.A2(n_469),
.B(n_464),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_489),
.A2(n_479),
.B(n_472),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_476),
.B(n_38),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_493),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_466),
.B(n_467),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_496),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_114),
.C(n_150),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_478),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_505),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_484),
.A2(n_462),
.B(n_471),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_498),
.A2(n_20),
.B(n_9),
.Y(n_516)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_499),
.A2(n_500),
.B(n_39),
.Y(n_520)
);

NOR3xp33_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_472),
.C(n_114),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_504),
.B(n_509),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_155),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_155),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_507),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_150),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_491),
.B(n_10),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_9),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_494),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_514),
.B(n_519),
.Y(n_521)
);

AOI322xp5_ASAP7_75t_L g513 ( 
.A1(n_500),
.A2(n_480),
.A3(n_488),
.B1(n_496),
.B2(n_486),
.C1(n_20),
.C2(n_102),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_513),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_508),
.A2(n_87),
.B(n_20),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_516),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_501),
.B(n_8),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_503),
.B(n_39),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_503),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_525),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_498),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_527),
.A3(n_519),
.B1(n_12),
.B2(n_9),
.C1(n_5),
.C2(n_1),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_9),
.C(n_3),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_517),
.A2(n_14),
.B(n_12),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_530),
.B(n_529),
.Y(n_533)
);

OA22x2_ASAP7_75t_L g531 ( 
.A1(n_521),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_522),
.B(n_5),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_533),
.B1(n_2),
.B2(n_6),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_534),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_2),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_2),
.B(n_6),
.Y(n_537)
);


endmodule