module fake_jpeg_11863_n_580 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_580);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_65),
.B(n_77),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_26),
.Y(n_68)
);

CKINVDCx9p33_ASAP7_75t_R g160 ( 
.A(n_68),
.Y(n_160)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_71),
.Y(n_161)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_24),
.B(n_16),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_88),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_27),
.B(n_2),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_2),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_96),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_2),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_21),
.A2(n_3),
.B(n_4),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_23),
.B(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_106),
.Y(n_128)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

CKINVDCx9p33_ASAP7_75t_R g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g206 ( 
.A(n_105),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_107),
.B(n_115),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_110),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_55),
.B(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_27),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_48),
.Y(n_153)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_20),
.Y(n_114)
);

INVx2_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_19),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_117),
.Y(n_170)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_120),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_47),
.B(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_5),
.Y(n_136)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

NOR2x1_ASAP7_75t_R g199 ( 
.A(n_122),
.B(n_125),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_123),
.B(n_124),
.Y(n_186)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_41),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_127),
.Y(n_188)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_136),
.B(n_200),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_100),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_141),
.B(n_143),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_40),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_67),
.B(n_36),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_144),
.B(n_167),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_73),
.A2(n_37),
.B1(n_47),
.B2(n_56),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_150),
.A2(n_182),
.B1(n_160),
.B2(n_178),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_34),
.C(n_31),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_83),
.A2(n_46),
.B1(n_37),
.B2(n_43),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_165),
.A2(n_187),
.B1(n_197),
.B2(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_86),
.B(n_40),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_123),
.B1(n_116),
.B2(n_115),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_181),
.B1(n_30),
.B2(n_59),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_83),
.B(n_43),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_175),
.B(n_190),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_109),
.B(n_36),
.C(n_60),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_180),
.B(n_5),
.C(n_11),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_110),
.A2(n_60),
.B1(n_38),
.B2(n_52),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_74),
.A2(n_48),
.B1(n_49),
.B2(n_56),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_88),
.B(n_51),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_183),
.B(n_185),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_90),
.B(n_51),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_69),
.A2(n_46),
.B1(n_58),
.B2(n_57),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_68),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_75),
.B(n_49),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_192),
.B(n_193),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_81),
.B(n_52),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_99),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_194),
.B(n_196),
.Y(n_271)
);

FAx1_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_46),
.CI(n_31),
.CON(n_195),
.SN(n_195)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_31),
.B(n_30),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_104),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_89),
.A2(n_53),
.B1(n_58),
.B2(n_57),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_95),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_97),
.A2(n_54),
.B1(n_53),
.B2(n_38),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_102),
.B(n_54),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_203),
.B(n_181),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_35),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_205),
.B(n_14),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_107),
.B(n_35),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_208),
.B(n_148),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_160),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_211),
.B(n_221),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_213),
.B(n_226),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_106),
.B1(n_105),
.B2(n_35),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_214),
.A2(n_257),
.B1(n_264),
.B2(n_265),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_128),
.B(n_34),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_215),
.Y(n_324)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_135),
.Y(n_217)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_217),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_141),
.B(n_34),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_219),
.B(n_130),
.C(n_139),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_222),
.A2(n_249),
.B(n_252),
.Y(n_299)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_223),
.Y(n_285)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_224),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_30),
.B1(n_59),
.B2(n_25),
.Y(n_225)
);

OAI22x1_ASAP7_75t_L g332 ( 
.A1(n_225),
.A2(n_227),
.B1(n_229),
.B2(n_239),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_59),
.B1(n_25),
.B2(n_7),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_131),
.A2(n_59),
.B1(n_25),
.B2(n_7),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_137),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_230),
.B(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_154),
.Y(n_233)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_137),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_235),
.Y(n_319)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_161),
.A2(n_59),
.B1(n_25),
.B2(n_8),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_183),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_241),
.B(n_248),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_161),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_191),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_244),
.A2(n_250),
.B1(n_254),
.B2(n_259),
.Y(n_286)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_157),
.Y(n_246)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_130),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_158),
.A2(n_11),
.B(n_12),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_191),
.A2(n_174),
.B1(n_138),
.B2(n_185),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_149),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_251),
.B(n_260),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_167),
.A2(n_11),
.B(n_12),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_174),
.A2(n_12),
.B1(n_14),
.B2(n_138),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_261),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_164),
.A2(n_171),
.B1(n_204),
.B2(n_169),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_157),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_258),
.B(n_232),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_132),
.A2(n_134),
.B1(n_147),
.B2(n_198),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_146),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_162),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_266),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_164),
.A2(n_204),
.B1(n_169),
.B2(n_148),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_143),
.A2(n_144),
.B1(n_136),
.B2(n_180),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_164),
.A2(n_199),
.B(n_209),
.C(n_129),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_267),
.A2(n_219),
.B(n_216),
.C(n_215),
.Y(n_313)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_166),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_280),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_170),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_269),
.B(n_272),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_147),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_166),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_179),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_275),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_210),
.A2(n_142),
.B1(n_188),
.B2(n_186),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_274),
.A2(n_219),
.B1(n_215),
.B2(n_253),
.Y(n_331)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_132),
.A2(n_134),
.B1(n_198),
.B2(n_149),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_276),
.A2(n_277),
.B1(n_258),
.B2(n_238),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_151),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_189),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_177),
.B(n_199),
.CI(n_129),
.CON(n_279),
.SN(n_279)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_279),
.B(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_281),
.B(n_156),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_289),
.B(n_292),
.Y(n_370)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_216),
.A2(n_133),
.A3(n_156),
.B1(n_139),
.B2(n_184),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_298),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_133),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_296),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_151),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_271),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_212),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_331),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_152),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_302),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_152),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_241),
.B(n_159),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_314),
.Y(n_377)
);

O2A1O1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_222),
.A2(n_157),
.B(n_155),
.C(n_184),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_310),
.B(n_330),
.Y(n_378)
);

NOR2x1_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_217),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_234),
.B(n_265),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_316),
.B(n_320),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_281),
.A2(n_159),
.B1(n_163),
.B2(n_155),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_317),
.A2(n_226),
.B1(n_213),
.B2(n_261),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_252),
.B(n_163),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_220),
.B(n_269),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_328),
.B(n_335),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_267),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_333),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_334),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_247),
.B(n_279),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_211),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_223),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_237),
.B(n_279),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_262),
.C(n_256),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_218),
.B1(n_282),
.B2(n_248),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_341),
.A2(n_348),
.B1(n_354),
.B2(n_356),
.Y(n_417)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_249),
.C(n_267),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_349),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_344),
.A2(n_346),
.B1(n_366),
.B2(n_372),
.Y(n_386)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_345),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_323),
.A2(n_233),
.B1(n_231),
.B2(n_280),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_301),
.B1(n_302),
.B2(n_296),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_293),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_350),
.A2(n_371),
.B(n_319),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_289),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_311),
.A2(n_277),
.B1(n_224),
.B2(n_240),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_240),
.B1(n_268),
.B2(n_266),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_300),
.B(n_272),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_357),
.B(n_364),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_323),
.A2(n_245),
.B1(n_278),
.B2(n_275),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

BUFx2_ASAP7_75t_SL g388 ( 
.A(n_360),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_330),
.A2(n_277),
.B1(n_228),
.B2(n_236),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_362),
.A2(n_367),
.B1(n_382),
.B2(n_336),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_243),
.C(n_235),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_381),
.C(n_334),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_323),
.A2(n_246),
.B1(n_251),
.B2(n_287),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_330),
.A2(n_299),
.B1(n_311),
.B2(n_294),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_298),
.B(n_321),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_368),
.Y(n_402)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_283),
.Y(n_369)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

OR2x2_ASAP7_75t_SL g371 ( 
.A(n_313),
.B(n_338),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_287),
.A2(n_330),
.B1(n_310),
.B2(n_314),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_337),
.A2(n_317),
.B1(n_291),
.B2(n_324),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_373),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_328),
.B(n_312),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_374),
.B(n_307),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_283),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_380),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_305),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_292),
.B(n_339),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_299),
.A2(n_309),
.B1(n_324),
.B2(n_314),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_290),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_383),
.B(n_394),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_385),
.B(n_353),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_387),
.A2(n_418),
.B(n_361),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_354),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_390),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_346),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_372),
.A2(n_286),
.B1(n_336),
.B2(n_332),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_398),
.B(n_412),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_379),
.A2(n_332),
.B1(n_290),
.B2(n_303),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_399),
.B(n_410),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_356),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_413),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_370),
.C(n_381),
.Y(n_422)
);

BUFx12_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_405),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_340),
.A2(n_307),
.B1(n_303),
.B2(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_406),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_369),
.Y(n_409)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_409),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_327),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_379),
.A2(n_306),
.B1(n_297),
.B2(n_288),
.Y(n_411)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_371),
.A2(n_306),
.B(n_285),
.C(n_288),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_284),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_297),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_378),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_345),
.B(n_315),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_416),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_378),
.A2(n_325),
.B1(n_315),
.B2(n_285),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_423),
.C(n_427),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_370),
.C(n_365),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_430),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_367),
.C(n_351),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_435),
.C(n_437),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_436),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_383),
.B(n_351),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_410),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_352),
.C(n_382),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_417),
.A2(n_366),
.B1(n_352),
.B2(n_377),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_438),
.A2(n_386),
.B1(n_399),
.B2(n_395),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_403),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_442),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_348),
.C(n_377),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_418),
.C(n_361),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_411),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_362),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_444),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_406),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_447),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_387),
.A2(n_350),
.B(n_392),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_446),
.B(n_350),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_398),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_400),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_400),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_396),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_451),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_443),
.B(n_396),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_447),
.B(n_402),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_452),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_414),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_470),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_421),
.A2(n_394),
.B1(n_395),
.B2(n_386),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_454),
.A2(n_459),
.B(n_466),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_392),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_463),
.Y(n_485)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_408),
.Y(n_457)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_457),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_458),
.A2(n_434),
.B1(n_439),
.B2(n_449),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_427),
.B(n_417),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_460),
.B(n_428),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_445),
.A2(n_401),
.B1(n_390),
.B2(n_409),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_434),
.B1(n_442),
.B2(n_444),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_415),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_423),
.B(n_363),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_477),
.Y(n_486)
);

A2O1A1Ixp33_ASAP7_75t_SL g466 ( 
.A1(n_424),
.A2(n_412),
.B(n_342),
.C(n_413),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_439),
.A2(n_419),
.B(n_424),
.Y(n_470)
);

XOR2x2_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_341),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_446),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_420),
.B(n_416),
.Y(n_474)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_430),
.C(n_449),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_426),
.B(n_384),
.Y(n_476)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_476),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_384),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_479),
.A2(n_502),
.B1(n_454),
.B2(n_472),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_481),
.A2(n_494),
.B1(n_470),
.B2(n_462),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_483),
.B(n_487),
.Y(n_522)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_470),
.Y(n_484)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_484),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_436),
.C(n_438),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_492),
.C(n_498),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_455),
.B(n_426),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_495),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_444),
.C(n_419),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_458),
.A2(n_342),
.B1(n_389),
.B2(n_448),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_460),
.B(n_428),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_475),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_425),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_425),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_500),
.C(n_477),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_440),
.C(n_429),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_461),
.A2(n_391),
.B1(n_431),
.B2(n_429),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_504),
.B(n_507),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_456),
.Y(n_505)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_505),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_506),
.B(n_517),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_508),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_484),
.A2(n_467),
.B(n_468),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_510),
.A2(n_521),
.B(n_480),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_487),
.A2(n_467),
.B1(n_473),
.B2(n_466),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_480),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_457),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_512),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_465),
.C(n_471),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_513),
.B(n_514),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_467),
.C(n_466),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_490),
.B(n_466),
.C(n_360),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_500),
.C(n_485),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_479),
.A2(n_344),
.B1(n_391),
.B2(n_388),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_375),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_520),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_482),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_497),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_481),
.A2(n_388),
.B1(n_393),
.B2(n_405),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_492),
.A2(n_405),
.B(n_393),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_530),
.Y(n_545)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_525),
.Y(n_544)
);

NOR2xp67_ASAP7_75t_SL g542 ( 
.A(n_529),
.B(n_531),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_491),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_505),
.B(n_493),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_538),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_510),
.A2(n_483),
.B(n_478),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_534),
.A2(n_535),
.B(n_514),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_516),
.A2(n_494),
.B(n_495),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_503),
.B(n_485),
.C(n_486),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_532),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_539),
.B(n_551),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_518),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_540),
.A2(n_546),
.B1(n_520),
.B2(n_496),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_503),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_541),
.B(n_547),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_536),
.A2(n_511),
.B(n_515),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_509),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_526),
.A2(n_527),
.B1(n_528),
.B2(n_537),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_524),
.B(n_521),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_524),
.B(n_531),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_322),
.Y(n_561)
);

AND2x4_ASAP7_75t_SL g555 ( 
.A(n_550),
.B(n_522),
.Y(n_555)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_528),
.Y(n_551)
);

AOI322xp5_ASAP7_75t_L g552 ( 
.A1(n_540),
.A2(n_534),
.A3(n_530),
.B1(n_506),
.B2(n_527),
.C1(n_517),
.C2(n_535),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_552),
.B(n_553),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_538),
.C(n_523),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_513),
.C(n_522),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_554),
.B(n_559),
.Y(n_562)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_555),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_557),
.A2(n_550),
.B(n_322),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_558),
.Y(n_564)
);

AOI322xp5_ASAP7_75t_L g559 ( 
.A1(n_544),
.A2(n_405),
.A3(n_393),
.B1(n_509),
.B2(n_486),
.C1(n_284),
.C2(n_329),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_561),
.B(n_542),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_545),
.C(n_546),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_566),
.B(n_568),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_567),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_564),
.B(n_556),
.C(n_560),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_569),
.B(n_570),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_562),
.B(n_556),
.C(n_552),
.Y(n_570)
);

AOI21xp33_ASAP7_75t_L g573 ( 
.A1(n_563),
.A2(n_329),
.B(n_308),
.Y(n_573)
);

AOI21xp33_ASAP7_75t_L g576 ( 
.A1(n_573),
.A2(n_308),
.B(n_572),
.Y(n_576)
);

OAI21x1_ASAP7_75t_SL g574 ( 
.A1(n_571),
.A2(n_565),
.B(n_564),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_574),
.Y(n_577)
);

FAx1_ASAP7_75t_SL g578 ( 
.A(n_576),
.B(n_569),
.CI(n_575),
.CON(n_578),
.SN(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_578),
.B(n_577),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_578),
.Y(n_580)
);


endmodule