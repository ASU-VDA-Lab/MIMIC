module real_jpeg_1036_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_249;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_295;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_1),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_29),
.B1(n_35),
.B2(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_46),
.B1(n_51),
.B2(n_75),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_44),
.B1(n_46),
.B2(n_51),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_2),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_44),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_46),
.B1(n_51),
.B2(n_73),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_73),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_5),
.A2(n_46),
.B1(n_51),
.B2(n_107),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_107),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_5),
.A2(n_29),
.B1(n_35),
.B2(n_107),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_6),
.A2(n_46),
.B1(n_51),
.B2(n_56),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_6),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_56),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_8),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_46),
.B1(n_51),
.B2(n_152),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_152),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_152),
.Y(n_263)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_12),
.A2(n_46),
.B1(n_51),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_12),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_88),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_88),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_13),
.A2(n_36),
.B1(n_65),
.B2(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_15),
.B(n_40),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_15),
.B(n_153),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_15),
.A2(n_51),
.B(n_83),
.C(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_15),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_15),
.B(n_85),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_15),
.A2(n_46),
.B1(n_51),
.B2(n_203),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_15),
.B(n_29),
.C(n_68),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_15),
.B(n_32),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_101),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_128),
.B1(n_300),
.B2(n_301),
.Y(n_18)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_19),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_126),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_21),
.B(n_111),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.C(n_92),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_22),
.A2(n_23),
.B1(n_77),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_60),
.B2(n_76),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_59),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_26),
.A2(n_38),
.B(n_76),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_26),
.A2(n_59),
.B1(n_61),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_27),
.A2(n_32),
.B1(n_97),
.B2(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_27),
.A2(n_203),
.B(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_28),
.A2(n_31),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_28),
.A2(n_31),
.B1(n_178),
.B2(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_28),
.B(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_28),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_28),
.A2(n_31),
.B1(n_234),
.B2(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_29),
.A2(n_35),
.B1(n_68),
.B2(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_29),
.B(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_31),
.A2(n_193),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_31),
.B(n_207),
.Y(n_236)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_32),
.A2(n_206),
.B(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B(n_53),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_39),
.A2(n_45),
.B1(n_108),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_41),
.B1(n_49),
.B2(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_41),
.A2(n_49),
.A3(n_51),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_41),
.A2(n_108),
.B(n_203),
.C(n_212),
.Y(n_211)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_45),
.B(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_45),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_45),
.A2(n_53),
.B(n_167),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_45)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_46),
.B(n_52),
.Y(n_175)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_49),
.Y(n_52)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_83),
.B(n_84),
.C(n_85),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_57),
.A2(n_106),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_61),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_70),
.B1(n_74),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_62),
.A2(n_70),
.B1(n_196),
.B2(n_230),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_62),
.A2(n_198),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_72),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_63),
.A2(n_101),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_63),
.A2(n_100),
.B1(n_101),
.B2(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_63),
.A2(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_63),
.B(n_199),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_64)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_66),
.B1(n_83),
.B2(n_86),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_65),
.A2(n_86),
.B(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_66),
.B(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_70),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_70),
.A2(n_219),
.B(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_91),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_80),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_89),
.B1(n_90),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_81),
.A2(n_169),
.B(n_171),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_81),
.A2(n_171),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_82),
.A2(n_85),
.B1(n_170),
.B2(n_187),
.Y(n_215)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_85),
.B(n_149),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_89),
.A2(n_103),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_89),
.A2(n_148),
.B(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_104),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_94),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_101),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_102),
.B(n_104),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_109),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_110),
.B(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_125),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_124),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_128),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_154),
.B(n_299),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_130),
.B(n_133),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_139),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.C(n_150),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_141),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_142),
.B(n_144),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_143),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_180),
.B(n_298),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_156),
.B(n_158),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.C(n_165),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_159),
.B(n_163),
.Y(n_283)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_165),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.C(n_172),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_166),
.B(n_168),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_172),
.B(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_176),
.B1(n_177),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI31xp33_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_280),
.A3(n_290),
.B(n_295),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_224),
.B(n_279),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_208),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_183),
.B(n_208),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.C(n_200),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_189),
.C(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_194),
.B(n_200),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_204),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_220),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_209),
.B(n_221),
.C(n_223),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_210),
.B(n_215),
.C(n_216),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_274),
.B(n_278),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_243),
.B(n_273),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_237),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.C(n_232),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_233),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_255),
.B(n_272),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_251),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_266),
.B(n_271),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_264),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_284),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_294),
.Y(n_296)
);


endmodule