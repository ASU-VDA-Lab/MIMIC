module real_jpeg_22862_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_0),
.B(n_47),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_0),
.B(n_66),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_0),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_1),
.B(n_33),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_1),
.B(n_52),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_1),
.B(n_49),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_1),
.B(n_47),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_1),
.B(n_66),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_2),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_2),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_33),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_2),
.B(n_52),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_7),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_7),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_7),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_7),
.B(n_33),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_7),
.B(n_52),
.Y(n_264)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_33),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_10),
.B(n_17),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_10),
.B(n_52),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_10),
.B(n_49),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_10),
.B(n_47),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_10),
.B(n_66),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_10),
.B(n_27),
.Y(n_278)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_12),
.B(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_12),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_12),
.B(n_33),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_12),
.B(n_52),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_12),
.B(n_49),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_12),
.B(n_47),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_12),
.B(n_66),
.Y(n_284)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_47),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_14),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_14),
.B(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_14),
.B(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_14),
.B(n_220),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_14),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_14),
.B(n_52),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_15),
.B(n_49),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_15),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_15),
.B(n_33),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_15),
.B(n_47),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_15),
.B(n_66),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_15),
.B(n_27),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_52),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_16),
.B(n_33),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_16),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_16),
.B(n_49),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_16),
.B(n_47),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_16),
.B(n_66),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_16),
.B(n_27),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_16),
.B(n_73),
.Y(n_298)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_17),
.Y(n_150)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_17),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.C(n_97),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_21),
.B(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.C(n_70),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_22),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_23),
.B(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_30),
.C(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_60),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_30),
.B(n_86),
.C(n_96),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_30),
.A2(n_38),
.B1(n_85),
.B2(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_32),
.B(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_36),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_36),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.C(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_39),
.B(n_45),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_40),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_41),
.A2(n_42),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_44),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_45),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.CI(n_51),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_48),
.C(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_52),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_54),
.B(n_70),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_55),
.A2(n_56),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.C(n_62),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_57),
.B(n_62),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_59),
.B(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_61),
.B(n_63),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_76),
.C(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_65),
.A2(n_69),
.B1(n_77),
.B2(n_337),
.Y(n_336)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_69),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_79),
.A2(n_80),
.B1(n_97),
.B2(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_91),
.C(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_83),
.B(n_86),
.C(n_87),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_88),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.C(n_94),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_93),
.CI(n_94),
.CON(n_102),
.SN(n_102)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_97),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_104),
.C(n_107),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.C(n_102),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_99),
.B(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_101),
.B(n_102),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_102),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_110),
.C(n_113),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_119),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_121),
.CI(n_122),
.CON(n_119),
.SN(n_119)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_348),
.C(n_349),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_340),
.C(n_341),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_324),
.C(n_325),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_300),
.C(n_301),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_267),
.C(n_268),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_235),
.C(n_236),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_214),
.C(n_215),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_194),
.C(n_195),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_172),
.C(n_173),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_158),
.C(n_163),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_154),
.B2(n_155),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_156),
.C(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.C(n_168),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_166),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_185),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_178),
.C(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_184),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_193),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_189),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_192),
.C(n_193),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_198),
.C(n_203),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_201),
.C(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_206),
.C(n_207),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_213),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_229),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_230),
.C(n_234),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_225),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_224),
.C(n_225),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_223),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_225),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.CI(n_228),
.CON(n_225),
.SN(n_225)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.CI(n_233),
.CON(n_230),
.SN(n_230)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_251),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_240),
.C(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_247),
.C(n_250),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_242),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.CI(n_245),
.CON(n_242),
.SN(n_242)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_258),
.C(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B1(n_265),
.B2(n_266),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_254),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_256),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_291),
.C(n_292),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_286)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_287),
.B2(n_299),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_288),
.C(n_289),
.Y(n_300)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_273),
.C(n_280),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_280),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_274),
.B(n_276),
.C(n_279),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_285),
.C(n_286),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_296),
.C(n_298),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_322),
.B2(n_323),
.Y(n_301)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_313),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_313),
.C(n_322),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_308),
.C(n_309),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_316),
.C(n_317),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_328),
.C(n_339),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_339),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_345),
.C(n_347),
.Y(n_348)
);


endmodule