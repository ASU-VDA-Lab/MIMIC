module fake_netlist_1_10415_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
AND2x4_ASAP7_75t_L g3 ( .A(n_0), .B(n_2), .Y(n_3) );
INVx1_ASAP7_75t_SL g4 ( .A(n_2), .Y(n_4) );
A2O1A1Ixp33_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .C(n_2), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
AOI22xp33_ASAP7_75t_L g7 ( .A1(n_6), .A2(n_3), .B1(n_4), .B2(n_0), .Y(n_7) );
INVxp67_ASAP7_75t_SL g8 ( .A(n_6), .Y(n_8) );
AOI222xp33_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_1), .B1(n_3), .B2(n_4), .C1(n_5), .C2(n_8), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
AOI21xp33_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_10), .B(n_8), .Y(n_12) );
endmodule