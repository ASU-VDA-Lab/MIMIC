module real_jpeg_26142_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_25),
.B1(n_43),
.B2(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_4),
.A2(n_20),
.B1(n_44),
.B2(n_56),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_121)
);

INVx8_ASAP7_75t_SL g78 ( 
.A(n_5),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_24),
.C(n_25),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_20),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_8),
.B(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_8),
.A2(n_25),
.B1(n_43),
.B2(n_57),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_8),
.B(n_30),
.C(n_47),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_8),
.A2(n_36),
.B(n_106),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_10),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_20),
.B1(n_39),
.B2(n_56),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_25),
.B1(n_39),
.B2(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_94),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_65),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_17),
.B(n_65),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.C(n_53),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_18),
.B(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_23),
.Y(n_19)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_20),
.A2(n_24),
.B1(n_56),
.B2(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_20),
.A2(n_56),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_25),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_25),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_28),
.A2(n_36),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_29),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_29),
.B(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_34),
.A2(n_121),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_36),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_40),
.A2(n_53),
.B1(n_54),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_40),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_42),
.A2(n_49),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_45),
.B(n_92),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_49),
.B(n_57),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_62),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_57),
.B(n_134),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_69),
.B(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_85),
.B2(n_86),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B(n_91),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_91),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_140),
.B(n_145),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_116),
.B(n_139),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_110),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_110),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_102),
.C(n_104),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_126),
.B(n_138),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_124),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_131),
.B(n_137),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_144),
.Y(n_145)
);


endmodule