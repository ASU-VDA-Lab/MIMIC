module real_aes_15744_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_883, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_883;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_119;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
AND2x4_ASAP7_75t_L g845 ( .A(n_0), .B(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_1), .A2(n_33), .B1(n_124), .B2(n_126), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_2), .A2(n_10), .B1(n_167), .B2(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g846 ( .A(n_3), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_4), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_5), .A2(n_11), .B1(n_169), .B2(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g815 ( .A(n_6), .Y(n_815) );
OR2x2_ASAP7_75t_L g825 ( .A(n_7), .B(n_30), .Y(n_825) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_8), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_9), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_12), .B(n_168), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_13), .A2(n_96), .B1(n_167), .B2(n_186), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_14), .A2(n_29), .B1(n_200), .B2(n_201), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_15), .B(n_168), .Y(n_241) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_16), .A2(n_46), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_17), .B(n_544), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_18), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_19), .A2(n_37), .B1(n_132), .B2(n_134), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_20), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_21), .A2(n_39), .B1(n_859), .B2(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g860 ( .A(n_21), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_22), .A2(n_44), .B1(n_134), .B2(n_167), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_23), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_24), .B(n_200), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_25), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_26), .B(n_224), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_27), .B(n_138), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_28), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_31), .A2(n_80), .B1(n_124), .B2(n_149), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_32), .A2(n_36), .B1(n_124), .B2(n_171), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_34), .A2(n_49), .B1(n_167), .B2(n_189), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_35), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_38), .Y(n_865) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_39), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g859 ( .A(n_39), .Y(n_859) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_40), .B(n_168), .Y(n_530) );
INVx2_ASAP7_75t_L g820 ( .A(n_41), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_42), .B(n_136), .Y(n_539) );
BUFx3_ASAP7_75t_L g823 ( .A(n_43), .Y(n_823) );
INVx1_ASAP7_75t_L g851 ( .A(n_43), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_45), .B(n_495), .Y(n_546) );
AND2x2_ASAP7_75t_L g494 ( .A(n_47), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_48), .B(n_202), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_50), .B(n_224), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_51), .B(n_132), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_52), .A2(n_68), .B1(n_132), .B2(n_189), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_53), .A2(n_71), .B1(n_124), .B2(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_54), .B(n_516), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_55), .A2(n_152), .B(n_471), .C(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_56), .A2(n_93), .B1(n_167), .B2(n_169), .Y(n_166) );
AND2x4_ASAP7_75t_L g120 ( .A(n_57), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g141 ( .A(n_58), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_59), .A2(n_60), .B1(n_134), .B2(n_205), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_61), .B(n_138), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_62), .B(n_495), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_63), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_64), .B(n_134), .Y(n_533) );
INVx1_ASAP7_75t_L g121 ( .A(n_65), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_66), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_67), .B(n_138), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_69), .B(n_124), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_70), .B(n_126), .C(n_136), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_72), .B(n_124), .Y(n_469) );
INVx2_ASAP7_75t_L g130 ( .A(n_73), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_74), .B(n_154), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_75), .B(n_168), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_76), .B(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_77), .A2(n_92), .B1(n_134), .B2(n_152), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_78), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_79), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_81), .A2(n_86), .B1(n_224), .B2(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_82), .B(n_168), .Y(n_563) );
NAND2xp33_ASAP7_75t_SL g504 ( .A(n_83), .B(n_133), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_84), .B(n_187), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_85), .B(n_138), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_87), .Y(n_228) );
INVx1_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_88), .B(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_89), .B(n_829), .Y(n_828) );
NAND2xp33_ASAP7_75t_L g244 ( .A(n_90), .B(n_168), .Y(n_244) );
NAND2xp33_ASAP7_75t_L g470 ( .A(n_91), .B(n_133), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_94), .B(n_495), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_95), .B(n_133), .C(n_154), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_97), .B(n_124), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_98), .B(n_224), .Y(n_514) );
OAI32xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_836), .A3(n_871), .B1(n_876), .B2(n_883), .Y(n_99) );
NAND3xp33_ASAP7_75t_L g100 ( .A(n_101), .B(n_826), .C(n_828), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_813), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2xp33_ASAP7_75t_L g826 ( .A(n_103), .B(n_827), .Y(n_826) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_455), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_110), .Y(n_104) );
INVx8_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx12f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g834 ( .A(n_108), .B(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g812 ( .A(n_109), .Y(n_812) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1p5_ASAP7_75t_L g111 ( .A(n_112), .B(n_365), .Y(n_111) );
NAND4xp75_ASAP7_75t_L g112 ( .A(n_113), .B(n_310), .C(n_330), .D(n_346), .Y(n_112) );
NOR2x1p5_ASAP7_75t_SL g113 ( .A(n_114), .B(n_280), .Y(n_113) );
NAND4xp75_ASAP7_75t_L g114 ( .A(n_115), .B(n_216), .C(n_257), .D(n_266), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_177), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_144), .Y(n_116) );
AND2x4_ASAP7_75t_L g390 ( .A(n_117), .B(n_317), .Y(n_390) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_118), .Y(n_233) );
INVx2_ASAP7_75t_L g251 ( .A(n_118), .Y(n_251) );
AND2x2_ASAP7_75t_L g274 ( .A(n_118), .B(n_236), .Y(n_274) );
OR2x2_ASAP7_75t_L g329 ( .A(n_118), .B(n_145), .Y(n_329) );
AO31x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_122), .A3(n_137), .B(n_142), .Y(n_118) );
INVx2_ASAP7_75t_L g174 ( .A(n_119), .Y(n_174) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_119), .A2(n_146), .A3(n_198), .B(n_206), .Y(n_197) );
AO31x2_ASAP7_75t_L g220 ( .A1(n_119), .A2(n_163), .A3(n_221), .B(n_227), .Y(n_220) );
AO31x2_ASAP7_75t_L g550 ( .A1(n_119), .A2(n_158), .A3(n_551), .B(n_555), .Y(n_550) );
BUFx10_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g156 ( .A(n_120), .Y(n_156) );
BUFx10_ASAP7_75t_L g480 ( .A(n_120), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B1(n_131), .B2(n_135), .Y(n_122) );
INVx1_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
INVx4_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
INVx1_ASAP7_75t_L g189 ( .A(n_124), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_124), .A2(n_134), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_125), .Y(n_126) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_125), .Y(n_134) );
INVx2_ASAP7_75t_L g150 ( .A(n_125), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
INVx1_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx1_ASAP7_75t_L g202 ( .A(n_125), .Y(n_202) );
INVx1_ASAP7_75t_L g205 ( .A(n_125), .Y(n_205) );
INVx1_ASAP7_75t_L g225 ( .A(n_125), .Y(n_225) );
INVx2_ASAP7_75t_L g516 ( .A(n_126), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_127), .A2(n_135), .B1(n_185), .B2(n_188), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_127), .A2(n_135), .B1(n_199), .B2(n_203), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_127), .A2(n_135), .B1(n_212), .B2(n_213), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_127), .B(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_127), .A2(n_135), .B1(n_552), .B2(n_554), .Y(n_551) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g517 ( .A(n_128), .Y(n_517) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g476 ( .A(n_129), .Y(n_476) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx8_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
INVx1_ASAP7_75t_L g472 ( .A(n_130), .Y(n_472) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_134), .A2(n_539), .B(n_540), .Y(n_538) );
INVx2_ASAP7_75t_L g553 ( .A(n_134), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_135), .A2(n_148), .B1(n_151), .B2(n_153), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_135), .A2(n_166), .B1(n_170), .B2(n_172), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_135), .A2(n_172), .B1(n_222), .B2(n_226), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_135), .A2(n_243), .B(n_244), .Y(n_242) );
INVx6_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_136), .A2(n_171), .B(n_240), .C(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_136), .A2(n_532), .B(n_533), .Y(n_531) );
O2A1O1Ixp5_ASAP7_75t_L g561 ( .A1(n_136), .A2(n_186), .B(n_562), .C(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_139), .B(n_143), .Y(n_142) );
BUFx3_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_139), .B(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_139), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_SL g237 ( .A(n_139), .Y(n_237) );
AND2x4_ASAP7_75t_SL g479 ( .A(n_139), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g497 ( .A(n_139), .Y(n_497) );
INVx2_ASAP7_75t_L g526 ( .A(n_139), .Y(n_526) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g159 ( .A(n_140), .Y(n_159) );
AND2x2_ASAP7_75t_L g247 ( .A(n_144), .B(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g397 ( .A(n_144), .B(n_274), .Y(n_397) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_161), .Y(n_144) );
OR2x2_ASAP7_75t_L g234 ( .A(n_145), .B(n_235), .Y(n_234) );
BUFx2_ASAP7_75t_L g265 ( .A(n_145), .Y(n_265) );
AND2x2_ASAP7_75t_L g271 ( .A(n_145), .B(n_162), .Y(n_271) );
INVx1_ASAP7_75t_L g289 ( .A(n_145), .Y(n_289) );
INVx2_ASAP7_75t_L g318 ( .A(n_145), .Y(n_318) );
AO31x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .A3(n_155), .B(n_157), .Y(n_145) );
INVx2_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_150), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g477 ( .A(n_152), .Y(n_477) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_SL g172 ( .A(n_154), .Y(n_172) );
INVx1_ASAP7_75t_L g545 ( .A(n_154), .Y(n_545) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_155), .A2(n_190), .A3(n_211), .B(n_214), .Y(n_210) );
INVx2_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_SL g245 ( .A(n_156), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
INVx2_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
NOR2xp33_ASAP7_75t_SL g227 ( .A(n_158), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g164 ( .A(n_159), .Y(n_164) );
INVx2_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
INVx3_ASAP7_75t_L g294 ( .A(n_161), .Y(n_294) );
INVx2_ASAP7_75t_L g299 ( .A(n_161), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_161), .B(n_250), .Y(n_304) );
AND2x2_ASAP7_75t_L g327 ( .A(n_161), .B(n_306), .Y(n_327) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_161), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_161), .B(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_L g316 ( .A(n_162), .Y(n_316) );
AND2x2_ASAP7_75t_L g364 ( .A(n_162), .B(n_318), .Y(n_364) );
AO31x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .A3(n_173), .B(n_175), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_164), .B(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_168), .A2(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g544 ( .A(n_168), .Y(n_544) );
AO31x2_ASAP7_75t_L g183 ( .A1(n_173), .A2(n_184), .A3(n_190), .B(n_192), .Y(n_183) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp67_ASAP7_75t_SL g485 ( .A(n_174), .B(n_191), .Y(n_485) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_195), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_179), .B(n_308), .Y(n_355) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_180), .B(n_308), .Y(n_352) );
INVx1_ASAP7_75t_L g453 ( .A(n_180), .Y(n_453) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g403 ( .A(n_181), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g256 ( .A(n_182), .Y(n_256) );
OR2x2_ASAP7_75t_L g337 ( .A(n_182), .B(n_209), .Y(n_337) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g279 ( .A(n_183), .Y(n_279) );
AND2x4_ASAP7_75t_L g285 ( .A(n_183), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_194), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g495 ( .A(n_194), .Y(n_495) );
INVx2_ASAP7_75t_L g518 ( .A(n_194), .Y(n_518) );
AOI32xp33_ASAP7_75t_L g423 ( .A1(n_195), .A2(n_326), .A3(n_424), .B1(n_426), .B2(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g372 ( .A(n_196), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_208), .Y(n_196) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_197), .Y(n_218) );
OR2x2_ASAP7_75t_L g254 ( .A(n_197), .B(n_210), .Y(n_254) );
INVx1_ASAP7_75t_L g269 ( .A(n_197), .Y(n_269) );
AND2x2_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g284 ( .A(n_197), .Y(n_284) );
INVx2_ASAP7_75t_L g309 ( .A(n_197), .Y(n_309) );
AND2x2_ASAP7_75t_L g428 ( .A(n_197), .B(n_220), .Y(n_428) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_208), .B(n_261), .Y(n_348) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g219 ( .A(n_210), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
INVx2_ASAP7_75t_L g286 ( .A(n_210), .Y(n_286) );
AND2x4_ASAP7_75t_L g308 ( .A(n_210), .B(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_210), .Y(n_400) );
AOI22x1_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_229), .B1(n_247), .B2(n_252), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
NAND4xp25_ASAP7_75t_L g377 ( .A(n_219), .B(n_378), .C(n_379), .D(n_380), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_219), .B(n_278), .Y(n_408) );
INVx4_ASAP7_75t_SL g261 ( .A(n_220), .Y(n_261) );
BUFx2_ASAP7_75t_L g324 ( .A(n_220), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_220), .B(n_269), .Y(n_387) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g349 ( .A(n_231), .B(n_298), .Y(n_349) );
NOR2x1_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x4_ASAP7_75t_L g272 ( .A(n_235), .B(n_250), .Y(n_272) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_236), .B(n_251), .Y(n_296) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_236) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_291) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_242), .B(n_245), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_248), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g314 ( .A(n_248), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g353 ( .A(n_249), .B(n_271), .Y(n_353) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g396 ( .A(n_251), .B(n_306), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_252), .A2(n_369), .B1(n_371), .B2(n_374), .C(n_376), .Y(n_368) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g262 ( .A(n_254), .Y(n_262) );
OR2x2_ASAP7_75t_L g362 ( .A(n_254), .B(n_301), .Y(n_362) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_263), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_258), .A2(n_384), .B1(n_388), .B2(n_391), .Y(n_383) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
AND2x4_ASAP7_75t_L g307 ( .A(n_259), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g419 ( .A(n_259), .B(n_337), .Y(n_419) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g267 ( .A(n_261), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g283 ( .A(n_261), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g342 ( .A(n_261), .B(n_279), .Y(n_342) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_261), .Y(n_359) );
INVx1_ASAP7_75t_L g373 ( .A(n_261), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_261), .B(n_286), .Y(n_416) );
AND2x4_ASAP7_75t_L g323 ( .A(n_262), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_265), .B(n_306), .Y(n_305) );
NAND2x1_ASAP7_75t_L g425 ( .A(n_265), .B(n_327), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B1(n_273), .B2(n_275), .Y(n_266) );
AND2x2_ASAP7_75t_L g292 ( .A(n_267), .B(n_285), .Y(n_292) );
INVx1_ASAP7_75t_L g333 ( .A(n_267), .Y(n_333) );
AND2x2_ASAP7_75t_L g440 ( .A(n_267), .B(n_301), .Y(n_440) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_SL g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_L g273 ( .A(n_271), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g413 ( .A(n_271), .Y(n_413) );
AND2x2_ASAP7_75t_L g430 ( .A(n_271), .B(n_290), .Y(n_430) );
AND2x2_ASAP7_75t_L g446 ( .A(n_271), .B(n_396), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_272), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g369 ( .A(n_272), .B(n_370), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_272), .A2(n_362), .B1(n_377), .B2(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g332 ( .A(n_274), .Y(n_332) );
AND2x2_ASAP7_75t_L g363 ( .A(n_274), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_274), .B(n_370), .Y(n_392) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g398 ( .A(n_278), .B(n_399), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_278), .A2(n_302), .B1(n_407), .B2(n_409), .Y(n_406) );
INVx3_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
AND2x2_ASAP7_75t_L g433 ( .A(n_279), .B(n_286), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_297), .Y(n_280) );
AOI32xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_287), .A3(n_290), .B1(n_292), .B2(n_293), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_284), .Y(n_379) );
INVx1_ASAP7_75t_L g404 ( .A(n_284), .Y(n_404) );
INVx3_ASAP7_75t_L g360 ( .A(n_285), .Y(n_360) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_288), .A2(n_436), .B1(n_437), .B2(n_438), .C(n_439), .Y(n_435) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g412 ( .A(n_290), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g448 ( .A(n_290), .B(n_409), .Y(n_448) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g306 ( .A(n_291), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_293), .B(n_321), .Y(n_320) );
AO22x1_ASAP7_75t_L g350 ( .A1(n_293), .A2(n_351), .B1(n_353), .B2(n_354), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_293), .B(n_321), .Y(n_454) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g370 ( .A(n_294), .Y(n_370) );
INVx1_ASAP7_75t_L g380 ( .A(n_294), .Y(n_380) );
AND2x2_ASAP7_75t_L g300 ( .A(n_295), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_296), .Y(n_382) );
INVx1_ASAP7_75t_L g422 ( .A(n_296), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_300), .B(n_302), .C(n_307), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NOR2x1p5_ASAP7_75t_L g409 ( .A(n_299), .B(n_329), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_300), .B(n_359), .Y(n_436) );
AOI31xp33_ASAP7_75t_L g319 ( .A1(n_301), .A2(n_320), .A3(n_322), .B(n_325), .Y(n_319) );
INVx4_ASAP7_75t_L g378 ( .A(n_301), .Y(n_378) );
OR2x2_ASAP7_75t_L g415 ( .A(n_301), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x4_ASAP7_75t_L g317 ( .A(n_306), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_308), .Y(n_313) );
AND2x2_ASAP7_75t_L g344 ( .A(n_308), .B(n_342), .Y(n_344) );
NOR2xp67_ASAP7_75t_L g310 ( .A(n_311), .B(n_319), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g437 ( .A(n_314), .Y(n_437) );
INVx1_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g375 ( .A(n_316), .Y(n_375) );
AND2x2_ASAP7_75t_L g374 ( .A(n_317), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI322xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .A3(n_334), .B1(n_338), .B2(n_341), .C1(n_343), .C2(n_345), .Y(n_331) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI211x1_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B(n_350), .C(n_356), .Y(n_346) );
INVx1_ASAP7_75t_L g451 ( .A(n_347), .Y(n_451) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g405 ( .A(n_349), .Y(n_405) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_361), .B(n_363), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g426 ( .A(n_360), .Y(n_426) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_364), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_434), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_401), .C(n_417), .Y(n_366) );
NAND3xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_383), .C(n_393), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_370), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_374), .A2(n_430), .B(n_431), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_378), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_378), .B(n_428), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_379), .B(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_380), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_390), .A2(n_440), .B(n_441), .Y(n_439) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B(n_406), .C(n_410), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_412), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_416), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B(n_423), .C(n_429), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_428), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g449 ( .A(n_428), .Y(n_449) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g445 ( .A(n_433), .Y(n_445) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_443), .C(n_450), .Y(n_434) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI21xp33_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_447), .B(n_449), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI21xp33_ASAP7_75t_R g450 ( .A1(n_451), .A2(n_452), .B(n_454), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_811), .Y(n_455) );
INVx1_ASAP7_75t_L g862 ( .A(n_457), .Y(n_862) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_691), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_599), .C(n_650), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_520), .B(n_568), .C(n_586), .Y(n_459) );
NAND3x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_481), .C(n_506), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g659 ( .A(n_462), .B(n_638), .Y(n_659) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND3x2_ASAP7_75t_L g579 ( .A(n_463), .B(n_580), .C(n_584), .Y(n_579) );
AND2x2_ASAP7_75t_L g614 ( .A(n_463), .B(n_598), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_463), .B(n_616), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_463), .B(n_584), .Y(n_761) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g663 ( .A(n_464), .B(n_584), .Y(n_663) );
AND2x2_ASAP7_75t_L g674 ( .A(n_464), .B(n_628), .Y(n_674) );
BUFx2_ASAP7_75t_L g680 ( .A(n_464), .Y(n_680) );
NAND2x1_ASAP7_75t_L g696 ( .A(n_464), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g702 ( .A(n_464), .B(n_703), .Y(n_702) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g596 ( .A(n_465), .Y(n_596) );
AND2x2_ASAP7_75t_L g627 ( .A(n_465), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g647 ( .A(n_465), .B(n_583), .Y(n_647) );
INVx1_ASAP7_75t_L g718 ( .A(n_465), .Y(n_718) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
OAI21x1_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_473), .B(n_479), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_471), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_471), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_471), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_471), .A2(n_529), .B(n_530), .Y(n_528) );
BUFx4f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_476), .B1(n_477), .B2(n_478), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_475), .A2(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
OAI21x1_ASAP7_75t_L g498 ( .A1(n_480), .A2(n_499), .B(n_502), .Y(n_498) );
OAI21x1_ASAP7_75t_L g509 ( .A1(n_480), .A2(n_510), .B(n_513), .Y(n_509) );
OAI21x1_ASAP7_75t_L g527 ( .A1(n_480), .A2(n_528), .B(n_531), .Y(n_527) );
OAI21x1_ASAP7_75t_L g537 ( .A1(n_480), .A2(n_538), .B(n_541), .Y(n_537) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_480), .A2(n_561), .B(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x6_ASAP7_75t_L g695 ( .A(n_482), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g597 ( .A(n_483), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_483), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
INVx2_ASAP7_75t_L g585 ( .A(n_484), .Y(n_585) );
INVx1_ASAP7_75t_L g639 ( .A(n_484), .Y(n_639) );
AOI21x1_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_494), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
INVx2_ASAP7_75t_L g617 ( .A(n_496), .Y(n_617) );
OAI21x1_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_505), .Y(n_496) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_507), .A2(n_799), .B(n_803), .Y(n_798) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g638 ( .A(n_508), .B(n_639), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_518), .B(n_519), .Y(n_508) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_509), .A2(n_518), .B(n_519), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_517), .Y(n_513) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_518), .A2(n_560), .B(n_567), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_518), .A2(n_560), .B(n_567), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_547), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_522), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2xp67_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
INVx3_ASAP7_75t_L g576 ( .A(n_524), .Y(n_576) );
AND2x2_ASAP7_75t_L g723 ( .A(n_524), .B(n_536), .Y(n_723) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g612 ( .A(n_525), .Y(n_612) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_534), .Y(n_525) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_526), .A2(n_537), .B(n_546), .Y(n_536) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_526), .A2(n_527), .B(n_534), .Y(n_591) );
OA21x2_ASAP7_75t_L g594 ( .A1(n_526), .A2(n_537), .B(n_546), .Y(n_594) );
AND2x4_ASAP7_75t_L g577 ( .A(n_535), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g636 ( .A(n_536), .Y(n_636) );
AND2x2_ASAP7_75t_L g653 ( .A(n_536), .B(n_550), .Y(n_653) );
AND2x2_ASAP7_75t_L g765 ( .A(n_536), .B(n_642), .Y(n_765) );
AND2x2_ASAP7_75t_L g787 ( .A(n_536), .B(n_558), .Y(n_787) );
AOI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_545), .Y(n_541) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_549), .B(n_557), .Y(n_548) );
INVx1_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_549), .B(n_797), .Y(n_796) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g578 ( .A(n_550), .Y(n_578) );
OR2x2_ASAP7_75t_L g593 ( .A(n_550), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g611 ( .A(n_550), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g665 ( .A(n_550), .B(n_591), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_550), .B(n_594), .Y(n_707) );
OR2x2_ASAP7_75t_L g777 ( .A(n_550), .B(n_591), .Y(n_777) );
INVx1_ASAP7_75t_L g605 ( .A(n_557), .Y(n_605) );
AND2x4_ASAP7_75t_L g623 ( .A(n_557), .B(n_577), .Y(n_623) );
AND2x2_ASAP7_75t_L g769 ( .A(n_557), .B(n_611), .Y(n_769) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx3_ASAP7_75t_L g571 ( .A(n_558), .Y(n_571) );
AND2x2_ASAP7_75t_L g631 ( .A(n_558), .B(n_590), .Y(n_631) );
INVx1_ASAP7_75t_L g684 ( .A(n_558), .Y(n_684) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_558), .Y(n_722) );
AND2x2_ASAP7_75t_L g725 ( .A(n_558), .B(n_594), .Y(n_725) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_558), .Y(n_735) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B(n_579), .Y(n_568) );
AND2x2_ASAP7_75t_L g767 ( .A(n_569), .B(n_672), .Y(n_767) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g634 ( .A(n_570), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_570), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_571), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g714 ( .A(n_571), .B(n_577), .Y(n_714) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_576), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g712 ( .A(n_576), .B(n_653), .Y(n_712) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_576), .Y(n_743) );
INVx2_ASAP7_75t_L g677 ( .A(n_577), .Y(n_677) );
AND2x2_ASAP7_75t_L g806 ( .A(n_578), .B(n_591), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_579), .A2(n_661), .B1(n_662), .B2(n_664), .C(n_666), .Y(n_660) );
AND2x2_ASAP7_75t_L g601 ( .A(n_580), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g662 ( .A(n_580), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx2_ASAP7_75t_L g598 ( .A(n_581), .Y(n_598) );
OR2x2_ASAP7_75t_L g731 ( .A(n_581), .B(n_616), .Y(n_731) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g628 ( .A(n_582), .Y(n_628) );
INVxp67_ASAP7_75t_L g658 ( .A(n_583), .Y(n_658) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g602 ( .A(n_585), .Y(n_602) );
AND2x2_ASAP7_75t_L g615 ( .A(n_585), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g622 ( .A(n_585), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_595), .Y(n_586) );
AND2x2_ASAP7_75t_L g745 ( .A(n_587), .B(n_746), .Y(n_745) );
AND2x4_ASAP7_75t_L g587 ( .A(n_588), .B(n_592), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g672 ( .A(n_589), .B(n_653), .Y(n_672) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_589), .Y(n_802) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g630 ( .A(n_592), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g780 ( .A(n_592), .Y(n_780) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g668 ( .A(n_593), .Y(n_668) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_593), .Y(n_742) );
AND2x2_ASAP7_75t_L g641 ( .A(n_594), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_595), .B(n_767), .Y(n_766) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g637 ( .A(n_596), .B(n_638), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_597), .A2(n_619), .B(n_623), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g599 ( .A(n_600), .B(n_618), .C(n_624), .D(n_632), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B(n_608), .Y(n_600) );
INVx2_ASAP7_75t_L g689 ( .A(n_602), .Y(n_689) );
AND2x2_ASAP7_75t_L g700 ( .A(n_602), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g710 ( .A(n_602), .B(n_627), .Y(n_710) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g786 ( .A(n_607), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_613), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI33xp33_ASAP7_75t_L g756 ( .A1(n_610), .A2(n_647), .A3(n_757), .B1(n_759), .B2(n_762), .B3(n_763), .Y(n_756) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g789 ( .A(n_611), .B(n_641), .Y(n_789) );
BUFx2_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_615), .B(n_627), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_616), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_617), .Y(n_670) );
INVx1_ASAP7_75t_L g703 ( .A(n_617), .Y(n_703) );
AND2x2_ASAP7_75t_L g717 ( .A(n_617), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g688 ( .A(n_620), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g740 ( .A(n_620), .Y(n_740) );
INVx1_ASAP7_75t_L g750 ( .A(n_621), .Y(n_750) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g626 ( .A(n_622), .Y(n_626) );
INVx1_ASAP7_75t_L g732 ( .A(n_622), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_629), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
OR2x2_ASAP7_75t_L g715 ( .A(n_626), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g686 ( .A(n_627), .B(n_670), .Y(n_686) );
AND2x2_ASAP7_75t_L g649 ( .A(n_628), .B(n_639), .Y(n_649) );
INVx2_ASAP7_75t_L g697 ( .A(n_628), .Y(n_697) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g690 ( .A(n_631), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_637), .B1(n_640), .B2(n_645), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_635), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_637), .A2(n_720), .B1(n_724), .B2(n_726), .C(n_728), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_638), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g774 ( .A(n_638), .Y(n_774) );
AND2x2_ASAP7_75t_L g793 ( .A(n_638), .B(n_717), .Y(n_793) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g762 ( .A(n_641), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_641), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g748 ( .A(n_642), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_643), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g736 ( .A(n_643), .B(n_677), .Y(n_736) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_645), .A2(n_791), .B1(n_793), .B2(n_794), .Y(n_790) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
OR2x2_ASAP7_75t_L g807 ( .A(n_648), .B(n_702), .Y(n_807) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g755 ( .A(n_649), .B(n_717), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B(n_660), .C(n_675), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_653), .Y(n_661) );
AND2x2_ASAP7_75t_L g734 ( .A(n_653), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g727 ( .A(n_659), .Y(n_727) );
BUFx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_665), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g724 ( .A(n_665), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g758 ( .A(n_665), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_665), .B(n_772), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B1(n_671), .B2(n_673), .Y(n_666) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI21xp33_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_678), .B(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B1(n_687), .B2(n_690), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_683), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI211xp5_ASAP7_75t_SL g768 ( .A1(n_686), .A2(n_769), .B(n_770), .C(n_778), .Y(n_768) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g783 ( .A(n_689), .B(n_717), .Y(n_783) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_751), .C(n_781), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_719), .C(n_739), .Y(n_692) );
O2A1O1Ixp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_698), .B(n_704), .C(n_708), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp33_ASAP7_75t_SL g770 ( .A1(n_696), .A2(n_771), .B1(n_773), .B2(n_775), .Y(n_770) );
INVx1_ASAP7_75t_SL g760 ( .A(n_697), .Y(n_760) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g773 ( .A(n_702), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B1(n_713), .B2(n_715), .Y(n_708) );
NAND2xp33_ASAP7_75t_SL g726 ( .A(n_709), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g792 ( .A(n_714), .Y(n_792) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g746 ( .A(n_717), .B(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_721), .B(n_755), .Y(n_754) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g797 ( .A(n_722), .Y(n_797) );
INVx1_ASAP7_75t_L g772 ( .A(n_725), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_733), .B1(n_736), .B2(n_737), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2x1p5_ASAP7_75t_SL g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g738 ( .A(n_731), .Y(n_738) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g744 ( .A(n_735), .Y(n_744) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_745), .C(n_749), .Y(n_739) );
NOR3x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .C(n_744), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_746), .B(n_801), .Y(n_800) );
AND2x2_ASAP7_75t_L g805 ( .A(n_747), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_766), .C(n_768), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NOR2xp67_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g810 ( .A(n_779), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_790), .C(n_798), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_788), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVxp67_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVxp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVxp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx6f_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NOR2xp33_ASAP7_75t_SL g813 ( .A(n_814), .B(n_816), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_815), .B(n_816), .Y(n_827) );
CKINVDCx16_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
BUFx12f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AND2x6_ASAP7_75t_SL g818 ( .A(n_819), .B(n_821), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_820), .B(n_833), .Y(n_832) );
INVx3_ASAP7_75t_L g842 ( .A(n_820), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_820), .B(n_847), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_823), .B(n_825), .Y(n_835) );
AND2x6_ASAP7_75t_SL g848 ( .A(n_824), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx10_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_852), .B1(n_860), .B2(n_868), .Y(n_836) );
INVx8_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_839), .Y(n_838) );
OR2x6_ASAP7_75t_L g839 ( .A(n_840), .B(n_847), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
BUFx6f_ASAP7_75t_L g875 ( .A(n_842), .Y(n_875) );
OR2x4_ASAP7_75t_L g869 ( .A(n_843), .B(n_870), .Y(n_869) );
BUFx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
AND2x2_ASAP7_75t_L g880 ( .A(n_845), .B(n_881), .Y(n_880) );
INVx2_ASAP7_75t_L g854 ( .A(n_847), .Y(n_854) );
INVx3_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx4_ASAP7_75t_L g867 ( .A(n_848), .Y(n_867) );
INVx5_ASAP7_75t_L g881 ( .A(n_848), .Y(n_881) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVxp67_ASAP7_75t_SL g852 ( .A(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_SL g872 ( .A(n_853), .B(n_873), .Y(n_872) );
OAI21xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B(n_863), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B1(n_861), .B2(n_862), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NOR2xp33_ASAP7_75t_SL g864 ( .A(n_865), .B(n_866), .Y(n_864) );
BUFx12f_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx4_ASAP7_75t_SL g868 ( .A(n_869), .Y(n_868) );
INVxp67_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
CKINVDCx11_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_877), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_878), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_879), .Y(n_878) );
CKINVDCx16_ASAP7_75t_R g879 ( .A(n_880), .Y(n_879) );
endmodule