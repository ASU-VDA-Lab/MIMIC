module real_jpeg_7119_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_0),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_0),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_0),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_0),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_0),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_0),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_0),
.B(n_63),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_0),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_1),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_1),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_1),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_1),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_1),
.B(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_2),
.Y(n_271)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_2),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_2),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_2),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_3),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_4),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_4),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_4),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_4),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_5),
.B(n_59),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_5),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_5),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_5),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_5),
.B(n_282),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_5),
.B(n_414),
.Y(n_413)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g405 ( 
.A(n_6),
.Y(n_405)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_7),
.Y(n_509)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g375 ( 
.A(n_8),
.Y(n_375)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_10),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_11),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_11),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_11),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_11),
.B(n_126),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_11),
.B(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_13),
.B(n_164),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_13),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_13),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_13),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_13),
.B(n_356),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_13),
.B(n_49),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_13),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_14),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_14),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_14),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_14),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_14),
.B(n_117),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_14),
.B(n_99),
.Y(n_390)
);

AND2x6_ASAP7_75t_SL g404 ( 
.A(n_14),
.B(n_405),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_15),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_15),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_15),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_15),
.B(n_316),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_15),
.B(n_381),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_15),
.B(n_375),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_16),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_16),
.B(n_42),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_16),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_16),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_16),
.B(n_282),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_16),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_16),
.B(n_132),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_16),
.B(n_117),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_17),
.Y(n_512)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_19),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_19),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_19),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_19),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_19),
.B(n_65),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_19),
.B(n_378),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_19),
.B(n_419),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_507),
.B(n_510),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_175),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_174),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_106),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_25),
.B(n_106),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_84),
.B1(n_85),
.B2(n_105),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_26),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_55),
.C(n_72),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_27),
.A2(n_28),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_30),
.B(n_34),
.C(n_40),
.Y(n_104)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_37),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_39),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_39),
.Y(n_301)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_39),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.C(n_51),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_41),
.B(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_43),
.Y(n_218)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_145)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_48),
.B(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_50),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_54),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_55),
.A2(n_72),
.B1(n_73),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.C(n_67),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_56),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_60),
.Y(n_197)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_60),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_61),
.A2(n_62),
.B1(n_139),
.B2(n_143),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_167)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_62),
.B(n_135),
.C(n_139),
.Y(n_168)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_66),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_66),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_68),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_78),
.C(n_83),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_71),
.Y(n_345)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_83),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_79),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_104),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_95),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_94),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_100),
.Y(n_275)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_165),
.C(n_170),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_107),
.A2(n_108),
.B1(n_493),
.B2(n_494),
.Y(n_492)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_144),
.C(n_146),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_109),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_122),
.C(n_134),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_110),
.A2(n_111),
.B1(n_122),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_116),
.C(n_119),
.Y(n_169)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_122),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.C(n_129),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_123),
.B(n_129),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_125),
.B(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_128),
.Y(n_320)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_133),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_134),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_139),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_149),
.C(n_153),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_139),
.A2(n_143),
.B1(n_149),
.B2(n_150),
.Y(n_243)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_141),
.Y(n_314)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_142),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_142),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_144),
.B(n_146),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_158),
.C(n_161),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_147),
.A2(n_148),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_149),
.A2(n_150),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_149),
.B(n_211),
.C(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_152),
.Y(n_325)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_152),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_153),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_158),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_158),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_158),
.A2(n_161),
.B1(n_220),
.B2(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_219),
.C(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_161),
.Y(n_253)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_165),
.B(n_170),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_166),
.B(n_499),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_168),
.B(n_169),
.Y(n_499)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_490),
.B(n_504),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_302),
.B(n_489),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_256),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_179),
.B(n_256),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_235),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_180),
.B(n_236),
.C(n_239),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_215),
.C(n_222),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_181),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_193),
.C(n_207),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_182),
.B(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_188),
.C(n_192),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_193),
.A2(n_194),
.B1(n_207),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_203),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_195),
.B(n_203),
.Y(n_465)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_198),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_202),
.Y(n_358)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_202),
.Y(n_414)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_207),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_222),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.C(n_232),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.C(n_229),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_224),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_229),
.Y(n_268)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_231),
.B(n_232),
.Y(n_288)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_248),
.B2(n_249),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_240),
.B(n_250),
.C(n_254),
.Y(n_500)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_246),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_258),
.B(n_261),
.Y(n_485)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_263),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_286),
.C(n_289),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_265),
.B(n_478),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_276),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_266),
.A2(n_267),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_269),
.A2(n_270),
.B(n_272),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_269),
.B(n_276),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_284),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_433)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx8_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_284),
.B(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_285),
.B(n_374),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_289),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.C(n_299),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_291),
.B(n_467),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_292),
.B(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_294),
.Y(n_446)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_298),
.B(n_299),
.Y(n_467)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_483),
.B(n_488),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_470),
.B(n_482),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_452),
.B(n_469),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_426),
.B(n_451),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_395),
.B(n_425),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_366),
.B(n_394),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_347),
.B(n_365),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_327),
.B(n_346),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_321),
.B(n_326),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_318),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_315),
.Y(n_328)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_329),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_335),
.B2(n_336),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_338),
.C(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_333),
.Y(n_353)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_364),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_364),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_354),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_353),
.C(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_352),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_385),
.C(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_369),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_383),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_370),
.B(n_384),
.C(n_387),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_373),
.C(n_376),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_379),
.B1(n_380),
.B2(n_382),
.Y(n_376)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_382),
.Y(n_406)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_391),
.C(n_392),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_390),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_391),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_424),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_424),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_408),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_407),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_398),
.B(n_407),
.C(n_450),
.Y(n_449)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_406),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_404),
.Y(n_399)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_400),
.Y(n_440)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_404),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_406),
.B(n_440),
.C(n_441),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_415),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_417),
.C(n_422),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_412),
.C(n_413),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_422),
.B2(n_423),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_420),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_449),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_449),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_438),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_430),
.C(n_438),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_434),
.B2(n_435),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_461),
.C(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_442),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_443),
.C(n_448),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_447),
.B2(n_448),
.Y(n_442)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_443),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_468),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_468),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_459),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_458),
.C(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_456),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_464),
.C(n_466),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_480),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_480),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_477),
.C(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_484),
.B(n_486),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_486),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_501),
.Y(n_490)
);

OAI21xp33_ASAP7_75t_L g504 ( 
.A1(n_491),
.A2(n_505),
.B(n_506),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_495),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_495),
.Y(n_506)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_493),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.C(n_500),
.Y(n_495)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_496),
.B(n_498),
.CI(n_500),
.CON(n_502),
.SN(n_502)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_502),
.B(n_503),
.Y(n_505)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_502),
.Y(n_513)
);

BUFx12f_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_508),
.Y(n_511)
);

INVx13_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);


endmodule