module fake_ibex_2_n_129 (n_7, n_20, n_17, n_25, n_18, n_3, n_22, n_28, n_4, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_14, n_0, n_9, n_12, n_15, n_24, n_31, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_129);

input n_7;
input n_20;
input n_17;
input n_25;
input n_18;
input n_3;
input n_22;
input n_28;
input n_4;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_14;
input n_0;
input n_9;
input n_12;
input n_15;
input n_24;
input n_31;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_129;

wire n_85;
wire n_128;
wire n_84;
wire n_64;
wire n_73;
wire n_65;
wire n_103;
wire n_95;
wire n_55;
wire n_63;
wire n_98;
wire n_106;
wire n_76;
wire n_118;
wire n_67;
wire n_38;
wire n_124;
wire n_37;
wire n_110;
wire n_47;
wire n_108;
wire n_82;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_69;
wire n_75;
wire n_109;
wire n_121;
wire n_127;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_39;
wire n_62;
wire n_71;
wire n_120;
wire n_93;
wire n_122;
wire n_116;
wire n_61;
wire n_94;
wire n_42;
wire n_77;
wire n_112;
wire n_88;
wire n_44;
wire n_51;
wire n_46;
wire n_80;
wire n_49;
wire n_40;
wire n_66;
wire n_74;
wire n_90;
wire n_58;
wire n_43;
wire n_119;
wire n_33;
wire n_100;
wire n_72;
wire n_114;
wire n_34;
wire n_97;
wire n_102;
wire n_123;
wire n_52;
wire n_99;
wire n_105;
wire n_126;
wire n_111;
wire n_36;
wire n_104;
wire n_41;
wire n_45;
wire n_89;
wire n_83;
wire n_32;
wire n_53;
wire n_107;
wire n_115;
wire n_50;
wire n_92;
wire n_101;
wire n_113;
wire n_96;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_35;
wire n_56;
wire n_91;
wire n_54;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_20),
.Y(n_34)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_9),
.Y(n_35)
);

AND2x4_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_29),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx8_ASAP7_75t_SL g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_8),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_10),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_11),
.B(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_55),
.Y(n_62)
);

NOR3xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_58),
.C(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_32),
.A2(n_43),
.B1(n_54),
.B2(n_33),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_41),
.Y(n_69)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_34),
.C(n_51),
.Y(n_70)
);

NOR2x1p5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_41),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_56),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_43),
.B1(n_76),
.B2(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_72),
.B(n_73),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_65),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_70),
.B1(n_62),
.B2(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_76),
.B1(n_70),
.B2(n_67),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_64),
.B(n_63),
.C(n_61),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_R g92 ( 
.A(n_68),
.B(n_60),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_72),
.B(n_73),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_72),
.B(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_64),
.B(n_63),
.C(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AO21x2_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_94),
.B(n_93),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_83),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_92),
.B1(n_88),
.B2(n_78),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_85),
.B1(n_87),
.B2(n_97),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_106),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_98),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

BUFx2_ASAP7_75t_SL g116 ( 
.A(n_111),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_105),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_105),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_99),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_107),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_R g125 ( 
.A(n_124),
.B(n_120),
.Y(n_125)
);

AO22x2_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_121),
.B1(n_115),
.B2(n_113),
.Y(n_126)
);

OR2x6_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_119),
.Y(n_128)
);

OR2x6_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_114),
.Y(n_129)
);


endmodule