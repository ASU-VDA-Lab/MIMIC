module real_jpeg_1062_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_249;
wire n_221;
wire n_215;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_238;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_267;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_75),
.B1(n_76),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_1),
.A2(n_60),
.B1(n_62),
.B2(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_86),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_1),
.A2(n_29),
.B1(n_36),
.B2(n_86),
.Y(n_179)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_3),
.A2(n_75),
.B1(n_76),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_3),
.A2(n_60),
.B1(n_62),
.B2(n_84),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_84),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_3),
.A2(n_29),
.B1(n_36),
.B2(n_84),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_4),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_4),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_4),
.A2(n_37),
.B1(n_60),
.B2(n_62),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_5),
.B(n_130),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_5),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_5),
.A2(n_75),
.B(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_5),
.B(n_64),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_5),
.A2(n_62),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_29),
.C(n_50),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_175),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_5),
.B(n_32),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_5),
.B(n_55),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_6),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_95)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_59),
.B1(n_75),
.B2(n_76),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_59),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_59),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_11),
.A2(n_54),
.B1(n_60),
.B2(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_11),
.A2(n_29),
.B1(n_36),
.B2(n_54),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_13),
.A2(n_75),
.B1(n_76),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_13),
.A2(n_60),
.B1(n_62),
.B2(n_149),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_149),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_13),
.A2(n_29),
.B1(n_36),
.B2(n_149),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_14),
.A2(n_75),
.B1(n_76),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_14),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_14),
.A2(n_60),
.B1(n_62),
.B2(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_129),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_14),
.A2(n_29),
.B1(n_36),
.B2(n_129),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_16),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_16),
.A2(n_47),
.B1(n_60),
.B2(n_62),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_16),
.A2(n_29),
.B1(n_36),
.B2(n_47),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_16),
.A2(n_47),
.B1(n_75),
.B2(n_76),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_267),
.B1(n_289),
.B2(n_290),
.Y(n_19)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_20),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_131),
.B(n_266),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_113),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_22),
.B(n_113),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_87),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_23),
.B(n_97),
.C(n_112),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_56),
.C(n_71),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_24),
.A2(n_25),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_151)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_28),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_28),
.A2(n_32),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_28),
.A2(n_32),
.B1(n_142),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_28),
.A2(n_32),
.B1(n_179),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_28),
.A2(n_32),
.B1(n_175),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_28),
.A2(n_32),
.B1(n_229),
.B2(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_29),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_31),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_31),
.A2(n_35),
.B1(n_101),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_31),
.A2(n_101),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_31),
.A2(n_101),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_43),
.A2(n_52),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AO22x2_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_45),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_44),
.B(n_67),
.Y(n_176)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_45),
.A2(n_62),
.A3(n_65),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_45),
.B(n_217),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_55),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_48),
.A2(n_53),
.B1(n_55),
.B2(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_48),
.A2(n_55),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_48),
.A2(n_55),
.B1(n_171),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_48),
.A2(n_55),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_48),
.A2(n_55),
.B1(n_199),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_48),
.A2(n_55),
.B(n_95),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_52),
.A2(n_122),
.B1(n_170),
.B2(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_71),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_58),
.A2(n_64),
.B1(n_91),
.B2(n_126),
.Y(n_125)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_62),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_60),
.B(n_78),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_60),
.B(n_175),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_76),
.A3(n_79),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_63),
.A2(n_70),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_63),
.A2(n_70),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_63),
.A2(n_70),
.B1(n_145),
.B2(n_161),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_63),
.A2(n_70),
.B1(n_160),
.B2(n_208),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_64),
.A2(n_91),
.B1(n_92),
.B2(n_282),
.Y(n_281)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_81),
.B1(n_82),
.B2(n_85),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_81),
.B1(n_85),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_81),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_72),
.A2(n_81),
.B1(n_148),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_72),
.A2(n_81),
.B1(n_110),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_83),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_81),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B1(n_98),
.B2(n_112),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B(n_96),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_93),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_96),
.A2(n_273),
.B1(n_285),
.B2(n_286),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_96),
.Y(n_285)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_105),
.B1(n_106),
.B2(n_111),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_107),
.A2(n_109),
.B(n_111),
.Y(n_271)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_118),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.C(n_127),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_120),
.B(n_123),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_127),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_154),
.B(n_265),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_152),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_133),
.B(n_152),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_151),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_134),
.B(n_151),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_136),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.C(n_147),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_137),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_141),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_144),
.B(n_147),
.Y(n_255)
);

AOI31xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_249),
.A3(n_258),
.B(n_262),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_194),
.B(n_248),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_181),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_157),
.B(n_181),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_168),
.C(n_172),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_158),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_163),
.C(n_167),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_168),
.B(n_172),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_183),
.B(n_184),
.C(n_185),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_189),
.C(n_193),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_243),
.B(n_247),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_212),
.B(n_242),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_204),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_201),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_207),
.C(n_210),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_223),
.B(n_241),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_235),
.B(n_240),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_230),
.B(n_234),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_246),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_253),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_257),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_267),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_288),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_287),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_287),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);


endmodule