module fake_jpeg_17103_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_62),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_49),
.B1(n_42),
.B2(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_70),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_47),
.B1(n_40),
.B2(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_38),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_83),
.Y(n_85)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_82),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_89),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_43),
.B1(n_71),
.B2(n_6),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_90),
.B1(n_13),
.B2(n_14),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_3),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_20),
.B1(n_36),
.B2(n_7),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_43),
.B(n_6),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_4),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_11),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_98),
.B(n_99),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_76),
.C(n_84),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_101),
.C(n_90),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_88),
.C(n_94),
.Y(n_103)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_109),
.B(n_110),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_106),
.C(n_16),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_112),
.B(n_108),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_21),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_31),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_32),
.Y(n_120)
);


endmodule