module fake_jpeg_20032_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_28),
.B1(n_23),
.B2(n_37),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_18),
.B1(n_27),
.B2(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_75),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_71),
.Y(n_96)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_18),
.B1(n_37),
.B2(n_28),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_35),
.B1(n_31),
.B2(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_73),
.Y(n_97)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_18),
.B1(n_37),
.B2(n_21),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_30),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_99),
.B1(n_72),
.B2(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_81),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_93),
.B1(n_98),
.B2(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_83),
.A2(n_109),
.B1(n_103),
.B2(n_84),
.Y(n_135)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_21),
.B1(n_19),
.B2(n_36),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_89),
.A2(n_97),
.B1(n_100),
.B2(n_102),
.Y(n_151)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_27),
.B1(n_32),
.B2(n_35),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_103),
.Y(n_130)
);

BUFx2_ASAP7_75t_SL g101 ( 
.A(n_68),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_68),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_104),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_55),
.A2(n_29),
.B1(n_34),
.B2(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_16),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_107),
.Y(n_147)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_60),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_44),
.A3(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_66),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_20),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_16),
.C(n_34),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_112),
.B1(n_108),
.B2(n_92),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_14),
.B(n_13),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_15),
.C(n_14),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_114),
.B(n_96),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_125),
.B(n_128),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_30),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_70),
.B1(n_69),
.B2(n_66),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_30),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_146),
.B1(n_1),
.B2(n_2),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_83),
.A2(n_80),
.B1(n_92),
.B2(n_93),
.Y(n_146)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_81),
.B1(n_76),
.B2(n_90),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_155),
.Y(n_203)
);

OAI211xp5_ASAP7_75t_L g217 ( 
.A1(n_153),
.A2(n_13),
.B(n_10),
.C(n_9),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_107),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_90),
.B1(n_91),
.B2(n_76),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_173),
.B1(n_184),
.B2(n_126),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_135),
.B1(n_118),
.B2(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_178),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_99),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_136),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_99),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_165),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_16),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_128),
.A2(n_26),
.B1(n_34),
.B2(n_29),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_117),
.A2(n_115),
.B1(n_110),
.B2(n_34),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_16),
.B(n_33),
.C(n_29),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_129),
.B(n_142),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_13),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_33),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_0),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_0),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_16),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_185),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_201),
.B(n_214),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_160),
.B1(n_172),
.B2(n_174),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_118),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_194),
.B(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_199),
.B1(n_208),
.B2(n_209),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_140),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_149),
.B1(n_145),
.B2(n_150),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_141),
.B(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_140),
.B1(n_144),
.B2(n_126),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_144),
.B1(n_142),
.B2(n_134),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_217),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_154),
.B(n_148),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_165),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_174),
.A2(n_139),
.B(n_119),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_177),
.B(n_179),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_155),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_225),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_192),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_158),
.B1(n_160),
.B2(n_167),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_212),
.B1(n_201),
.B2(n_215),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_237),
.B(n_239),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_180),
.B1(n_163),
.B2(n_162),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_228),
.A2(n_230),
.B1(n_243),
.B2(n_5),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_163),
.B1(n_162),
.B2(n_176),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_200),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_232),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_200),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_139),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_186),
.A2(n_153),
.B1(n_170),
.B2(n_9),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_186),
.B(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_170),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_8),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_2),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_194),
.A2(n_203),
.B(n_215),
.C(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_1),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_1),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_242),
.B1(n_191),
.B2(n_211),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_187),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_248),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_192),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_258),
.B1(n_242),
.B2(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_261),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_196),
.B1(n_206),
.B2(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

XOR2x2_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_213),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_259),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_189),
.B1(n_199),
.B2(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_237),
.A2(n_190),
.B1(n_197),
.B2(n_5),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_8),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_2),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_241),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_221),
.B(n_6),
.CI(n_3),
.CON(n_262),
.SN(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_224),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_235),
.C(n_219),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_273),
.C(n_259),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_268),
.B(n_258),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_240),
.B1(n_264),
.B2(n_234),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_219),
.C(n_229),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_232),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_274),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_226),
.B1(n_255),
.B2(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_268),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_227),
.B1(n_218),
.B2(n_239),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_281),
.B1(n_263),
.B2(n_262),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_257),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_283),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_230),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_222),
.B(n_260),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_231),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_218),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_289),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_244),
.B(n_253),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_284),
.B(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_293),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_244),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_295),
.C(n_280),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_282),
.A2(n_249),
.B1(n_222),
.B2(n_225),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_6),
.C(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_270),
.B(n_281),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_297),
.B(n_265),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_292),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_284),
.B(n_275),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_315),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_298),
.B(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_314),
.Y(n_319)
);

OAI211xp5_ASAP7_75t_SL g314 ( 
.A1(n_304),
.A2(n_287),
.B(n_293),
.C(n_279),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_271),
.B1(n_279),
.B2(n_291),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_307),
.B1(n_266),
.B2(n_314),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_308),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_322),
.B(n_317),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_305),
.C(n_280),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_318),
.B(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

NAND2x1_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_302),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_328),
.Y(n_329)
);

AOI21x1_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_323),
.B(n_265),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_289),
.C(n_269),
.Y(n_331)
);


endmodule