module fake_jpeg_27899_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_33),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_81),
.Y(n_85)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_62),
.B1(n_52),
.B2(n_61),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_66),
.C(n_65),
.Y(n_97)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_94),
.Y(n_96)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_64),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_69),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_75),
.B(n_74),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_58),
.B1(n_53),
.B2(n_70),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_60),
.B1(n_59),
.B2(n_73),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_89),
.B1(n_68),
.B2(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_54),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_84),
.B1(n_87),
.B2(n_66),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_115),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_23),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_117),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_63),
.B1(n_56),
.B2(n_55),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_119),
.B1(n_67),
.B2(n_53),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_95),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_70),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_5),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_128),
.B1(n_130),
.B2(n_132),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_19),
.B1(n_46),
.B2(n_45),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_21),
.B(n_28),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_17),
.B1(n_39),
.B2(n_37),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_15),
.C(n_30),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_2),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_113),
.B1(n_112),
.B2(n_109),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_142),
.B1(n_143),
.B2(n_10),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_141),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_137),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_125),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_4),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_6),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_6),
.B(n_8),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_142),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_134),
.C(n_133),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_147),
.C(n_149),
.Y(n_156)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_156),
.A2(n_146),
.B(n_150),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_22),
.B(n_12),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_24),
.A3(n_13),
.B1(n_16),
.B2(n_20),
.C(n_47),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_162),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_146),
.CI(n_25),
.CON(n_164),
.SN(n_164)
);


endmodule