module fake_jpeg_31661_n_529 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_529);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_529;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_58),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_73),
.Y(n_106)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_31),
.B(n_16),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_15),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_101),
.Y(n_108)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_96),
.Y(n_148)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_100),
.Y(n_134)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_103),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_33),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_104),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_30),
.B1(n_46),
.B2(n_25),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_112),
.A2(n_27),
.B1(n_38),
.B2(n_45),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_132),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_31),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_31),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_156),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_38),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_22),
.B(n_29),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_153),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_61),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_62),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_34),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_50),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_75),
.A2(n_52),
.B1(n_48),
.B2(n_47),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_68),
.B1(n_65),
.B2(n_60),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_27),
.Y(n_165)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_175),
.B1(n_185),
.B2(n_186),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_176),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_108),
.A2(n_85),
.B1(n_95),
.B2(n_92),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_187),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_104),
.B1(n_88),
.B2(n_86),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_180),
.A2(n_218),
.B1(n_119),
.B2(n_158),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_20),
.B1(n_84),
.B2(n_77),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_181),
.A2(n_200),
.B1(n_202),
.B2(n_207),
.Y(n_230)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_58),
.B1(n_57),
.B2(n_59),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_108),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_190),
.Y(n_237)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_126),
.Y(n_190)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_192),
.B(n_193),
.Y(n_257)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_198),
.Y(n_227)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_196),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_106),
.B(n_45),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_201),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_20),
.B1(n_46),
.B2(n_30),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_203),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_106),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_208),
.Y(n_250)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_206),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_209),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_127),
.A2(n_56),
.B1(n_53),
.B2(n_30),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_157),
.B1(n_147),
.B2(n_141),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_138),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_148),
.Y(n_244)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_113),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_149),
.A2(n_20),
.B1(n_46),
.B2(n_47),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_217),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_220),
.Y(n_231)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_128),
.A2(n_48),
.B1(n_47),
.B2(n_41),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_219),
.A2(n_115),
.B1(n_20),
.B2(n_4),
.Y(n_255)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_162),
.B1(n_131),
.B2(n_136),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_222),
.A2(n_229),
.B1(n_232),
.B2(n_240),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_147),
.B1(n_165),
.B2(n_141),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_144),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_241),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_119),
.B1(n_123),
.B2(n_144),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_239),
.A2(n_247),
.B1(n_252),
.B2(n_4),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_191),
.A2(n_210),
.B1(n_186),
.B2(n_172),
.Y(n_240)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_188),
.A2(n_158),
.B1(n_145),
.B2(n_120),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_4),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_123),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_256),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_194),
.B(n_15),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_225),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_216),
.A2(n_145),
.B1(n_110),
.B2(n_22),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_172),
.A2(n_48),
.B1(n_41),
.B2(n_29),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_253),
.A2(n_258),
.B1(n_259),
.B2(n_200),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_1),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_180),
.A2(n_115),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_197),
.A2(n_205),
.B1(n_218),
.B2(n_178),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_206),
.C(n_193),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_266),
.C(n_280),
.Y(n_323)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_219),
.C(n_207),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_268),
.B(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_202),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_273),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_225),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_241),
.A2(n_171),
.B1(n_181),
.B2(n_168),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_274),
.B1(n_294),
.B2(n_261),
.Y(n_321)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_189),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_245),
.A2(n_214),
.B(n_167),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_277),
.A2(n_284),
.B(n_297),
.Y(n_326)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_203),
.C(n_183),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_235),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_281),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_231),
.B(n_2),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_288),
.Y(n_310)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_283),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_237),
.A2(n_196),
.B(n_5),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_259),
.B1(n_221),
.B2(n_229),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_290),
.Y(n_325)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_240),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_235),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_289),
.Y(n_305)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_250),
.B(n_5),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_255),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_221),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_295),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_244),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_296),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_231),
.A2(n_7),
.B(n_8),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_298),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_301),
.B(n_284),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_270),
.B(n_227),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_306),
.A2(n_319),
.B1(n_329),
.B2(n_307),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_239),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_277),
.C(n_266),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_241),
.Y(n_311)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_241),
.Y(n_314)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_279),
.B(n_269),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_316),
.A2(n_300),
.B(n_301),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g318 ( 
.A(n_278),
.B(n_262),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_262),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_285),
.A2(n_230),
.B1(n_236),
.B2(n_247),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_288),
.A2(n_224),
.B(n_228),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_320),
.A2(n_292),
.B(n_297),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_321),
.A2(n_296),
.B1(n_273),
.B2(n_264),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_251),
.Y(n_322)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_288),
.A2(n_253),
.B1(n_254),
.B2(n_248),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_295),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_309),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_261),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_323),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_333),
.A2(n_358),
.B1(n_356),
.B2(n_306),
.Y(n_378)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_335),
.B(n_342),
.Y(n_385)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_315),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_304),
.B(n_289),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_339),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_309),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_349),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_343),
.B(n_354),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_326),
.A2(n_320),
.B(n_300),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_344),
.A2(n_356),
.B(n_360),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_315),
.A2(n_276),
.B1(n_272),
.B2(n_248),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_345),
.A2(n_363),
.B1(n_319),
.B2(n_325),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_346),
.B(n_351),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_347),
.A2(n_350),
.B(n_353),
.Y(n_390)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_326),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_302),
.A2(n_305),
.B(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_302),
.B(n_281),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_305),
.A2(n_329),
.B(n_310),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_282),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_355),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_314),
.A2(n_274),
.B(n_263),
.Y(n_356)
);

NAND2x1_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_282),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_SL g371 ( 
.A(n_357),
.B(n_303),
.C(n_324),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_321),
.A2(n_263),
.B1(n_275),
.B2(n_265),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_308),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_359),
.B(n_332),
.Y(n_383)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_268),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_313),
.C(n_312),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_331),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_353),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_368),
.B(n_388),
.C(n_391),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_312),
.Y(n_369)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_364),
.B(n_322),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_370),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_371),
.B(n_360),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_378),
.A2(n_392),
.B1(n_363),
.B2(n_343),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_311),
.Y(n_379)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_324),
.Y(n_381)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_381),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_382),
.A2(n_357),
.B1(n_283),
.B2(n_295),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_383),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_355),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_386),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_350),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_317),
.C(n_260),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_317),
.C(n_260),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_358),
.A2(n_327),
.B1(n_330),
.B2(n_328),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_254),
.C(n_332),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_340),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_327),
.Y(n_394)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_396),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_360),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_399),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_390),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_377),
.B(n_364),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_401),
.B(n_403),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_340),
.Y(n_402)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_404),
.A2(n_384),
.B1(n_380),
.B2(n_396),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_386),
.A2(n_349),
.B(n_344),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_406),
.A2(n_410),
.B(n_392),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_411),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_380),
.A2(n_333),
.B(n_347),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_365),
.Y(n_414)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_414),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_375),
.B(n_348),
.Y(n_416)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_416),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_385),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_400),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_373),
.Y(n_420)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_420),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_357),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_423),
.Y(n_428)
);

INVx13_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_424),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_391),
.C(n_385),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_429),
.C(n_442),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_388),
.C(n_393),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_379),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_399),
.B1(n_406),
.B2(n_405),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_422),
.A2(n_390),
.B1(n_378),
.B2(n_374),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_437),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_389),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_440),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_368),
.C(n_408),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_389),
.C(n_394),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_428),
.Y(n_454)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_447),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_397),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_452),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_409),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_428),
.A2(n_417),
.B1(n_415),
.B2(n_403),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_453),
.A2(n_456),
.B1(n_365),
.B2(n_387),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_462),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_426),
.A2(n_417),
.B1(n_415),
.B2(n_412),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_457),
.A2(n_433),
.B1(n_434),
.B2(n_430),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_422),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_463),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_398),
.Y(n_461)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_405),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_399),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_442),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_412),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_429),
.C(n_418),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_421),
.B1(n_414),
.B2(n_418),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_466),
.A2(n_440),
.B1(n_425),
.B2(n_446),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_475),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_472),
.A2(n_473),
.B1(n_480),
.B2(n_283),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_451),
.A2(n_434),
.B1(n_439),
.B2(n_395),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_453),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_474),
.B(n_476),
.Y(n_484)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_459),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_SL g477 ( 
.A(n_458),
.B(n_427),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_477),
.A2(n_483),
.B(n_450),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_224),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_463),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_455),
.A2(n_376),
.B1(n_387),
.B2(n_366),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_456),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_482),
.Y(n_486)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_424),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_458),
.C(n_450),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_491),
.C(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_487),
.B(n_495),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_471),
.Y(n_489)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_489),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_493),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_448),
.C(n_460),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_468),
.B(n_448),
.C(n_376),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_366),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_473),
.Y(n_494)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_494),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_290),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_496),
.A2(n_498),
.B(n_490),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_480),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_287),
.B(n_242),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_505),
.Y(n_511)
);

OAI321xp33_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_474),
.A3(n_468),
.B1(n_223),
.B2(n_242),
.C(n_243),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_9),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_486),
.A2(n_249),
.B1(n_246),
.B2(n_243),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_504),
.B(n_13),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_485),
.A2(n_249),
.B1(n_238),
.B2(n_243),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_491),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_488),
.A2(n_238),
.B1(n_243),
.B2(n_11),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_509),
.B(n_492),
.Y(n_510)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_510),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_488),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_512),
.A2(n_513),
.B(n_514),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_10),
.C(n_11),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_515),
.A2(n_506),
.B(n_503),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g517 ( 
.A1(n_516),
.A2(n_501),
.B(n_499),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_517),
.A2(n_519),
.B(n_510),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_500),
.C(n_12),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_518),
.B(n_511),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_504),
.B(n_509),
.Y(n_523)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_523),
.Y(n_525)
);

MAJx2_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_524),
.C(n_12),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_11),
.B(n_12),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_12),
.Y(n_528)
);

FAx1_ASAP7_75t_SL g529 ( 
.A(n_528),
.B(n_13),
.CI(n_524),
.CON(n_529),
.SN(n_529)
);


endmodule