module fake_jpeg_25248_n_291 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_284;
wire n_288;
wire n_272;
wire n_234;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_8),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_49),
.B(n_19),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_28),
.B1(n_22),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_28),
.B1(n_33),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_23),
.B1(n_33),
.B2(n_30),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_36),
.B1(n_29),
.B2(n_34),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_36),
.B1(n_29),
.B2(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_18),
.B1(n_31),
.B2(n_27),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_18),
.B1(n_27),
.B2(n_30),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_41),
.B1(n_20),
.B2(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_46),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_77),
.B(n_81),
.Y(n_135)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_88),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_17),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx5_ASAP7_75t_SL g94 ( 
.A(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_99),
.Y(n_115)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_17),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_37),
.B(n_30),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_79),
.B(n_101),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_105),
.Y(n_122)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_27),
.B1(n_43),
.B2(n_40),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_56),
.B(n_24),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_60),
.B1(n_46),
.B2(n_65),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_109),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_55),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_60),
.B1(n_74),
.B2(n_41),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_128),
.B1(n_141),
.B2(n_82),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_39),
.C(n_42),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_134),
.C(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_112),
.B1(n_94),
.B2(n_98),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_13),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_19),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_42),
.B1(n_39),
.B2(n_21),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_42),
.C(n_39),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_42),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_32),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_32),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_21),
.B1(n_32),
.B2(n_20),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_142),
.B(n_153),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_97),
.B1(n_84),
.B2(n_91),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_149),
.B(n_159),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_102),
.B1(n_98),
.B2(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_95),
.B1(n_88),
.B2(n_110),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_162),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_24),
.Y(n_158)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_114),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_78),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_21),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_120),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_92),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_167),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_109),
.B1(n_104),
.B2(n_76),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_128),
.B1(n_119),
.B2(n_113),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_76),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_65),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_113),
.B(n_126),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_32),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_162),
.C(n_143),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_115),
.C(n_122),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.C(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_183),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_117),
.C(n_119),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_156),
.C(n_19),
.Y(n_211)
);

BUFx12f_ASAP7_75t_SL g219 ( 
.A(n_186),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_117),
.B1(n_127),
.B2(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_121),
.B1(n_104),
.B2(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_20),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_152),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_138),
.B1(n_116),
.B2(n_46),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_145),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_149),
.A2(n_20),
.A3(n_138),
.B1(n_116),
.B2(n_19),
.C1(n_5),
.C2(n_6),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_9),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_5),
.C2(n_7),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_19),
.B(n_0),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_1),
.B(n_2),
.Y(n_218)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_205),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_164),
.B(n_151),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_217),
.B(n_221),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_150),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_148),
.B(n_146),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_218),
.B(n_197),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_177),
.C(n_173),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_194),
.B1(n_187),
.B2(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_10),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_10),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_216),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_0),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_196),
.Y(n_220)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_210),
.A2(n_174),
.B1(n_176),
.B2(n_191),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_202),
.B1(n_201),
.B2(n_221),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_235),
.B(n_219),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_1),
.C(n_3),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_205),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_173),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_236),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_180),
.B(n_178),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_175),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_209),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_174),
.B1(n_181),
.B2(n_185),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_199),
.B1(n_202),
.B2(n_200),
.Y(n_242)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_246),
.B(n_248),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_249),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_251),
.B(n_252),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_245),
.B1(n_253),
.B2(n_235),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_201),
.B1(n_211),
.B2(n_215),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_224),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_231),
.C(n_11),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_206),
.C(n_184),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_254),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_218),
.B(n_214),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_226),
.B1(n_227),
.B2(n_233),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_231),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_259),
.B(n_246),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_238),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_236),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_228),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_R g275 ( 
.A(n_266),
.B(n_258),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_249),
.C(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_268),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_279),
.B(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_262),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_257),
.B(n_263),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_267),
.C(n_271),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_256),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_265),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_5),
.C2(n_16),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_270),
.B1(n_248),
.B2(n_275),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_14),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_285),
.B(n_14),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_287),
.A2(n_288),
.B(n_286),
.C(n_16),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_14),
.B(n_16),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_234),
.Y(n_291)
);


endmodule