module fake_aes_2403_n_27 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_14), .Y(n_18) );
AO31x2_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_12), .A3(n_13), .B(n_2), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_19), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_15), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_20), .Y(n_22) );
AOI221x1_ASAP7_75t_SL g23 ( .A1(n_22), .A2(n_1), .B1(n_13), .B2(n_7), .C(n_8), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_23), .B(n_1), .Y(n_24) );
INVx2_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_26), .B(n_24), .Y(n_27) );
endmodule