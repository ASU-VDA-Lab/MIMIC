module fake_jpeg_17603_n_83 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_10),
.B(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_9),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_40),
.B1(n_39),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_59),
.B1(n_32),
.B2(n_23),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_5),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_53),
.B(n_54),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_58),
.B1(n_60),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_35),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_25),
.B(n_38),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_56),
.B(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_6),
.B1(n_9),
.B2(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_22),
.B1(n_42),
.B2(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_30),
.B1(n_32),
.B2(n_45),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_65),
.Y(n_74)
);

XOR2x2_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_61),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_75),
.C(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_69),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

AOI221xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_73),
.B1(n_75),
.B2(n_68),
.C(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_68),
.C(n_67),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_81),
.B(n_57),
.C(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.Y(n_83)
);


endmodule