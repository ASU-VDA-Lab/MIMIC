module fake_jpeg_4951_n_92 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_92);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_92;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx5_ASAP7_75t_SL g29 ( 
.A(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_36),
.B(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_9),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_9),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_18),
.B1(n_30),
.B2(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_28),
.B1(n_29),
.B2(n_26),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_26),
.B(n_27),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_34),
.B(n_22),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_11),
.B1(n_14),
.B2(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_46),
.B(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_48),
.C(n_51),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_41),
.B1(n_22),
.B2(n_11),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_15),
.B(n_13),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_41),
.A3(n_14),
.B1(n_15),
.B2(n_17),
.C1(n_13),
.C2(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_67),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_13),
.B(n_10),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_57),
.B(n_10),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_55),
.B(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_61),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_67),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_80),
.C(n_74),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_6),
.B(n_8),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_57),
.Y(n_80)
);

OA21x2_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_82),
.B(n_1),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_23),
.C(n_6),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_77),
.Y(n_85)
);

AOI21x1_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_1),
.B(n_4),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_4),
.B(n_5),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_88),
.B(n_89),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_86),
.C(n_5),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_23),
.Y(n_92)
);


endmodule