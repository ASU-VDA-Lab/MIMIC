module fake_ibex_775_n_913 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_913);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_913;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_510;
wire n_193;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_894;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVxp33_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_51),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_70),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_72),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_28),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_166),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_52),
.B(n_47),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_12),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_58),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_97),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_24),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_9),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_43),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_29),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_24),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_74),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_31),
.Y(n_212)
);

BUFx2_ASAP7_75t_SL g213 ( 
.A(n_119),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_13),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_49),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_53),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_99),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_75),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_76),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_2),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_121),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_89),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_78),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_80),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_92),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_45),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_158),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_159),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_102),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_30),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_96),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_0),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_152),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_19),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_16),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_17),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_113),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_88),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_7),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_81),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_98),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_59),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_40),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_83),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_106),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_108),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_38),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_164),
.B(n_73),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_105),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_136),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_125),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_5),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_94),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_162),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_118),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_46),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_63),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_134),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_5),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_122),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_29),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_20),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_95),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_153),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_18),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_141),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_41),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_38),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_133),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_150),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_32),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_167),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

AND2x4_ASAP7_75t_SL g291 ( 
.A(n_190),
.B(n_44),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_50),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_239),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_177),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_187),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_176),
.B(n_2),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_203),
.A2(n_84),
.B(n_173),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_187),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_203),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_215),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_215),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_4),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

INVxp33_ASAP7_75t_SL g310 ( 
.A(n_178),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_193),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_180),
.B(n_6),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_197),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_242),
.B(n_7),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g319 ( 
.A(n_194),
.B(n_54),
.Y(n_319)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_194),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_197),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_202),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_179),
.B(n_10),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_238),
.A2(n_87),
.B(n_172),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_202),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_181),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_206),
.B(n_245),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_245),
.B(n_13),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_274),
.B(n_14),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_190),
.Y(n_332)
);

OAI22x1_ASAP7_75t_R g333 ( 
.A1(n_274),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_182),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_207),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_207),
.B(n_269),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_276),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_284),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_183),
.B(n_56),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_276),
.B(n_21),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_275),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_277),
.Y(n_346)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_234),
.Y(n_348)
);

AND2x2_ASAP7_75t_SL g349 ( 
.A(n_192),
.B(n_57),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_186),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_234),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_184),
.B(n_23),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_319),
.B(n_255),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_188),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_332),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_191),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_311),
.B(n_195),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

BUFx8_ASAP7_75t_SL g361 ( 
.A(n_332),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

BUFx4f_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_327),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_198),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_352),
.Y(n_369)
);

OR2x6_ASAP7_75t_L g370 ( 
.A(n_315),
.B(n_213),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_352),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_338),
.A2(n_255),
.B1(n_278),
.B2(n_280),
.Y(n_373)
);

AND3x2_ASAP7_75t_L g374 ( 
.A(n_315),
.B(n_346),
.C(n_307),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_350),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_199),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_310),
.B(n_201),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_319),
.B(n_278),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_289),
.B(n_204),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_329),
.B(n_293),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_313),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_352),
.Y(n_386)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_298),
.B(n_205),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_349),
.A2(n_250),
.B1(n_185),
.B2(n_209),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_316),
.B(n_195),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_316),
.B(n_208),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_291),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_289),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_290),
.Y(n_393)
);

OR2x6_ASAP7_75t_L g394 ( 
.A(n_321),
.B(n_200),
.Y(n_394)
);

BUFx6f_ASAP7_75t_SL g395 ( 
.A(n_337),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

INVx8_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_L g399 ( 
.A(n_330),
.B(n_224),
.C(n_210),
.Y(n_399)
);

OR2x6_ASAP7_75t_L g400 ( 
.A(n_314),
.B(n_241),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_295),
.B(n_211),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_243),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_337),
.B(n_216),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_331),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_292),
.B(n_217),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_218),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_302),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_302),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_303),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_304),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_336),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_291),
.B(n_244),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_304),
.B(n_221),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_306),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_319),
.A2(n_246),
.B1(n_254),
.B2(n_283),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_296),
.B(n_223),
.Y(n_423)
);

BUFx12f_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

NOR2x1p5_ASAP7_75t_L g425 ( 
.A(n_296),
.B(n_257),
.Y(n_425)
);

OAI22x1_ASAP7_75t_L g426 ( 
.A1(n_333),
.A2(n_214),
.B1(n_265),
.B2(n_282),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_301),
.B(n_225),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_317),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_305),
.B(n_226),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_328),
.A2(n_249),
.B1(n_228),
.B2(n_281),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_301),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_334),
.B(n_229),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_339),
.B(n_344),
.Y(n_436)
);

AO22x2_ASAP7_75t_L g437 ( 
.A1(n_339),
.A2(n_270),
.B1(n_230),
.B2(n_231),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_324),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_365),
.A2(n_344),
.B1(n_345),
.B2(n_352),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

OR2x6_ASAP7_75t_L g442 ( 
.A(n_370),
.B(n_400),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_219),
.Y(n_443)
);

AND2x6_ASAP7_75t_SL g444 ( 
.A(n_394),
.B(n_361),
.Y(n_444)
);

NOR3xp33_ASAP7_75t_L g445 ( 
.A(n_373),
.B(n_236),
.C(n_233),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_397),
.B(n_342),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_385),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_367),
.B(n_220),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_370),
.B(n_189),
.Y(n_449)
);

NOR2x1p5_ASAP7_75t_L g450 ( 
.A(n_357),
.B(n_222),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_355),
.A2(n_347),
.B1(n_341),
.B2(n_300),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_240),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

NOR3xp33_ASAP7_75t_SL g454 ( 
.A(n_373),
.B(n_258),
.C(n_287),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_388),
.A2(n_267),
.B1(n_248),
.B2(n_288),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_375),
.B(n_248),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_355),
.A2(n_347),
.B1(n_341),
.B2(n_300),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_424),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_414),
.B(n_253),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_414),
.B(n_258),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_380),
.B(n_263),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_432),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_390),
.B(n_263),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_268),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_421),
.B(n_251),
.Y(n_469)
);

OAI22xp33_ASAP7_75t_L g470 ( 
.A1(n_394),
.A2(n_279),
.B1(n_287),
.B2(n_256),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_366),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_421),
.B(n_398),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_387),
.B(n_232),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_356),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_356),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_428),
.B(n_259),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_428),
.B(n_264),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_387),
.B(n_235),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_388),
.A2(n_196),
.B1(n_271),
.B2(n_237),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_425),
.B(n_300),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_400),
.B(n_325),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_374),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_387),
.B(n_227),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_394),
.B(n_23),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_364),
.B(n_325),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

INVx8_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_413),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_426),
.B(n_261),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_391),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_359),
.B(n_341),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_404),
.B(n_312),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_355),
.A2(n_351),
.B1(n_348),
.B2(n_312),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_404),
.B(n_312),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_377),
.B(n_379),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_381),
.B(n_348),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_407),
.B(n_348),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_355),
.A2(n_351),
.B1(n_318),
.B2(n_309),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_354),
.B(n_297),
.Y(n_503)
);

NOR2x2_ASAP7_75t_L g504 ( 
.A(n_418),
.B(n_25),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_358),
.B(n_368),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

AND2x6_ASAP7_75t_SL g507 ( 
.A(n_423),
.B(n_25),
.Y(n_507)
);

OR2x6_ASAP7_75t_SL g508 ( 
.A(n_391),
.B(n_26),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_406),
.B(n_299),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_364),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_434),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_438),
.A2(n_505),
.B(n_471),
.C(n_466),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_447),
.B(n_382),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_389),
.B(n_382),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_468),
.B(n_437),
.Y(n_515)
);

AOI221xp5_ASAP7_75t_L g516 ( 
.A1(n_445),
.A2(n_399),
.B1(n_429),
.B2(n_376),
.C(n_431),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_442),
.B(n_383),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_490),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_448),
.B(n_406),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_448),
.B(n_406),
.Y(n_523)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_438),
.A2(n_429),
.B(n_427),
.C(n_401),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_500),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_490),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_508),
.Y(n_527)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_483),
.A2(n_419),
.B(n_435),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_452),
.B(n_419),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_456),
.A2(n_395),
.B1(n_435),
.B2(n_422),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_446),
.A2(n_433),
.B(n_378),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_477),
.A2(n_396),
.B(n_417),
.C(n_416),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_489),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_459),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_449),
.B(n_27),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_SL g536 ( 
.A1(n_503),
.A2(n_402),
.B(n_412),
.C(n_411),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_449),
.B(n_28),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_472),
.A2(n_386),
.B(n_372),
.Y(n_539)
);

CKINVDCx8_ASAP7_75t_R g540 ( 
.A(n_444),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_482),
.A2(n_430),
.B1(n_386),
.B2(n_372),
.Y(n_541)
);

AOI22x1_ASAP7_75t_L g542 ( 
.A1(n_483),
.A2(n_386),
.B1(n_372),
.B2(n_369),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

O2A1O1Ixp33_ASAP7_75t_SL g544 ( 
.A1(n_503),
.A2(n_109),
.B(n_174),
.C(n_171),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_472),
.A2(n_369),
.B(n_318),
.Y(n_545)
);

A2O1A1Ixp33_ASAP7_75t_L g546 ( 
.A1(n_477),
.A2(n_318),
.B(n_309),
.C(n_299),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_443),
.Y(n_547)
);

A2O1A1Ixp33_ASAP7_75t_L g548 ( 
.A1(n_478),
.A2(n_318),
.B(n_309),
.C(n_299),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_486),
.B(n_299),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g550 ( 
.A(n_507),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_496),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_451),
.A2(n_103),
.B(n_165),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_494),
.B(n_510),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_498),
.Y(n_554)
);

A2O1A1Ixp33_ASAP7_75t_L g555 ( 
.A1(n_481),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_484),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_463),
.B(n_467),
.Y(n_557)
);

A2O1A1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_493),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_485),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_458),
.A2(n_114),
.B(n_163),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_40),
.Y(n_561)
);

AOI33xp33_ASAP7_75t_L g562 ( 
.A1(n_470),
.A2(n_41),
.A3(n_42),
.B1(n_60),
.B2(n_61),
.B3(n_62),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_475),
.Y(n_563)
);

AOI22x1_ASAP7_75t_L g564 ( 
.A1(n_488),
.A2(n_440),
.B1(n_441),
.B2(n_453),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_455),
.A2(n_470),
.B1(n_454),
.B2(n_465),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_458),
.A2(n_117),
.B(n_64),
.Y(n_566)
);

AOI33xp33_ASAP7_75t_L g567 ( 
.A1(n_439),
.A2(n_42),
.A3(n_65),
.B1(n_66),
.B2(n_67),
.B3(n_68),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_506),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_473),
.B(n_69),
.Y(n_569)
);

BUFx8_ASAP7_75t_L g570 ( 
.A(n_504),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_461),
.B(n_77),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_462),
.B(n_79),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_492),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_479),
.B(n_82),
.Y(n_574)
);

AO32x1_ASAP7_75t_L g575 ( 
.A1(n_511),
.A2(n_85),
.A3(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_480),
.B(n_168),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_469),
.B(n_460),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_497),
.B(n_104),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_497),
.B(n_112),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_492),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_534),
.Y(n_581)
);

OAI221xp5_ASAP7_75t_L g582 ( 
.A1(n_557),
.A2(n_492),
.B1(n_439),
.B2(n_469),
.C(n_501),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_512),
.A2(n_495),
.B(n_457),
.C(n_464),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_529),
.B(n_450),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_564),
.A2(n_545),
.B(n_566),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_518),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_568),
.Y(n_587)
);

A2O1A1Ixp33_ASAP7_75t_L g588 ( 
.A1(n_524),
.A2(n_495),
.B(n_509),
.C(n_502),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_553),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_543),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_522),
.A2(n_523),
.B(n_514),
.Y(n_592)
);

INVx6_ASAP7_75t_SL g593 ( 
.A(n_561),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_531),
.A2(n_126),
.B(n_127),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_516),
.B(n_129),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_518),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_513),
.A2(n_131),
.B(n_132),
.Y(n_597)
);

AO31x2_ASAP7_75t_L g598 ( 
.A1(n_528),
.A2(n_135),
.A3(n_138),
.B(n_139),
.Y(n_598)
);

AOI31xp67_ASAP7_75t_L g599 ( 
.A1(n_569),
.A2(n_574),
.A3(n_576),
.B(n_578),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_540),
.B(n_140),
.Y(n_601)
);

AO31x2_ASAP7_75t_L g602 ( 
.A1(n_546),
.A2(n_143),
.A3(n_145),
.B(n_146),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_551),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_553),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_577),
.A2(n_154),
.B(n_155),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_565),
.B(n_554),
.Y(n_606)
);

AO31x2_ASAP7_75t_L g607 ( 
.A1(n_548),
.A2(n_552),
.A3(n_560),
.B(n_515),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_525),
.A2(n_571),
.B(n_572),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_517),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_570),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_519),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_535),
.A2(n_538),
.B1(n_518),
.B2(n_561),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_549),
.A2(n_536),
.B(n_530),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_SL g615 ( 
.A1(n_579),
.A2(n_558),
.B(n_555),
.C(n_541),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_561),
.B(n_520),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_556),
.Y(n_617)
);

AO31x2_ASAP7_75t_L g618 ( 
.A1(n_567),
.A2(n_575),
.A3(n_562),
.B(n_544),
.Y(n_618)
);

AO21x2_ASAP7_75t_L g619 ( 
.A1(n_575),
.A2(n_573),
.B(n_559),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_521),
.B(n_526),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_526),
.Y(n_621)
);

INVx3_ASAP7_75t_SL g622 ( 
.A(n_526),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_550),
.B(n_537),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_537),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_568),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_534),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_542),
.A2(n_539),
.B(n_564),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g630 ( 
.A(n_540),
.B(n_332),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_529),
.B(n_505),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_521),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_512),
.A2(n_557),
.B(n_438),
.C(n_524),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_529),
.B(n_505),
.Y(n_634)
);

BUFx10_ASAP7_75t_L g635 ( 
.A(n_553),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_521),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_529),
.B(n_505),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_527),
.A2(n_447),
.B(n_374),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_SL g639 ( 
.A1(n_512),
.A2(n_524),
.B(n_532),
.C(n_569),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_529),
.B(n_447),
.Y(n_640)
);

AO31x2_ASAP7_75t_L g641 ( 
.A1(n_528),
.A2(n_512),
.A3(n_545),
.B(n_546),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_529),
.B(n_505),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_518),
.B(n_447),
.Y(n_643)
);

CKINVDCx8_ASAP7_75t_R g644 ( 
.A(n_573),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_542),
.A2(n_539),
.B(n_564),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_547),
.B(n_447),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_521),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_529),
.B(n_505),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_529),
.B(n_447),
.Y(n_649)
);

AO31x2_ASAP7_75t_L g650 ( 
.A1(n_528),
.A2(n_512),
.A3(n_545),
.B(n_546),
.Y(n_650)
);

AO31x2_ASAP7_75t_L g651 ( 
.A1(n_528),
.A2(n_512),
.A3(n_545),
.B(n_546),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_529),
.B(n_447),
.Y(n_652)
);

AO31x2_ASAP7_75t_L g653 ( 
.A1(n_528),
.A2(n_512),
.A3(n_545),
.B(n_546),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_542),
.A2(n_539),
.B(n_564),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_534),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_529),
.B(n_447),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_542),
.A2(n_539),
.B(n_564),
.Y(n_657)
);

AO31x2_ASAP7_75t_L g658 ( 
.A1(n_592),
.A2(n_633),
.A3(n_614),
.B(n_595),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_630),
.A2(n_593),
.B1(n_631),
.B2(n_634),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_637),
.B(n_642),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_648),
.B(n_606),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_640),
.B(n_649),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_603),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_626),
.B(n_617),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_584),
.A2(n_593),
.B1(n_652),
.B2(n_656),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_612),
.A2(n_626),
.B1(n_586),
.B2(n_643),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_587),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_629),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g669 ( 
.A1(n_585),
.A2(n_657),
.B(n_654),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_609),
.B(n_643),
.Y(n_670)
);

NOR2x1_ASAP7_75t_SL g671 ( 
.A(n_647),
.B(n_632),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_588),
.B(n_615),
.C(n_583),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_616),
.B(n_590),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_609),
.B(n_596),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_647),
.B(n_613),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_635),
.B(n_622),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_611),
.B(n_580),
.Y(n_677)
);

AOI221xp5_ASAP7_75t_L g678 ( 
.A1(n_638),
.A2(n_655),
.B1(n_582),
.B2(n_604),
.C(n_627),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_589),
.B(n_591),
.Y(n_679)
);

AO21x2_ASAP7_75t_L g680 ( 
.A1(n_594),
.A2(n_597),
.B(n_605),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_600),
.Y(n_681)
);

BUFx8_ASAP7_75t_L g682 ( 
.A(n_625),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_619),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_641),
.B(n_653),
.Y(n_684)
);

INVx4_ASAP7_75t_SL g685 ( 
.A(n_602),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_641),
.B(n_653),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_624),
.Y(n_687)
);

AO21x2_ASAP7_75t_L g688 ( 
.A1(n_618),
.A2(n_598),
.B(n_599),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_620),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_647),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_613),
.Y(n_691)
);

AO21x2_ASAP7_75t_L g692 ( 
.A1(n_618),
.A2(n_598),
.B(n_651),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_635),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_636),
.A2(n_621),
.B(n_650),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_581),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_636),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_650),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_623),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_601),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_610),
.B(n_607),
.Y(n_700)
);

A2O1A1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_644),
.A2(n_633),
.B(n_512),
.C(n_365),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_622),
.Y(n_702)
);

OA21x2_ASAP7_75t_L g703 ( 
.A1(n_585),
.A2(n_645),
.B(n_628),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_603),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_646),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_603),
.Y(n_706)
);

BUFx8_ASAP7_75t_L g707 ( 
.A(n_625),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_610),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_603),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_631),
.B(n_634),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_633),
.A2(n_512),
.B(n_606),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_603),
.Y(n_712)
);

AO31x2_ASAP7_75t_L g713 ( 
.A1(n_592),
.A2(n_528),
.A3(n_633),
.B(n_614),
.Y(n_713)
);

INVx11_ASAP7_75t_L g714 ( 
.A(n_622),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_608),
.A2(n_639),
.B(n_633),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_603),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_593),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_610),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_633),
.B(n_631),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_633),
.B(n_631),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_593),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_603),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_631),
.B(n_634),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_647),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_603),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_603),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_584),
.A2(n_365),
.B1(n_447),
.B2(n_445),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_633),
.B(n_631),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_633),
.B(n_631),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_633),
.B(n_631),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_694),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_704),
.B(n_706),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_723),
.B(n_660),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_695),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_694),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_664),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_663),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_709),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_712),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_714),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_722),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_662),
.Y(n_742)
);

AOI222xp33_ASAP7_75t_L g743 ( 
.A1(n_660),
.A2(n_710),
.B1(n_661),
.B2(n_659),
.C1(n_666),
.C2(n_727),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_679),
.B(n_716),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_666),
.B(n_700),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_725),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_726),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_691),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_691),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_700),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_711),
.B(n_715),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_661),
.B(n_674),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_711),
.B(n_667),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_675),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_690),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_681),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_668),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_684),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_719),
.B(n_720),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_728),
.B(n_729),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_675),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_686),
.A2(n_672),
.B(n_683),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_702),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_691),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_728),
.B(n_730),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_729),
.B(n_730),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_670),
.B(n_673),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_678),
.A2(n_705),
.B1(n_665),
.B2(n_699),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_697),
.Y(n_769)
);

INVx11_ASAP7_75t_L g770 ( 
.A(n_682),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_689),
.Y(n_771)
);

AO21x2_ASAP7_75t_L g772 ( 
.A1(n_688),
.A2(n_669),
.B(n_692),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_677),
.B(n_692),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_701),
.B(n_687),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_713),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_724),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_703),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_658),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_671),
.B(n_696),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_676),
.Y(n_780)
);

INVxp67_ASAP7_75t_R g781 ( 
.A(n_718),
.Y(n_781)
);

AOI21x1_ASAP7_75t_L g782 ( 
.A1(n_685),
.A2(n_693),
.B(n_680),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_685),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_708),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_777),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_750),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_758),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_736),
.B(n_698),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_753),
.B(n_717),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_753),
.B(n_721),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_744),
.B(n_682),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_744),
.B(n_707),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_759),
.B(n_765),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_773),
.B(n_707),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_765),
.B(n_751),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_751),
.B(n_745),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_783),
.B(n_745),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_773),
.B(n_750),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_751),
.B(n_745),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_733),
.B(n_752),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_769),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

NOR2xp67_ASAP7_75t_L g803 ( 
.A(n_783),
.B(n_748),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_745),
.B(n_752),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_767),
.B(n_742),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_751),
.B(n_737),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_738),
.B(n_739),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_754),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_760),
.B(n_766),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_746),
.B(n_747),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_746),
.B(n_747),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_754),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_732),
.B(n_741),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_795),
.B(n_731),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_795),
.B(n_735),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_798),
.B(n_735),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_793),
.B(n_762),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_793),
.B(n_806),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_802),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_785),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_802),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_797),
.B(n_782),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_796),
.B(n_772),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_801),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_794),
.B(n_768),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_797),
.B(n_799),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_799),
.B(n_807),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_787),
.B(n_774),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_807),
.B(n_775),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_810),
.B(n_811),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_798),
.B(n_778),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_804),
.B(n_778),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_822),
.B(n_797),
.Y(n_833)
);

AOI21xp33_ASAP7_75t_L g834 ( 
.A1(n_825),
.A2(n_794),
.B(n_743),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_819),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_819),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_825),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_828),
.B(n_800),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_830),
.B(n_813),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_821),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_818),
.B(n_789),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_818),
.B(n_830),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_829),
.B(n_813),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_824),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_828),
.B(n_800),
.Y(n_845)
);

NOR2x1_ASAP7_75t_L g846 ( 
.A(n_822),
.B(n_791),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_816),
.B(n_805),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_L g848 ( 
.A(n_822),
.B(n_791),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_822),
.B(n_786),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_821),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_826),
.B(n_797),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_820),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_826),
.B(n_823),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_844),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_852),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_844),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_842),
.B(n_817),
.Y(n_857)
);

OAI22xp33_ASAP7_75t_L g858 ( 
.A1(n_846),
.A2(n_804),
.B1(n_812),
.B2(n_786),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_835),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_847),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_848),
.Y(n_861)
);

OAI22xp33_ASAP7_75t_L g862 ( 
.A1(n_849),
.A2(n_812),
.B1(n_808),
.B2(n_805),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_836),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_840),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_838),
.B(n_817),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_859),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_859),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_855),
.Y(n_868)
);

OAI221xp5_ASAP7_75t_L g869 ( 
.A1(n_861),
.A2(n_834),
.B1(n_837),
.B2(n_849),
.C(n_845),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_858),
.A2(n_849),
.B1(n_853),
.B2(n_851),
.Y(n_870)
);

OAI21xp33_ASAP7_75t_L g871 ( 
.A1(n_865),
.A2(n_838),
.B(n_845),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_854),
.B(n_833),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_854),
.B(n_833),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_860),
.A2(n_833),
.B1(n_792),
.B2(n_853),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_864),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_862),
.A2(n_824),
.B(n_808),
.Y(n_876)
);

OAI322xp33_ASAP7_75t_L g877 ( 
.A1(n_856),
.A2(n_839),
.A3(n_843),
.B1(n_816),
.B2(n_832),
.C1(n_831),
.C2(n_841),
.Y(n_877)
);

AOI221xp5_ASAP7_75t_L g878 ( 
.A1(n_877),
.A2(n_856),
.B1(n_863),
.B2(n_864),
.C(n_857),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_869),
.A2(n_853),
.B1(n_792),
.B2(n_851),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_874),
.A2(n_857),
.B1(n_851),
.B2(n_826),
.Y(n_880)
);

AOI221x1_ASAP7_75t_SL g881 ( 
.A1(n_871),
.A2(n_788),
.B1(n_781),
.B2(n_809),
.C(n_756),
.Y(n_881)
);

AOI222xp33_ASAP7_75t_L g882 ( 
.A1(n_870),
.A2(n_734),
.B1(n_789),
.B2(n_790),
.C1(n_823),
.C2(n_788),
.Y(n_882)
);

AOI221xp5_ASAP7_75t_L g883 ( 
.A1(n_866),
.A2(n_763),
.B1(n_850),
.B2(n_814),
.C(n_815),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_876),
.A2(n_781),
.B(n_755),
.Y(n_884)
);

OAI211xp5_ASAP7_75t_L g885 ( 
.A1(n_879),
.A2(n_884),
.B(n_878),
.C(n_882),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_880),
.A2(n_776),
.B(n_881),
.C(n_780),
.Y(n_886)
);

AOI322xp5_ASAP7_75t_L g887 ( 
.A1(n_883),
.A2(n_873),
.A3(n_872),
.B1(n_827),
.B2(n_867),
.C1(n_875),
.C2(n_790),
.Y(n_887)
);

OAI211xp5_ASAP7_75t_L g888 ( 
.A1(n_885),
.A2(n_740),
.B(n_784),
.C(n_770),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_886),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_889),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_888),
.A2(n_740),
.B(n_873),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_890),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_891),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_893),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_892),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_894),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_895),
.B(n_770),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_894),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_896),
.A2(n_889),
.B1(n_887),
.B2(n_780),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_898),
.B(n_872),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_897),
.A2(n_761),
.B1(n_774),
.B2(n_771),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_896),
.B(n_868),
.Y(n_902)
);

OAI21x1_ASAP7_75t_L g903 ( 
.A1(n_896),
.A2(n_756),
.B(n_757),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_900),
.B(n_757),
.Y(n_904)
);

OA21x2_ASAP7_75t_L g905 ( 
.A1(n_903),
.A2(n_771),
.B(n_779),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_901),
.Y(n_906)
);

AOI21xp33_ASAP7_75t_L g907 ( 
.A1(n_899),
.A2(n_764),
.B(n_749),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_SL g908 ( 
.A(n_902),
.B(n_764),
.Y(n_908)
);

AO21x2_ASAP7_75t_L g909 ( 
.A1(n_906),
.A2(n_803),
.B(n_779),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_904),
.Y(n_910)
);

NAND2x1_ASAP7_75t_L g911 ( 
.A(n_905),
.B(n_748),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_910),
.B(n_907),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_912),
.A2(n_908),
.B1(n_909),
.B2(n_911),
.Y(n_913)
);


endmodule