module fake_netlist_1_4121_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
OAI22xp5_ASAP7_75t_SL g12 ( .A1(n_8), .A2(n_3), .B1(n_4), .B2(n_10), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_11), .B(n_1), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_13), .B(n_1), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_2), .B1(n_5), .B2(n_6), .Y(n_18) );
AO31x2_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_14), .A3(n_15), .B(n_11), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
OAI21xp5_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_21), .B(n_17), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_19), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_12), .B1(n_18), .B2(n_14), .Y(n_29) );
INVxp67_ASAP7_75t_SL g30 ( .A(n_27), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_19), .Y(n_31) );
NOR4xp75_ASAP7_75t_L g32 ( .A(n_29), .B(n_2), .C(n_5), .D(n_6), .Y(n_32) );
INVx1_ASAP7_75t_SL g33 ( .A(n_32), .Y(n_33) );
XNOR2xp5_ASAP7_75t_L g34 ( .A(n_30), .B(n_19), .Y(n_34) );
OAI22x1_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_31), .B1(n_19), .B2(n_9), .Y(n_35) );
AOI22xp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_33), .B1(n_34), .B2(n_7), .Y(n_36) );
endmodule