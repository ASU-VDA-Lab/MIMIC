module fake_jpeg_25032_n_257 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_6),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_39),
.Y(n_40)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_21),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_50),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_21),
.B1(n_25),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_28),
.B1(n_38),
.B2(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_59),
.B1(n_64),
.B2(n_66),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_38),
.B1(n_28),
.B2(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_17),
.B1(n_28),
.B2(n_27),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_68),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_28),
.B1(n_17),
.B2(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_17),
.B1(n_27),
.B2(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_17),
.B1(n_34),
.B2(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_75),
.Y(n_81)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_22),
.B1(n_23),
.B2(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_76),
.B1(n_20),
.B2(n_26),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_34),
.B1(n_15),
.B2(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_25),
.B1(n_29),
.B2(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_55),
.B1(n_26),
.B2(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_20),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_14),
.B1(n_19),
.B2(n_11),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_0),
.B(n_1),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_14),
.B(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_16),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_14),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_104),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_59),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_22),
.C(n_23),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_110),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_62),
.B1(n_67),
.B2(n_69),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_116),
.B1(n_87),
.B2(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_57),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_123),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_121),
.B(n_85),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_70),
.B1(n_71),
.B2(n_65),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_119),
.B1(n_99),
.B2(n_22),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_103),
.B1(n_104),
.B2(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_82),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_70),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_16),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_126),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_132),
.B(n_137),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_121),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_97),
.C(n_90),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_151),
.C(n_122),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_85),
.B(n_90),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_142),
.B(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_121),
.B1(n_118),
.B2(n_125),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_90),
.C(n_100),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_150),
.B1(n_115),
.B2(n_120),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_96),
.B(n_14),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_146),
.Y(n_169)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_149),
.B1(n_127),
.B2(n_112),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_99),
.B1(n_35),
.B2(n_37),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_23),
.B1(n_22),
.B2(n_14),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_16),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_6),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_46),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_136),
.B1(n_129),
.B2(n_151),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_172),
.B(n_167),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_35),
.Y(n_194)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_112),
.B1(n_110),
.B2(n_128),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_37),
.B1(n_35),
.B2(n_7),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_134),
.B1(n_142),
.B2(n_132),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_46),
.C(n_54),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_154),
.C(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_148),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_166),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_182),
.B1(n_191),
.B2(n_194),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_144),
.C(n_153),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_46),
.C(n_54),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_170),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_172),
.B1(n_171),
.B2(n_165),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_46),
.C(n_37),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_195),
.C(n_162),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_161),
.B1(n_157),
.B2(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_159),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_196),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_207),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_205),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_164),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_209),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_210),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_160),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_173),
.C(n_172),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_184),
.C(n_195),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_218),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_211),
.A2(n_188),
.B1(n_185),
.B2(n_163),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_168),
.B1(n_158),
.B2(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_194),
.B(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_171),
.B(n_159),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_221),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_171),
.B(n_179),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_216),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_3),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_210),
.B1(n_193),
.B2(n_203),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_4),
.B1(n_9),
.B2(n_8),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_203),
.C(n_204),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_228),
.C(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_5),
.C(n_10),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_5),
.C(n_10),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_221),
.B(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_233),
.A2(n_220),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_212),
.B1(n_4),
.B2(n_3),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_240),
.C(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_225),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_245),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_230),
.A3(n_227),
.B1(n_8),
.B2(n_12),
.C1(n_2),
.C2(n_1),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_0),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_230),
.C(n_1),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_242),
.C(n_246),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_250),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_2),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_249),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_253),
.B(n_248),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_251),
.Y(n_256)
);

XNOR2x2_ASAP7_75t_SL g257 ( 
.A(n_256),
.B(n_2),
.Y(n_257)
);


endmodule