module real_jpeg_1481_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_167;
wire n_128;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_2),
.A2(n_39),
.B1(n_59),
.B2(n_61),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_2),
.B(n_57),
.C(n_59),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_39),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_39),
.B1(n_63),
.B2(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_2),
.B(n_55),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_40),
.C(n_74),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_2),
.B(n_24),
.C(n_46),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_72),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_2),
.B(n_31),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_2),
.B(n_50),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_65),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_65),
.Y(n_217)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_35),
.B1(n_63),
.B2(n_66),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_10),
.A2(n_35),
.B1(n_59),
.B2(n_61),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_135),
.B1(n_253),
.B2(n_254),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_134),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_109),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_17),
.B(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_82),
.C(n_100),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_18),
.A2(n_19),
.B1(n_100),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_20),
.B(n_71),
.C(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_21),
.B(n_36),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_32),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_22),
.A2(n_30),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_24),
.B(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_29),
.B(n_34),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_29),
.A2(n_30),
.B(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_29),
.B(n_108),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_29),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_30),
.B(n_217),
.Y(n_231)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_31),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_32),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_33),
.B(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_49),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_37),
.B(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_38),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_38),
.B(n_50),
.Y(n_188)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_42),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_40),
.B(n_211),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_43),
.B(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_43),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_43),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

OAI21x1_ASAP7_75t_SL g131 ( 
.A1(n_49),
.A2(n_103),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_49),
.B(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_50),
.B(n_190),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_71),
.B1(n_80),
.B2(n_81),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_67),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_54),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_62),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_55),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_57),
.B1(n_63),
.B2(n_66),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_61),
.B1(n_74),
.B2(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_59),
.B(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_97),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_79),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_72),
.B(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_76),
.B(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_77),
.B(n_124),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_94),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_91),
.B(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_99),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_105),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

AOI21x1_ASAP7_75t_SL g151 ( 
.A1(n_102),
.A2(n_132),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_104),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_106),
.B(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_127),
.B2(n_128),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_129),
.A2(n_130),
.B1(n_183),
.B2(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_157),
.B(n_250),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_137),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_138),
.B(n_141),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_145),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_153),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_175),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_159),
.B(n_161),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_163),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_231),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_194),
.B(n_249),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_191),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_177),
.B(n_191),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_186),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_179),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21x1_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_205),
.B(n_248),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_204),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_203),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_246),
.Y(n_245)
);

OAI21x1_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_243),
.B(n_247),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_225),
.B(n_242),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B1(n_219),
.B2(n_224),
.Y(n_213)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.C(n_224),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_241),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_229),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_237),
.B(n_240),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);


endmodule