module real_jpeg_30795_n_20 (n_17, n_8, n_0, n_2, n_692, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_692;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_578;
wire n_332;
wire n_366;
wire n_149;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_611;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_689;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_690;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_0),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_0),
.Y(n_275)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_0),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_179),
.B1(n_180),
.B2(n_185),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_1),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_1),
.A2(n_179),
.B1(n_238),
.B2(n_243),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_1),
.A2(n_179),
.B1(n_391),
.B2(n_395),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_1),
.A2(n_179),
.B1(n_643),
.B2(n_645),
.Y(n_642)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_2),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_4),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_4),
.A2(n_130),
.B1(n_291),
.B2(n_295),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_4),
.A2(n_130),
.B1(n_402),
.B2(n_404),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_4),
.A2(n_130),
.B1(n_267),
.B2(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_5),
.A2(n_164),
.B1(n_169),
.B2(n_170),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_5),
.A2(n_169),
.B1(n_337),
.B2(n_341),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_5),
.A2(n_169),
.B1(n_448),
.B2(n_450),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_5),
.A2(n_169),
.B1(n_201),
.B2(n_639),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_6),
.A2(n_55),
.B(n_219),
.Y(n_288)
);

INVx2_ASAP7_75t_R g326 ( 
.A(n_6),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_6),
.A2(n_326),
.B1(n_517),
.B2(n_519),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_6),
.B(n_113),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_6),
.A2(n_189),
.B1(n_589),
.B2(n_593),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_67),
.B1(n_71),
.B2(n_74),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_7),
.A2(n_74),
.B1(n_352),
.B2(n_355),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_7),
.A2(n_74),
.B1(n_439),
.B2(n_443),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_7),
.A2(n_74),
.B1(n_629),
.B2(n_632),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_9),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_10),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_10),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_11),
.A2(n_64),
.B1(n_266),
.B2(n_271),
.Y(n_265)
);

AOI22x1_ASAP7_75t_L g416 ( 
.A1(n_11),
.A2(n_64),
.B1(n_417),
.B2(n_419),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_11),
.A2(n_64),
.B1(n_367),
.B2(n_624),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_12),
.A2(n_136),
.B1(n_142),
.B2(n_146),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_12),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_12),
.A2(n_146),
.B1(n_374),
.B2(n_376),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_12),
.A2(n_146),
.B1(n_480),
.B2(n_485),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_12),
.A2(n_146),
.B1(n_530),
.B2(n_532),
.Y(n_529)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_13),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_14),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_14),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_14),
.A2(n_261),
.B1(n_319),
.B2(n_323),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_14),
.A2(n_261),
.B1(n_366),
.B2(n_369),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_14),
.A2(n_61),
.B1(n_95),
.B2(n_261),
.Y(n_457)
);

AOI22x1_ASAP7_75t_SL g93 ( 
.A1(n_15),
.A2(n_94),
.B1(n_98),
.B2(n_101),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_15),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_15),
.A2(n_101),
.B1(n_279),
.B2(n_284),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_15),
.A2(n_101),
.B1(n_243),
.B2(n_511),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_15),
.A2(n_101),
.B1(n_581),
.B2(n_583),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_21),
.B(n_689),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_16),
.B(n_690),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_17),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_17),
.A2(n_107),
.B1(n_308),
.B2(n_314),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_17),
.A2(n_107),
.B1(n_258),
.B2(n_538),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_17),
.A2(n_107),
.B1(n_590),
.B2(n_592),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_18),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_18),
.Y(n_125)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_18),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_18),
.Y(n_513)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_19),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_19),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_19),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_81),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_76),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_24),
.B(n_681),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_24),
.B(n_681),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_25),
.B(n_77),
.Y(n_81)
);

NAND4xp25_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_53),
.C(n_65),
.D(n_75),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_49),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_27),
.A2(n_49),
.B1(n_638),
.B2(n_641),
.Y(n_637)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_28),
.A2(n_50),
.B1(n_457),
.B2(n_642),
.Y(n_654)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_29),
.A2(n_51),
.B1(n_104),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_29),
.A2(n_51),
.B1(n_93),
.B2(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_29),
.A2(n_51),
.B1(n_373),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_34),
.Y(n_204)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_34),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_36),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_37),
.Y(n_403)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_37),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_37),
.Y(n_646)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_42),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_43),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_43),
.Y(n_635)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_46),
.Y(n_152)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_46),
.Y(n_627)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_66),
.B(n_78),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_91),
.B(n_102),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_49),
.A2(n_54),
.B1(n_78),
.B2(n_638),
.Y(n_650)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22x1_ASAP7_75t_L g456 ( 
.A1(n_50),
.A2(n_79),
.B1(n_401),
.B2(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2x1_ASAP7_75t_R g325 ( 
.A(n_51),
.B(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_56),
.Y(n_220)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_58),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_59),
.Y(n_375)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_63),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_617),
.B(n_682),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_469),
.B(n_612),
.Y(n_84)
);

NAND4xp25_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_329),
.C(n_426),
.D(n_461),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_299),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_87),
.B(n_299),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_221),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_88),
.A2(n_463),
.B(n_464),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_159),
.Y(n_88)
);

XNOR2x1_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_111),
.Y(n_89)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_90),
.Y(n_332)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_111),
.B(n_159),
.C(n_332),
.Y(n_331)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_126),
.B1(n_135),
.B2(n_147),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_112),
.A2(n_135),
.B1(n_147),
.B2(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_112),
.A2(n_278),
.B(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_112),
.A2(n_126),
.B1(n_147),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_112),
.A2(n_147),
.B1(n_307),
.B2(n_516),
.Y(n_515)
);

OAI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_112),
.A2(n_147),
.B1(n_623),
.B2(n_628),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g655 ( 
.A1(n_112),
.A2(n_147),
.B1(n_623),
.B2(n_656),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22x1_ASAP7_75t_SL g388 ( 
.A1(n_113),
.A2(n_305),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_113),
.A2(n_305),
.B1(n_390),
.B2(n_447),
.Y(n_446)
);

OAI21xp33_ASAP7_75t_SL g648 ( 
.A1(n_113),
.A2(n_305),
.B(n_649),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AO21x2_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_148),
.B(n_153),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B1(n_121),
.B2(n_124),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_119),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_119),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_120),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_120),
.Y(n_343)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_120),
.Y(n_442)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_124),
.B(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_124),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_124),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_125),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_125),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_125),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_129),
.Y(n_451)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_134),
.Y(n_286)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_134),
.Y(n_631)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_141),
.Y(n_283)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_144),
.Y(n_449)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_145),
.Y(n_520)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_147),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_153),
.A2(n_490),
.B(n_495),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_155),
.Y(n_314)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_195),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_160),
.A2(n_161),
.B1(n_195),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_172),
.B1(n_178),
.B2(n_188),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_163),
.A2(n_189),
.B1(n_265),
.B2(n_273),
.Y(n_264)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_168),
.Y(n_531)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_171),
.Y(n_272)
);

BUFx2_ASAP7_75t_SL g324 ( 
.A(n_171),
.Y(n_324)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_173),
.B(n_326),
.Y(n_595)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_177),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_177),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_178),
.A2(n_188),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_184),
.Y(n_562)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g499 ( 
.A1(n_188),
.A2(n_318),
.B1(n_500),
.B2(n_504),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_188),
.A2(n_346),
.B1(n_578),
.B2(n_579),
.Y(n_577)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_189),
.A2(n_265),
.B(n_345),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_189),
.A2(n_351),
.B(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_189),
.A2(n_525),
.B1(n_528),
.B2(n_529),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_189),
.A2(n_525),
.B1(n_580),
.B2(n_589),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_192),
.Y(n_584)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_193),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_194),
.Y(n_504)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_194),
.Y(n_593)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_195),
.Y(n_328)
);

OAI22x1_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_205),
.B1(n_208),
.B2(n_218),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_217),
.Y(n_397)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_276),
.B1(n_297),
.B2(n_298),
.Y(n_221)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_264),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_223),
.B(n_264),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_237),
.B1(n_246),
.B2(n_257),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_224),
.A2(n_237),
.B1(n_246),
.B2(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_224),
.A2(n_246),
.B1(n_510),
.B2(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_226),
.Y(n_296)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AO21x2_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_247),
.B(n_253),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_230),
.Y(n_564)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_SL g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_257),
.B1(n_290),
.B2(n_296),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_246),
.A2(n_296),
.B1(n_336),
.B2(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_246),
.Y(n_436)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_246),
.A2(n_296),
.B(n_438),
.Y(n_636)
);

AOI21xp33_ASAP7_75t_SL g653 ( 
.A1(n_246),
.A2(n_296),
.B(n_438),
.Y(n_653)
);

NAND2xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_251),
.Y(n_486)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_251),
.Y(n_555)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_252),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_252),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_253),
.Y(n_568)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_260),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_270),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_270),
.Y(n_357)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_270),
.Y(n_503)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_270),
.Y(n_598)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_271),
.Y(n_532)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_273),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_287),
.C(n_289),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_289),
.Y(n_301)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_283),
.Y(n_518)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_290),
.A2(n_296),
.B1(n_478),
.B2(n_487),
.Y(n_477)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_296),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_296),
.B(n_326),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g463 ( 
.A(n_297),
.B(n_298),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_R g464 ( 
.A(n_297),
.B(n_298),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_327),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g608 ( 
.A(n_300),
.B(n_609),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_302),
.B(n_327),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_315),
.C(n_325),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_303),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_310),
.Y(n_498)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_315),
.A2(n_316),
.B1(n_325),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_325),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_326),
.B(n_491),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_326),
.B(n_496),
.C(n_498),
.Y(n_495)
);

OAI21xp33_ASAP7_75t_SL g549 ( 
.A1(n_326),
.A2(n_550),
.B(n_552),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_326),
.B(n_553),
.Y(n_552)
);

A2O1A1O1Ixp25_ASAP7_75t_L g612 ( 
.A1(n_329),
.A2(n_426),
.B(n_613),
.C(n_615),
.D(n_616),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_382),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_330),
.B(n_382),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.C(n_358),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_331),
.B(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_334),
.A2(n_359),
.B1(n_360),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_334),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_344),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g385 ( 
.A(n_335),
.B(n_344),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_350),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_353),
.Y(n_567)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_357),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_361),
.B2(n_381),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_359),
.B(n_363),
.C(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_361),
.B(n_467),
.Y(n_466)
);

AO21x1_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_371),
.B(n_380),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_371),
.Y(n_380)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_408),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_409),
.C(n_428),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_406),
.B2(n_407),
.Y(n_384)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_385),
.Y(n_407)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_388),
.B1(n_398),
.B2(n_399),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_407),
.C(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_424),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_414),
.B(n_423),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_SL g423 ( 
.A(n_410),
.B(n_415),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_410),
.A2(n_411),
.B1(n_455),
.B2(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_415),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_411),
.Y(n_668)
);

INVx8_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_416),
.Y(n_435)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

BUFx2_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_424),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_427),
.B(n_429),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_430),
.B(n_460),
.C(n_673),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_453),
.B1(n_459),
.B2(n_460),
.Y(n_432)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_446),
.B(n_452),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_446),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_437),
.B2(n_445),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_436),
.Y(n_487)
);

AOI22x1_ASAP7_75t_L g508 ( 
.A1(n_436),
.A2(n_445),
.B1(n_479),
.B2(n_509),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_436),
.A2(n_445),
.B1(n_537),
.B2(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_441),
.Y(n_551)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_447),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx8_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_452),
.Y(n_664)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_453),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_453),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_458),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_456),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_458),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_462),
.B(n_465),
.C(n_614),
.Y(n_613)
);

AOI21x1_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_607),
.B(n_611),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_521),
.B(n_606),
.Y(n_470)
);

NOR2x1_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_505),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_472),
.B(n_505),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_476),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_473),
.B(n_477),
.C(n_488),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_488),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_499),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_489),
.B(n_499),
.Y(n_506)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_494),
.Y(n_497)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_502),
.Y(n_592)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_503),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.C(n_514),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_506),
.B(n_541),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_508),
.A2(n_514),
.B(n_542),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_515),
.Y(n_543)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

AOI31xp67_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_544),
.A3(n_572),
.B(n_605),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_540),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_523),
.B(n_540),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_533),
.C(n_534),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_524),
.B(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g578 ( 
.A(n_529),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_531),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_533),
.B(n_535),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_571),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_569),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_546),
.B(n_569),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_556),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_557),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_547),
.A2(n_557),
.B(n_576),
.Y(n_604)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_548),
.B(n_556),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_551),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_552),
.Y(n_565)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_558),
.A2(n_565),
.B1(n_566),
.B2(n_568),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_559),
.B(n_563),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_573),
.C(n_585),
.Y(n_572)
);

AO21x1_ASAP7_75t_L g573 ( 
.A1(n_574),
.A2(n_575),
.B(n_577),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_577),
.B(n_604),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_603),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_587),
.A2(n_599),
.B(n_602),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_588),
.B(n_594),
.Y(n_587)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_595),
.B(n_596),
.Y(n_594)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_601),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_600),
.B(n_601),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_608),
.B(n_610),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g611 ( 
.A(n_608),
.B(n_610),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_660),
.C(n_680),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_619),
.A2(n_684),
.B(n_687),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_620),
.B(n_651),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_620),
.B(n_651),
.Y(n_687)
);

XNOR2xp5_ASAP7_75t_SL g620 ( 
.A(n_621),
.B(n_647),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_621),
.B(n_648),
.C(n_650),
.Y(n_681)
);

MAJx2_ASAP7_75t_L g621 ( 
.A(n_622),
.B(n_636),
.C(n_637),
.Y(n_621)
);

OA22x2_ASAP7_75t_L g658 ( 
.A1(n_622),
.A2(n_636),
.B1(n_653),
.B2(n_659),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_622),
.Y(n_659)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_628),
.Y(n_649)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_636),
.A2(n_653),
.B1(n_655),
.B2(n_671),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_637),
.B(n_658),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g679 ( 
.A(n_637),
.B(n_654),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_648),
.B(n_650),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_652),
.B(n_654),
.C(n_657),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_652),
.B(n_678),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_653),
.B(n_654),
.C(n_655),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_654),
.B(n_670),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_655),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g678 ( 
.A(n_658),
.B(n_679),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_661),
.B(n_674),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_672),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_662),
.B(n_672),
.Y(n_685)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_663),
.B(n_669),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_664),
.B(n_665),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_664),
.B(n_665),
.C(n_669),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_SL g665 ( 
.A1(n_666),
.A2(n_667),
.B1(n_668),
.B2(n_692),
.Y(n_665)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_675),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_675),
.A2(n_685),
.B(n_686),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_676),
.B(n_677),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_676),
.B(n_677),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_680),
.A2(n_683),
.B(n_688),
.Y(n_682)
);


endmodule