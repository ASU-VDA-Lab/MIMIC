module fake_jpeg_23492_n_41 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp33_ASAP7_75t_SL g7 ( 
.A(n_3),
.B(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_12),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

AND2x6_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_2),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_27),
.C(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_26),
.Y(n_31)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_6),
.C(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_8),
.A2(n_6),
.B(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_32),
.C(n_28),
.Y(n_39)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_38),
.A3(n_36),
.B1(n_32),
.B2(n_35),
.C1(n_30),
.C2(n_20),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_33),
.B(n_16),
.Y(n_41)
);


endmodule