module fake_jpeg_19216_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_11),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_1),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_1),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_8),
.B1(n_12),
.B2(n_10),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_27),
.B(n_1),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_31),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_8),
.B1(n_10),
.B2(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_12),
.B1(n_7),
.B2(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_31),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_26),
.C(n_29),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_32),
.B1(n_39),
.B2(n_28),
.Y(n_44)
);

AOI222xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_42),
.B1(n_43),
.B2(n_25),
.C1(n_35),
.C2(n_2),
.Y(n_45)
);


endmodule