module fake_jpeg_19118_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_34),
.B1(n_21),
.B2(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_55),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_52),
.A2(n_21),
.B1(n_17),
.B2(n_26),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_41),
.B1(n_37),
.B2(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_83),
.Y(n_117)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_55),
.B(n_50),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_85),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_24),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_89),
.B1(n_85),
.B2(n_17),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_79),
.B1(n_98),
.B2(n_60),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_34),
.B1(n_25),
.B2(n_35),
.Y(n_79)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_34),
.B1(n_43),
.B2(n_40),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_97),
.B1(n_52),
.B2(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_81),
.Y(n_131)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_86),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_43),
.C(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_60),
.B1(n_67),
.B2(n_63),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_48),
.B1(n_39),
.B2(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_102),
.A2(n_33),
.B1(n_22),
.B2(n_30),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_129),
.B1(n_80),
.B2(n_74),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_54),
.B1(n_24),
.B2(n_27),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_20),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_17),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_27),
.B1(n_35),
.B2(n_21),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_23),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_45),
.B1(n_39),
.B2(n_36),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_26),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_26),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_120),
.B1(n_111),
.B2(n_113),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_106),
.B1(n_133),
.B2(n_111),
.Y(n_178)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_154),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_152),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_93),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_139),
.A2(n_33),
.B(n_30),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_80),
.B1(n_69),
.B2(n_101),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_148),
.B1(n_160),
.B2(n_161),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_145),
.B1(n_153),
.B2(n_158),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_91),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_68),
.B1(n_92),
.B2(n_72),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_68),
.B1(n_72),
.B2(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_33),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_23),
.B1(n_95),
.B2(n_94),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_121),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_121),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_28),
.B1(n_33),
.B2(n_10),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_28),
.B1(n_33),
.B2(n_10),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_131),
.C(n_121),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_175),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_106),
.B1(n_120),
.B2(n_104),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_177),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_172),
.B(n_176),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_156),
.B(n_135),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_191),
.B(n_156),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_126),
.B(n_108),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_178),
.B(n_188),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_121),
.C(n_114),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_138),
.B(n_137),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_111),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_104),
.B1(n_122),
.B2(n_114),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_110),
.B1(n_32),
.B2(n_30),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_141),
.A2(n_122),
.B1(n_110),
.B2(n_119),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_33),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_133),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_187),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_108),
.B(n_105),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_105),
.B(n_1),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_136),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_201),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_196),
.A2(n_202),
.B(n_4),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_138),
.B(n_142),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_189),
.B(n_176),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

AOI21x1_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_158),
.B(n_142),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_110),
.B1(n_9),
.B2(n_11),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_205),
.B1(n_179),
.B2(n_185),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_208),
.B1(n_210),
.B2(n_169),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_32),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_207),
.A2(n_215),
.B(n_3),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_22),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_175),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_1),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_1),
.B(n_2),
.Y(n_215)
);

AO22x1_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_3),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_165),
.B1(n_177),
.B2(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_3),
.Y(n_241)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_233),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_228),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_163),
.C(n_164),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_164),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_199),
.C(n_198),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_237),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_250),
.B1(n_215),
.B2(n_203),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_209),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_238),
.A2(n_249),
.B(n_207),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_186),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_244),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_181),
.B1(n_191),
.B2(n_182),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_240),
.A2(n_205),
.B1(n_202),
.B2(n_214),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_241),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_248),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_181),
.C(n_11),
.Y(n_244)
);

AOI22x1_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_181),
.B1(n_4),
.B2(n_6),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_16),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_195),
.B(n_13),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_247),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_222),
.Y(n_248)
);

BUFx12f_ASAP7_75t_SL g254 ( 
.A(n_249),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

BUFx12f_ASAP7_75t_SL g257 ( 
.A(n_229),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_194),
.B(n_217),
.Y(n_278)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_223),
.B1(n_213),
.B2(n_210),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_240),
.B1(n_235),
.B2(n_244),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_227),
.B(n_196),
.Y(n_264)
);

OAI221xp5_ASAP7_75t_SL g282 ( 
.A1(n_264),
.A2(n_237),
.B1(n_239),
.B2(n_245),
.C(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_269),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_217),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_204),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_279),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_236),
.B1(n_194),
.B2(n_224),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_233),
.B1(n_250),
.B2(n_232),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_228),
.C(n_230),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_260),
.C(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_243),
.B1(n_238),
.B2(n_226),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_254),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_252),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_253),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_219),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_259),
.A2(n_221),
.B1(n_7),
.B2(n_8),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_267),
.B1(n_261),
.B2(n_258),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_256),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_293),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_292),
.B(n_305),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_285),
.C(n_287),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_270),
.C(n_251),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_301),
.C(n_304),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_251),
.C(n_262),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_271),
.C(n_266),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_272),
.C(n_281),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_314),
.C(n_317),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_301),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_298),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_281),
.C(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_277),
.C(n_289),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_297),
.A2(n_302),
.B1(n_294),
.B2(n_293),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_326),
.B(n_12),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_322),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_312),
.A2(n_277),
.B1(n_288),
.B2(n_299),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_291),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_308),
.B(n_11),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_12),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_310),
.B1(n_317),
.B2(n_314),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_329),
.Y(n_335)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_307),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_324),
.B(n_320),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_307),
.C(n_12),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_13),
.C(n_7),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_332),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_336),
.A2(n_337),
.B(n_338),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_328),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_335),
.B(n_337),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_333),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_13),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_8),
.C(n_6),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_6),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_7),
.Y(n_346)
);


endmodule