module fake_jpeg_21848_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_3),
.B(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_12),
.B(n_8),
.Y(n_19)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_15),
.A2(n_18),
.B1(n_0),
.B2(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_6),
.Y(n_16)
);

NOR2x1_ASAP7_75t_R g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_7),
.B1(n_10),
.B2(n_6),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_18),
.C(n_9),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_17),
.C(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_22),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.C(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_20),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_19),
.B1(n_15),
.B2(n_13),
.Y(n_34)
);


endmodule