module real_jpeg_4946_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_1),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_1),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_1),
.A2(n_123),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_1),
.A2(n_123),
.B1(n_195),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_1),
.A2(n_123),
.B1(n_167),
.B2(n_279),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_2),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_2),
.A2(n_193),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_2),
.A2(n_193),
.B1(n_410),
.B2(n_412),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_2),
.A2(n_193),
.B1(n_465),
.B2(n_470),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_4),
.A2(n_46),
.B1(n_92),
.B2(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_4),
.A2(n_46),
.B1(n_52),
.B2(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_4),
.A2(n_46),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_274),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_5),
.A2(n_273),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_5),
.B(n_198),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_5),
.B(n_43),
.C(n_383),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g386 ( 
.A1(n_5),
.A2(n_387),
.B1(n_388),
.B2(n_390),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_5),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_5),
.B(n_144),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_5),
.A2(n_32),
.B1(n_431),
.B2(n_434),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_6),
.A2(n_264),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_6),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_6),
.A2(n_292),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_6),
.A2(n_292),
.B1(n_394),
.B2(n_397),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_6),
.A2(n_292),
.B1(n_415),
.B2(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_7),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_7),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_7),
.A2(n_297),
.B1(n_328),
.B2(n_332),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_7),
.A2(n_297),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_7),
.A2(n_166),
.B1(n_297),
.B2(n_421),
.Y(n_420)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_9),
.Y(n_313)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_9),
.Y(n_348)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_9),
.Y(n_436)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_10),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_10),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_83),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_10),
.A2(n_83),
.B1(n_166),
.B2(n_171),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_10),
.A2(n_83),
.B1(n_124),
.B2(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_13),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_13),
.Y(n_217)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_13),
.Y(n_246)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_14),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_17),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_17),
.A2(n_50),
.B1(n_146),
.B2(n_150),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_17),
.A2(n_50),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_17),
.A2(n_50),
.B1(n_284),
.B2(n_287),
.Y(n_283)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_512),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_502),
.B(n_511),
.Y(n_25)
);

OAI31xp33_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_222),
.A3(n_247),
.B(n_499),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_204),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_28),
.B(n_204),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_117),
.C(n_160),
.Y(n_28)
);

FAx1_ASAP7_75t_L g373 ( 
.A(n_29),
.B(n_117),
.CI(n_160),
.CON(n_373),
.SN(n_373)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_86),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_30),
.A2(n_31),
.B(n_88),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_47),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_31),
.A2(n_87),
.B1(n_88),
.B2(n_116),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_31),
.A2(n_47),
.B1(n_87),
.B2(n_365),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_38),
.B(n_40),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_32),
.B(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_32),
.A2(n_277),
.B1(n_282),
.B2(n_283),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_32),
.A2(n_283),
.B(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_32),
.A2(n_174),
.B(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_32),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_32),
.A2(n_420),
.B1(n_431),
.B2(n_434),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_32),
.A2(n_40),
.B(n_312),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_35),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_37),
.Y(n_425)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_70)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_47),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_60),
.B(n_76),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_49),
.A2(n_61),
.B1(n_77),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_54),
.Y(n_396)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_54),
.Y(n_453)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_55),
.Y(n_469)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_56),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_56),
.Y(n_389)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_56),
.Y(n_392)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_59),
.A2(n_127),
.B1(n_129),
.B2(n_132),
.Y(n_126)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_60),
.B(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_60),
.A2(n_78),
.B(n_154),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_60),
.A2(n_78),
.B1(n_158),
.B2(n_182),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_60),
.A2(n_76),
.B(n_154),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_60),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_61),
.A2(n_77),
.B1(n_386),
.B2(n_393),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_61),
.A2(n_77),
.B1(n_393),
.B2(n_404),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_61),
.A2(n_77),
.B1(n_404),
.B2(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_62)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_63),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_69),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_73),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_73),
.Y(n_411)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_73),
.Y(n_415)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_75),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_78),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_78),
.B(n_387),
.Y(n_429)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_82),
.Y(n_405)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_85),
.Y(n_184)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_107),
.B(n_109),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_89),
.B(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_89),
.A2(n_198),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_89),
.A2(n_198),
.B1(n_289),
.B2(n_293),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_90),
.A2(n_190),
.B(n_197),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_90),
.A2(n_115),
.B1(n_190),
.B2(n_294),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_90),
.A2(n_115),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_90),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_91)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_99),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_102),
.Y(n_263)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_103),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_103),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_109),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_112),
.Y(n_296)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_114),
.Y(n_299)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_115),
.A2(n_215),
.B(n_218),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_152),
.B(n_159),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_152),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_125),
.B1(n_144),
.B2(n_145),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_120),
.A2(n_126),
.B(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_121),
.Y(n_255)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_125),
.B(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_125),
.A2(n_145),
.B(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_125),
.A2(n_233),
.B(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_125),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_125),
.A2(n_144),
.B1(n_353),
.B2(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_125),
.A2(n_144),
.B(n_506),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_134),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_126),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_126),
.A2(n_307),
.B1(n_327),
.B2(n_335),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_126),
.A2(n_307),
.B1(n_327),
.B2(n_352),
.Y(n_351)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_129),
.Y(n_454)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_131),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_140),
.B2(n_143),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_144),
.B(n_202),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_SL g462 ( 
.A1(n_146),
.A2(n_387),
.B(n_455),
.Y(n_462)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_148),
.Y(n_354)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_153),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_159),
.B(n_205),
.CI(n_221),
.CON(n_204),
.SN(n_204)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_188),
.C(n_199),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_161),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_179),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_162),
.A2(n_179),
.B1(n_180),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_162),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_164),
.A2(n_278),
.B(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_165),
.Y(n_314)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_168),
.Y(n_433)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_169),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_170),
.Y(n_286)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_172),
.B(n_440),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_178),
.Y(n_282)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_188),
.A2(n_189),
.B1(n_199),
.B2(n_200),
.Y(n_367)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_197),
.B(n_218),
.Y(n_514)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_204),
.B(n_224),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_214),
.B2(n_220),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_213),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_208),
.B(n_230),
.C(n_240),
.Y(n_510)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_213),
.C(n_214),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_211),
.A2(n_234),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_220),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_214),
.B(n_225),
.C(n_228),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_216),
.Y(n_264)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_223),
.A2(n_500),
.B(n_501),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_240),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_234),
.Y(n_506)
);

INVx8_ASAP7_75t_L g450 ( 
.A(n_235),
.Y(n_450)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_239),
.Y(n_331)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_239),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_242),
.Y(n_508)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_374),
.B(n_493),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_359),
.C(n_371),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_337),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_250),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_316),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_251),
.B(n_316),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_300),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_252),
.B(n_301),
.C(n_303),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.C(n_288),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_253),
.B(n_288),
.Y(n_318)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_254),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_259),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_276),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_260),
.B(n_276),
.Y(n_340)
);

OAI32xp33_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_264),
.A3(n_265),
.B1(n_269),
.B2(n_272),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g356 ( 
.A(n_263),
.Y(n_356)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_281),
.Y(n_421)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_305),
.B(n_309),
.C(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_315),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.C(n_336),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_336),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.C(n_326),
.Y(n_319)
);

FAx1_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_321),
.CI(n_326),
.CON(n_339),
.SN(n_339)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_332),
.B(n_387),
.Y(n_455)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_357),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_338),
.B(n_357),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.C(n_341),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_339),
.B(n_491),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_339),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_340),
.B(n_341),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_349),
.C(n_351),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_342),
.A2(n_343),
.B1(n_349),
.B2(n_350),
.Y(n_478)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_345),
.B(n_387),
.Y(n_440)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_351),
.B(n_478),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

A2O1A1O1Ixp25_ASAP7_75t_L g493 ( 
.A1(n_359),
.A2(n_371),
.B(n_494),
.C(n_497),
.D(n_498),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_370),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_360),
.B(n_370),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_364),
.C(n_369),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_366),
.B1(n_368),
.B2(n_369),
.Y(n_363)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_364),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_366),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_372),
.B(n_373),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g519 ( 
.A(n_373),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_488),
.B(n_492),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_473),
.B(n_487),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_444),
.B(n_472),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_416),
.B(n_443),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_399),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_379),
.B(n_399),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_385),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_385),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_408),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_403),
.B2(n_407),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_407),
.C(n_408),
.Y(n_445)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_403),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_406),
.B(n_457),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_427),
.B(n_442),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_426),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_426),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_422),
.B1(n_423),
.B2(n_424),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_437),
.B(n_441),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_429),
.B(n_430),
.Y(n_441)
);

INVx4_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_446),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_460),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_461),
.C(n_463),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_459),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_459),
.Y(n_481)
);

OAI32xp33_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_451),
.A3(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_475),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_479),
.B2(n_480),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_482),
.C(n_485),
.Y(n_489)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_481),
.A2(n_482),
.B1(n_485),
.B2(n_486),
.Y(n_480)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_481),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_482),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_489),
.B(n_490),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_503),
.B(n_504),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_504),
.B(n_514),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_504),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g504 ( 
.A(n_505),
.B(n_507),
.CI(n_510),
.CON(n_504),
.SN(n_504)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_515),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_514),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);


endmodule