module real_jpeg_11898_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_200),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_200),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_3),
.A2(n_43),
.B1(n_48),
.B2(n_200),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_4),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_4),
.A2(n_33),
.B1(n_35),
.B2(n_173),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_4),
.A2(n_43),
.B1(n_48),
.B2(n_173),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_6),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_6),
.A2(n_59),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_6),
.B(n_83),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_6),
.B(n_28),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_6),
.A2(n_33),
.B1(n_35),
.B2(n_192),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_6),
.A2(n_35),
.B(n_47),
.C(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_6),
.B(n_74),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_6),
.B(n_100),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_6),
.B(n_41),
.Y(n_290)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_6),
.A2(n_28),
.B(n_249),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_7),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_108),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_108),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_7),
.A2(n_43),
.B1(n_48),
.B2(n_108),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_8),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_8),
.A2(n_37),
.B1(n_43),
.B2(n_48),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_68),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_10),
.A2(n_43),
.B1(n_48),
.B2(n_68),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_12),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_145),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_145),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_12),
.A2(n_43),
.B1(n_48),
.B2(n_145),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_13),
.A2(n_33),
.B1(n_35),
.B2(n_63),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_43),
.B1(n_48),
.B2(n_63),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_15),
.A2(n_39),
.B1(n_43),
.B2(n_48),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_16),
.A2(n_33),
.B1(n_35),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_16),
.A2(n_43),
.B1(n_48),
.B2(n_65),
.Y(n_164)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_75),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_75),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.C(n_69),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_22),
.A2(n_66),
.B1(n_116),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_22),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_52),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_25),
.B(n_40),
.C(n_53),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_25)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_26),
.A2(n_32),
.B1(n_113),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_26),
.A2(n_32),
.B1(n_142),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_26),
.A2(n_32),
.B1(n_195),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_26),
.A2(n_32),
.B1(n_224),
.B2(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_28),
.A2(n_29),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_28),
.B(n_56),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_28),
.A2(n_30),
.A3(n_33),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_29),
.A2(n_57),
.A3(n_59),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_31),
.B(n_35),
.Y(n_250)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_66),
.C(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_40),
.A2(n_52),
.B1(n_70),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B(n_51),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_41),
.A2(n_49),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_41),
.A2(n_49),
.B1(n_51),
.B2(n_105),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_41),
.A2(n_49),
.B1(n_104),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_41),
.A2(n_49),
.B1(n_167),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_41),
.A2(n_49),
.B1(n_216),
.B2(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_41),
.A2(n_49),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_41),
.A2(n_49),
.B1(n_264),
.B2(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_42),
.A2(n_140),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_42),
.A2(n_168),
.B1(n_243),
.B2(n_301),
.Y(n_300)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_42)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_43),
.B(n_287),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_46),
.A2(n_48),
.B(n_192),
.Y(n_266)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_49),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_54),
.A2(n_55),
.B1(n_67),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_54),
.A2(n_55),
.B1(n_107),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_54),
.A2(n_55),
.B1(n_144),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_54),
.A2(n_55),
.B1(n_199),
.B2(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_60),
.B(n_192),
.Y(n_191)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_74),
.B(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_72),
.A2(n_74),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_72),
.A2(n_74),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_86),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_81),
.A2(n_83),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_151),
.B(n_321),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_146),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_122),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_92),
.B(n_122),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_109),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_115),
.C(n_120),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B(n_106),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_95),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_97),
.B1(n_106),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_98),
.A2(n_100),
.B1(n_164),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_98),
.A2(n_100),
.B1(n_188),
.B2(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_98),
.A2(n_100),
.B1(n_228),
.B2(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_98),
.A2(n_100),
.B1(n_252),
.B2(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_98),
.A2(n_100),
.B1(n_192),
.B2(n_285),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_98),
.A2(n_100),
.B1(n_278),
.B2(n_285),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_99),
.A2(n_136),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_99),
.A2(n_162),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_111),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.C(n_130),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_141),
.C(n_143),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_132),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_146),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_147),
.B(n_148),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_176),
.B(n_320),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_174),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_153),
.B(n_174),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_158),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_169),
.C(n_171),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_160),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_161),
.B(n_165),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_171),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_204),
.B(n_319),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_202),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_178),
.B(n_202),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_184),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_183),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_184),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_193),
.C(n_197),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_197),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_235),
.B(n_313),
.C(n_318),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_229),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_206),
.B(n_229),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_219),
.C(n_221),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_207),
.A2(n_208),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_213),
.C(n_218),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_221),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_227),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_231),
.B(n_232),
.C(n_233),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_312),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_256),
.B(n_311),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_253),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_238),
.B(n_253),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_244),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_241),
.A2(n_244),
.B1(n_245),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_251),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_246),
.A2(n_247),
.B1(n_251),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_305),
.B(n_310),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_294),
.B(n_304),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_274),
.B(n_293),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_260),
.B(n_267),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_270),
.C(n_272),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_273),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_282),
.B(n_292),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_280),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_288),
.B(n_291),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_296),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_300),
.C(n_302),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);


endmodule