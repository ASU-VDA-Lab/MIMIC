module fake_netlist_1_12754_n_720 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_720);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_720;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g106 ( .A(n_79), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_91), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_81), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_24), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_22), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_92), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_63), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_56), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_32), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_54), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_19), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_102), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_42), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_93), .Y(n_119) );
BUFx8_ASAP7_75t_SL g120 ( .A(n_105), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_86), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_57), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_60), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_62), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_48), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_41), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_77), .Y(n_128) );
BUFx10_ASAP7_75t_L g129 ( .A(n_23), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_7), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_88), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_18), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_53), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_1), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_17), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_19), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_65), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_66), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_38), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_39), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_68), .Y(n_143) );
CKINVDCx14_ASAP7_75t_R g144 ( .A(n_5), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_76), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_45), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_26), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_16), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_114), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_117), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_129), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_129), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_135), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_106), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_129), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
AOI22x1_ASAP7_75t_SL g164 ( .A1(n_110), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_137), .B(n_0), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_108), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_110), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_131), .B(n_3), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_162), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_154), .B(n_112), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_153), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_163), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_154), .B(n_116), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_151), .B(n_109), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_151), .B(n_115), .Y(n_182) );
BUFx10_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
INVxp33_ASAP7_75t_L g186 ( .A(n_165), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_154), .B(n_121), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
BUFx8_ASAP7_75t_SL g190 ( .A(n_155), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_156), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_155), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_157), .B(n_123), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_177), .A2(n_167), .B1(n_157), .B2(n_166), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_192), .B(n_155), .Y(n_196) );
INVx5_ASAP7_75t_L g197 ( .A(n_177), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_170), .B(n_155), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_186), .B(n_161), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_179), .B(n_168), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_185), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_179), .B(n_159), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_170), .B(n_159), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_183), .B(n_107), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_185), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_183), .B(n_107), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_183), .B(n_113), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_188), .B(n_159), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_180), .B(n_166), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_183), .B(n_113), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_180), .B(n_166), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_194), .A2(n_162), .B(n_139), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_182), .B(n_118), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_177), .A2(n_122), .B1(n_133), .B2(n_152), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_177), .A2(n_167), .B1(n_164), .B2(n_111), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_175), .B(n_118), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_175), .B(n_136), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_182), .B(n_125), .Y(n_218) );
NOR3xp33_ASAP7_75t_L g219 ( .A(n_194), .B(n_136), .C(n_138), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_181), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_177), .A2(n_164), .B1(n_126), .B2(n_132), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_177), .B(n_125), .Y(n_222) );
NOR2xp33_ASAP7_75t_SL g223 ( .A(n_175), .B(n_147), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_169), .A2(n_152), .B1(n_158), .B2(n_160), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_181), .A2(n_138), .B1(n_149), .B2(n_140), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_175), .B(n_128), .Y(n_227) );
NOR3xp33_ASAP7_75t_SL g228 ( .A(n_190), .B(n_149), .C(n_134), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_169), .B(n_128), .Y(n_229) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_223), .B(n_193), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_217), .A2(n_169), .B1(n_191), .B2(n_187), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_220), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_198), .B(n_187), .Y(n_234) );
NAND2x1_ASAP7_75t_L g235 ( .A(n_220), .B(n_191), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_197), .B(n_193), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_197), .A2(n_189), .B1(n_184), .B2(n_140), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_198), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_198), .B(n_184), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_197), .B(n_185), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_203), .A2(n_171), .B(n_172), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_198), .B(n_158), .Y(n_242) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_222), .B(n_184), .Y(n_243) );
AOI22x1_ASAP7_75t_L g244 ( .A1(n_201), .A2(n_185), .B1(n_189), .B2(n_176), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_199), .A2(n_178), .B(n_176), .C(n_171), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_217), .A2(n_134), .B1(n_145), .B2(n_189), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_209), .A2(n_160), .B(n_124), .C(n_146), .Y(n_247) );
OR2x6_ASAP7_75t_L g248 ( .A(n_216), .B(n_127), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_225), .B(n_185), .Y(n_249) );
OA22x2_ASAP7_75t_L g250 ( .A1(n_215), .A2(n_145), .B1(n_130), .B2(n_141), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_201), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_208), .A2(n_172), .B(n_174), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_211), .A2(n_174), .B(n_173), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_200), .B(n_120), .Y(n_254) );
NOR2xp67_ASAP7_75t_SL g255 ( .A(n_197), .B(n_142), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_213), .B(n_143), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_218), .B(n_148), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_202), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_229), .A2(n_173), .B(n_176), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_195), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_244), .A2(n_205), .B(n_226), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_242), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_259), .A2(n_197), .B(n_196), .Y(n_264) );
O2A1O1Ixp5_ASAP7_75t_SL g265 ( .A1(n_260), .A2(n_178), .B(n_212), .C(n_210), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_236), .Y(n_266) );
AO31x2_ASAP7_75t_L g267 ( .A1(n_233), .A2(n_205), .A3(n_226), .B(n_195), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_258), .B(n_225), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_252), .A2(n_224), .B(n_214), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_241), .A2(n_219), .B(n_204), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_247), .A2(n_215), .B(n_221), .C(n_178), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_245), .A2(n_207), .B(n_206), .C(n_227), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_253), .A2(n_178), .B(n_221), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_235), .A2(n_50), .B(n_104), .Y(n_274) );
AO21x1_ASAP7_75t_L g275 ( .A1(n_247), .A2(n_4), .B(n_5), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_245), .A2(n_51), .B(n_103), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_238), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_232), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_251), .A2(n_49), .B(n_101), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_251), .A2(n_47), .B(n_100), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_239), .A2(n_228), .B(n_46), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_230), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_230), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_277), .Y(n_285) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_276), .A2(n_257), .B(n_256), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_267), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_268), .B(n_231), .Y(n_288) );
CKINVDCx6p67_ASAP7_75t_R g289 ( .A(n_278), .Y(n_289) );
AO31x2_ASAP7_75t_L g290 ( .A1(n_275), .A2(n_234), .A3(n_237), .B(n_254), .Y(n_290) );
AOI21xp33_ASAP7_75t_L g291 ( .A1(n_284), .A2(n_250), .B(n_249), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_278), .B(n_232), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_262), .B(n_243), .Y(n_293) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_274), .A2(n_240), .B(n_246), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_267), .Y(n_295) );
AND2x6_ASAP7_75t_L g296 ( .A(n_282), .B(n_232), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_265), .A2(n_240), .B(n_250), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_272), .A2(n_243), .B(n_248), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_267), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_274), .A2(n_255), .B(n_248), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_261), .A2(n_232), .B(n_248), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_267), .Y(n_302) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_275), .A2(n_44), .B(n_98), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_263), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_261), .A2(n_43), .B(n_97), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_292), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_295), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_287), .B(n_271), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_301), .A2(n_281), .B(n_270), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_289), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_301), .A2(n_280), .B(n_279), .Y(n_311) );
AO31x2_ASAP7_75t_L g312 ( .A1(n_287), .A2(n_271), .A3(n_273), .B(n_264), .Y(n_312) );
AO31x2_ASAP7_75t_L g313 ( .A1(n_302), .A2(n_272), .A3(n_269), .B(n_9), .Y(n_313) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_301), .A2(n_269), .B(n_283), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_302), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_295), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_295), .B(n_266), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_299), .B(n_6), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_289), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_299), .B(n_8), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_285), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_288), .B(n_10), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_296), .B(n_55), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_305), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_289), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
OAI21xp5_ASAP7_75t_SL g332 ( .A1(n_298), .A2(n_10), .B(n_11), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_307), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_307), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_315), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_316), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_308), .B(n_303), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_330), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_308), .B(n_303), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_330), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_308), .B(n_303), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_319), .B(n_303), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_319), .B(n_303), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_319), .B(n_303), .Y(n_345) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_327), .B(n_304), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_319), .B(n_290), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_316), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_330), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_317), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_317), .Y(n_352) );
INVx4_ASAP7_75t_L g353 ( .A(n_330), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_323), .B(n_305), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_331), .B(n_288), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_323), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_327), .B(n_290), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_314), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_318), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_306), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_314), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_306), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_326), .A2(n_296), .B1(n_298), .B2(n_294), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_310), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_314), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_326), .A2(n_296), .B1(n_288), .B2(n_291), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_318), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_325), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_314), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_320), .B(n_290), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_377), .B(n_320), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_377), .B(n_320), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_377), .B(n_322), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_347), .B(n_322), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_361), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_353), .Y(n_384) );
INVx4_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_347), .B(n_322), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_312), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_361), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_358), .B(n_312), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_336), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_335), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_342), .B(n_331), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_347), .B(n_314), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_362), .B(n_312), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_359), .B(n_327), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_342), .B(n_325), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_348), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_362), .B(n_312), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_348), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_360), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_365), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_363), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_374), .B(n_312), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_370), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_370), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_374), .B(n_312), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_375), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_365), .Y(n_413) );
AND2x4_ASAP7_75t_SL g414 ( .A(n_353), .B(n_310), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_375), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_336), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_333), .B(n_312), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_359), .B(n_312), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_359), .B(n_313), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_350), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_333), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_359), .B(n_313), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_359), .B(n_327), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_355), .B(n_333), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_350), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_356), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_334), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_334), .B(n_326), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_351), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_357), .B(n_313), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_357), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_368), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_351), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_352), .B(n_313), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_371), .B(n_321), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_337), .B(n_313), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_340), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_368), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_337), .B(n_313), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_337), .B(n_313), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_352), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_356), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_339), .B(n_313), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_385), .B(n_353), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_414), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_425), .B(n_339), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_379), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_385), .B(n_353), .Y(n_450) );
AOI32xp33_ASAP7_75t_L g451 ( .A1(n_414), .A2(n_371), .A3(n_346), .B1(n_349), .B2(n_338), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_430), .B(n_356), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_433), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_430), .B(n_356), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_390), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_379), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_382), .B(n_346), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_425), .B(n_332), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_391), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_385), .B(n_338), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_397), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_382), .B(n_346), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_397), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_399), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_394), .B(n_339), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_399), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_439), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_394), .B(n_341), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_386), .B(n_355), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_398), .B(n_341), .Y(n_472) );
AND2x4_ASAP7_75t_SL g473 ( .A(n_385), .B(n_306), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_386), .B(n_346), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_398), .B(n_341), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_392), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_378), .B(n_364), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_414), .B(n_340), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_429), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_407), .B(n_368), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_378), .B(n_364), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_420), .A2(n_373), .B1(n_296), .B2(n_367), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_407), .B(n_372), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_380), .B(n_366), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_380), .B(n_366), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_381), .B(n_366), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_384), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_392), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_381), .B(n_364), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_411), .B(n_366), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_429), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_416), .B(n_338), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_437), .B(n_332), .C(n_291), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_400), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_384), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_395), .B(n_338), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_426), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_429), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_428), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_416), .B(n_349), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_411), .B(n_372), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_387), .B(n_349), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_400), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_419), .B(n_349), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_402), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_383), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_419), .B(n_373), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_428), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_402), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_404), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_404), .Y(n_511) );
NAND2x1_ASAP7_75t_L g512 ( .A(n_395), .B(n_327), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_405), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_405), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_383), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_395), .B(n_367), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_393), .B(n_372), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_383), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_406), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_393), .B(n_376), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_395), .B(n_343), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_406), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_408), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_439), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_408), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_417), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_424), .B(n_343), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_424), .B(n_343), .Y(n_528) );
AOI21x1_ASAP7_75t_SL g529 ( .A1(n_424), .A2(n_344), .B(n_345), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_476), .B(n_438), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_446), .B(n_424), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_517), .B(n_387), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_488), .B(n_438), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_448), .B(n_441), .Y(n_534) );
AOI32xp33_ASAP7_75t_L g535 ( .A1(n_450), .A2(n_423), .A3(n_420), .B1(n_445), .B2(n_442), .Y(n_535) );
NAND2x2_ASAP7_75t_L g536 ( .A(n_447), .B(n_389), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_448), .B(n_441), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_455), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_493), .B(n_306), .C(n_297), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_504), .B(n_423), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_506), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_449), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_467), .B(n_442), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_459), .B(n_445), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_484), .B(n_428), .Y(n_545) );
NAND2x1_ASAP7_75t_SL g546 ( .A(n_446), .B(n_428), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_467), .B(n_389), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_456), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_470), .B(n_421), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_458), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_517), .B(n_417), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_460), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_485), .B(n_432), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_463), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_520), .B(n_388), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_470), .B(n_421), .Y(n_556) );
INVxp33_ASAP7_75t_L g557 ( .A(n_450), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_459), .A2(n_396), .B1(n_443), .B2(n_427), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_472), .B(n_427), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_465), .Y(n_560) );
NAND3xp33_ASAP7_75t_SL g561 ( .A(n_451), .B(n_432), .C(n_436), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_506), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_486), .B(n_444), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_466), .Y(n_564) );
OAI31xp33_ASAP7_75t_L g565 ( .A1(n_493), .A2(n_444), .A3(n_443), .B(n_435), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_457), .B(n_409), .Y(n_566) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_478), .B(n_431), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_468), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_487), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_471), .B(n_396), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_462), .B(n_409), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_516), .A2(n_296), .B1(n_306), .B2(n_436), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_464), .B(n_410), .Y(n_573) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_461), .B(n_297), .C(n_410), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_520), .B(n_388), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_512), .A2(n_435), .B1(n_431), .B2(n_415), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_453), .Y(n_577) );
OAI31xp33_ASAP7_75t_L g578 ( .A1(n_473), .A2(n_412), .A3(n_415), .B(n_344), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_474), .B(n_412), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_490), .B(n_388), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_472), .B(n_401), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_521), .B(n_401), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_494), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_503), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_527), .B(n_401), .Y(n_585) );
NAND4xp25_ASAP7_75t_L g586 ( .A(n_482), .B(n_293), .C(n_344), .D(n_345), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_528), .B(n_403), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_461), .B(n_440), .C(n_434), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_505), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
NAND2xp33_ASAP7_75t_SL g591 ( .A(n_462), .B(n_403), .Y(n_591) );
AOI32xp33_ASAP7_75t_L g592 ( .A1(n_507), .A2(n_345), .A3(n_434), .B1(n_418), .B2(n_413), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_495), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_496), .B(n_403), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_509), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_510), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_475), .B(n_413), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_511), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_496), .B(n_413), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_477), .B(n_434), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_513), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_526), .A2(n_296), .B(n_297), .Y(n_603) );
O2A1O1Ixp5_ASAP7_75t_R g604 ( .A1(n_480), .A2(n_293), .B(n_12), .C(n_13), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_514), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_519), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_558), .B(n_526), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_540), .B(n_524), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_555), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_586), .A2(n_482), .B1(n_489), .B2(n_481), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_569), .B(n_469), .Y(n_612) );
AOI322xp5_ASAP7_75t_L g613 ( .A1(n_604), .A2(n_475), .A3(n_497), .B1(n_501), .B2(n_480), .C1(n_483), .C2(n_469), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_SL g614 ( .A1(n_539), .A2(n_508), .B(n_491), .C(n_498), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_532), .B(n_483), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_544), .B(n_497), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_577), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_593), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_545), .B(n_501), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_551), .B(n_502), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_558), .B(n_522), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_549), .Y(n_622) );
OAI322xp33_ASAP7_75t_L g623 ( .A1(n_547), .A2(n_452), .A3(n_454), .B1(n_500), .B2(n_492), .C1(n_525), .C2(n_523), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_578), .B(n_499), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_557), .A2(n_518), .B(n_508), .C(n_479), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_582), .B(n_499), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_547), .B(n_440), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_549), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_567), .B(n_300), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_536), .A2(n_529), .B1(n_440), .B2(n_418), .Y(n_630) );
NOR2xp33_ASAP7_75t_R g631 ( .A(n_591), .B(n_11), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_585), .B(n_587), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_581), .B(n_418), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_556), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_546), .A2(n_529), .B(n_354), .C(n_376), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_581), .B(n_376), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_561), .B(n_311), .C(n_329), .Y(n_637) );
AOI21xp33_ASAP7_75t_L g638 ( .A1(n_565), .A2(n_12), .B(n_13), .Y(n_638) );
AOI321xp33_ASAP7_75t_L g639 ( .A1(n_574), .A2(n_354), .A3(n_329), .B1(n_328), .B2(n_296), .C(n_290), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_556), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_598), .B(n_575), .Y(n_641) );
OAI321xp33_ASAP7_75t_L g642 ( .A1(n_535), .A2(n_292), .A3(n_328), .B1(n_329), .B2(n_296), .C(n_290), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_598), .B(n_543), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_543), .B(n_290), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_559), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_534), .B(n_290), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_559), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g648 ( .A1(n_576), .A2(n_354), .A3(n_328), .B1(n_311), .B2(n_296), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_586), .A2(n_354), .B(n_15), .C(n_16), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_597), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_592), .A2(n_354), .B1(n_15), .B2(n_17), .C(n_18), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_534), .B(n_309), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_570), .A2(n_14), .B1(n_20), .B2(n_21), .C(n_22), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_542), .Y(n_654) );
XOR2x2_ASAP7_75t_L g655 ( .A(n_531), .B(n_14), .Y(n_655) );
AOI222xp33_ASAP7_75t_L g656 ( .A1(n_530), .A2(n_296), .B1(n_311), .B2(n_290), .C1(n_20), .C2(n_21), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_612), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_624), .A2(n_649), .B(n_613), .C(n_625), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_608), .B(n_537), .Y(n_659) );
OAI322xp33_ASAP7_75t_L g660 ( .A1(n_616), .A2(n_537), .A3(n_533), .B1(n_530), .B2(n_602), .C1(n_548), .C2(n_550), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_622), .B(n_533), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_626), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_611), .A2(n_571), .B1(n_531), .B2(n_594), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_649), .A2(n_588), .B(n_571), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g665 ( .A1(n_637), .A2(n_553), .A3(n_579), .B1(n_566), .B2(n_573), .C1(n_580), .C2(n_563), .Y(n_665) );
AOI21xp5_ASAP7_75t_R g666 ( .A1(n_630), .A2(n_603), .B(n_572), .Y(n_666) );
OA21x2_ASAP7_75t_SL g667 ( .A1(n_618), .A2(n_603), .B(n_600), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_610), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_623), .A2(n_606), .B1(n_605), .B2(n_552), .C(n_599), .Y(n_669) );
OAI31xp33_ASAP7_75t_L g670 ( .A1(n_614), .A2(n_584), .A3(n_596), .B(n_595), .Y(n_670) );
AOI322xp5_ASAP7_75t_L g671 ( .A1(n_621), .A2(n_601), .A3(n_560), .B1(n_589), .B2(n_583), .C1(n_568), .C2(n_564), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_628), .B(n_554), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_638), .A2(n_562), .B(n_541), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_623), .A2(n_590), .B(n_300), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g675 ( .A1(n_631), .A2(n_309), .B(n_300), .C(n_294), .Y(n_675) );
AOI32xp33_ASAP7_75t_L g676 ( .A1(n_625), .A2(n_300), .A3(n_309), .B1(n_294), .B2(n_292), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_648), .A2(n_309), .B1(n_300), .B2(n_292), .C(n_294), .Y(n_677) );
AOI31xp33_ASAP7_75t_L g678 ( .A1(n_651), .A2(n_309), .A3(n_300), .B(n_294), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_639), .A2(n_309), .B1(n_294), .B2(n_286), .C(n_29), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_642), .A2(n_25), .B1(n_27), .B2(n_28), .C(n_31), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_634), .B(n_286), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_641), .B(n_286), .Y(n_682) );
AOI21xp33_ASAP7_75t_SL g683 ( .A1(n_656), .A2(n_33), .B(n_34), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_655), .A2(n_286), .B(n_36), .Y(n_684) );
NOR4xp25_ASAP7_75t_SL g685 ( .A(n_607), .B(n_286), .C(n_37), .D(n_40), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_640), .A2(n_35), .B1(n_52), .B2(n_58), .C(n_59), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_643), .B(n_286), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_646), .A2(n_61), .B(n_64), .C(n_67), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_645), .A2(n_69), .B1(n_70), .B2(n_71), .C(n_72), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_635), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_639), .B(n_80), .C(n_82), .Y(n_691) );
NAND4xp25_ASAP7_75t_L g692 ( .A(n_653), .B(n_84), .C(n_85), .D(n_87), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_629), .A2(n_89), .B1(n_90), .B2(n_94), .Y(n_693) );
NAND2x1_ASAP7_75t_L g694 ( .A(n_609), .B(n_99), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_620), .A2(n_95), .B1(n_96), .B2(n_615), .Y(n_695) );
AOI222xp33_ASAP7_75t_L g696 ( .A1(n_644), .A2(n_647), .B1(n_654), .B2(n_617), .C1(n_627), .C2(n_619), .Y(n_696) );
OAI21xp5_ASAP7_75t_L g697 ( .A1(n_629), .A2(n_636), .B(n_652), .Y(n_697) );
CKINVDCx16_ASAP7_75t_R g698 ( .A(n_695), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_696), .B(n_671), .Y(n_699) );
NOR4xp75_ASAP7_75t_L g700 ( .A(n_664), .B(n_660), .C(n_694), .D(n_666), .Y(n_700) );
NOR4xp25_ASAP7_75t_L g701 ( .A(n_658), .B(n_669), .C(n_657), .D(n_667), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_670), .A2(n_683), .B(n_673), .C(n_684), .Y(n_702) );
AOI211x1_ASAP7_75t_SL g703 ( .A1(n_691), .A2(n_697), .B(n_659), .C(n_692), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_668), .A2(n_678), .B1(n_674), .B2(n_663), .C(n_677), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g705 ( .A(n_698), .B(n_690), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_702), .B(n_680), .C(n_693), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_699), .B(n_675), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g708 ( .A(n_704), .B(n_686), .C(n_689), .Y(n_708) );
AND3x1_ASAP7_75t_L g709 ( .A(n_706), .B(n_701), .C(n_700), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_707), .B(n_662), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_708), .B(n_672), .Y(n_711) );
XNOR2xp5_ASAP7_75t_L g712 ( .A(n_709), .B(n_703), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_710), .A2(n_705), .B1(n_679), .B2(n_682), .Y(n_713) );
INVx4_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_713), .A2(n_711), .B1(n_710), .B2(n_688), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_711), .B1(n_661), .B2(n_687), .Y(n_716) );
OAI222xp33_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_714), .B1(n_711), .B2(n_676), .C1(n_650), .C2(n_665), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_711), .B(n_678), .Y(n_718) );
AO21x1_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_681), .B(n_632), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_685), .B(n_633), .Y(n_720) );
endmodule