module real_jpeg_24216_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_0),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_0),
.B(n_53),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_0),
.B(n_50),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_0),
.B(n_32),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_0),
.B(n_17),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_0),
.B(n_48),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_0),
.B(n_68),
.Y(n_272)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_2),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_32),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_53),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_2),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_2),
.B(n_50),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_2),
.B(n_48),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_2),
.B(n_68),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_3),
.B(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_3),
.B(n_68),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_32),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_3),
.B(n_53),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_3),
.B(n_50),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_4),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_4),
.B(n_17),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_4),
.B(n_32),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_4),
.B(n_53),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_53),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_68),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_5),
.B(n_271),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_8),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_50),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_8),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_8),
.B(n_48),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_53),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_13),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_13),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_13),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_13),
.B(n_32),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_13),
.B(n_53),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_14),
.B(n_48),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_14),
.B(n_68),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_14),
.B(n_50),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_14),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_14),
.B(n_32),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_14),
.B(n_27),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_44),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_16),
.B(n_50),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_16),
.B(n_48),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_16),
.B(n_53),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_16),
.B(n_32),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_16),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_16),
.B(n_68),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_16),
.B(n_27),
.Y(n_260)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_17),
.Y(n_174)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_17),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_148),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.C(n_91),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_21),
.B(n_79),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_56),
.C(n_73),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_46),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_23),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_29),
.C(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_62),
.Y(n_125)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_29),
.A2(n_39),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g132 ( 
.A(n_29),
.B(n_81),
.C(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_30),
.B(n_63),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_31),
.B(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_34),
.A2(n_38),
.B1(n_41),
.B2(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_41),
.C(n_42),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_40),
.B(n_46),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_41),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_42),
.A2(n_43),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_44),
.Y(n_276)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_45),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_46),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.CI(n_52),
.CON(n_46),
.SN(n_46)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_49),
.C(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_53),
.Y(n_216)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_73),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_67),
.C(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_57),
.A2(n_58),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_64),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_61),
.CI(n_64),
.CON(n_93),
.SN(n_93)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_71),
.B1(n_77),
.B2(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_67),
.B(n_76),
.C(n_78),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_71),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_86),
.C(n_87),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_84),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_87),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.CI(n_90),
.CON(n_87),
.SN(n_87)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_91),
.B(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_104),
.C(n_108),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_92),
.B(n_104),
.CI(n_108),
.CON(n_325),
.SN(n_325)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.C(n_100),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_93),
.B(n_309),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_93),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_94),
.B(n_100),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_97),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_116),
.C(n_117),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_109),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_109),
.B(n_315),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_112),
.CI(n_115),
.CON(n_109),
.SN(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_116),
.B(n_117),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_133),
.B2(n_134),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_129),
.B2(n_130),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_127),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_327),
.C(n_328),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_318),
.C(n_319),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_304),
.C(n_305),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_282),
.C(n_283),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_250),
.C(n_251),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_225),
.C(n_226),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_186),
.C(n_198),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_169),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_164),
.C(n_169),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_159),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_167),
.C(n_168),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_178),
.C(n_179),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_174),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_185),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_185),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_197),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_191),
.B1(n_197),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_221),
.C(n_222),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.C(n_212),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_205),
.C(n_206),
.Y(n_221)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.C(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_215),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_239),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_240),
.C(n_249),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_235),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_234),
.C(n_235),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_233),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_235),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.CI(n_238),
.CON(n_235),
.SN(n_235)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_249),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_243),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_246),
.C(n_248),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_266),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_255),
.C(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_262),
.C(n_265),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_257),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.CI(n_260),
.CON(n_257),
.SN(n_257)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_274),
.C(n_280),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B1(n_280),
.B2(n_281),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_272),
.B(n_273),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_272),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_301),
.C(n_302),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_274),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_278),
.C(n_279),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_297),
.B2(n_303),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_298),
.C(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_295),
.C(n_296),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_316),
.B2(n_317),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_310),
.C(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_322),
.C(n_326),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_325),
.Y(n_330)
);


endmodule