module fake_jpeg_25953_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_60),
.Y(n_86)
);

BUFx2_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_18),
.Y(n_100)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_31),
.B1(n_17),
.B2(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_82),
.B1(n_93),
.B2(n_50),
.Y(n_112)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_78),
.Y(n_104)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_31),
.B1(n_17),
.B2(n_46),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_87),
.Y(n_123)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_34),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_42),
.B1(n_31),
.B2(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_34),
.B1(n_27),
.B2(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_27),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_22),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_35),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_35),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_118),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_78),
.B1(n_79),
.B2(n_87),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_54),
.B1(n_32),
.B2(n_20),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_117),
.B1(n_129),
.B2(n_85),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_43),
.C(n_45),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_109),
.C(n_118),
.Y(n_146)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_72),
.Y(n_135)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_35),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_54),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_81),
.A2(n_32),
.B1(n_20),
.B2(n_25),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_131),
.A2(n_144),
.B(n_119),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_127),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_96),
.B1(n_91),
.B2(n_76),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_150),
.B1(n_125),
.B2(n_120),
.Y(n_169)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_107),
.B(n_23),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_71),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_9),
.C(n_15),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_145),
.Y(n_175)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_19),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_105),
.B(n_19),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_85),
.B1(n_99),
.B2(n_88),
.Y(n_150)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_156),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_102),
.B(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_26),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_30),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_158),
.Y(n_188)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_173),
.C(n_180),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_84),
.B1(n_106),
.B2(n_108),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_183),
.B1(n_0),
.B2(n_1),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_121),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_170),
.B1(n_186),
.B2(n_131),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_119),
.B1(n_106),
.B2(n_125),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_124),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_191),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_174),
.B(n_155),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_120),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_20),
.B(n_32),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_103),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_1),
.B(n_5),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_30),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_130),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_73),
.C(n_108),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_187),
.C(n_156),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_107),
.B1(n_25),
.B2(n_23),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_133),
.Y(n_187)
);

NAND2x1p5_ASAP7_75t_L g189 ( 
.A(n_131),
.B(n_44),
.Y(n_189)
);

NAND2x1p5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_28),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_205),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_194),
.A2(n_195),
.B(n_214),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_134),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_198),
.B(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_202),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_201),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

CKINVDCx12_ASAP7_75t_R g205 ( 
.A(n_164),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_216),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_143),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_152),
.B1(n_28),
.B2(n_4),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_217),
.B1(n_189),
.B2(n_174),
.Y(n_223)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_28),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_219),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_184),
.B1(n_179),
.B2(n_172),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_9),
.C(n_4),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_163),
.B1(n_171),
.B2(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_5),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_161),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_191),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_232),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_235),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_6),
.C(n_7),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_179),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_211),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_248),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_207),
.C(n_203),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_262),
.C(n_228),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_202),
.B1(n_196),
.B2(n_215),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_256),
.A2(n_263),
.B1(n_268),
.B2(n_239),
.Y(n_283)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_198),
.B(n_220),
.C(n_203),
.D(n_210),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_243),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_204),
.C(n_194),
.Y(n_262)
);

NAND2xp67_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_212),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_264),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_232),
.A2(n_200),
.B1(n_192),
.B2(n_9),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_239),
.B1(n_237),
.B2(n_246),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_6),
.B(n_8),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_10),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_262),
.C(n_261),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_226),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_287),
.Y(n_291)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_285),
.Y(n_303)
);

HAxp5_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_252),
.CON(n_299),
.SN(n_299)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_267),
.B1(n_260),
.B2(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_235),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_286),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_226),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_228),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_292),
.B(n_296),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_252),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_272),
.Y(n_304)
);

BUFx12_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_275),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_266),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_253),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_281),
.Y(n_308)
);

BUFx12_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_302),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_251),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_303),
.B1(n_289),
.B2(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_307),
.A2(n_247),
.B1(n_302),
.B2(n_240),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_314),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_272),
.C(n_271),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_313),
.C(n_296),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_274),
.B(n_231),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_274),
.B(n_231),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_245),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_258),
.C(n_225),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_268),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_259),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_317),
.B(n_304),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_320),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_305),
.A2(n_302),
.B1(n_257),
.B2(n_241),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_313),
.C(n_309),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_225),
.B1(n_234),
.B2(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_312),
.Y(n_327)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_234),
.B(n_12),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_319),
.B(n_326),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_334),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_335),
.B(n_331),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_321),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_332),
.B1(n_318),
.B2(n_322),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_11),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_320),
.C2(n_325),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_11),
.B(n_12),
.Y(n_342)
);


endmodule