module fake_jpeg_14368_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_60),
.B(n_65),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_24),
.Y(n_61)
);

CKINVDCx6p67_ASAP7_75t_R g154 ( 
.A(n_61),
.Y(n_154)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_16),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_20),
.B(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_88),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_24),
.Y(n_82)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_84),
.B(n_92),
.Y(n_135)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx4f_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_94),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_91),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_24),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_15),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_97),
.Y(n_116)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_99),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_102),
.Y(n_140)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_25),
.Y(n_141)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_49),
.B1(n_29),
.B2(n_46),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_105),
.A2(n_134),
.B1(n_144),
.B2(n_54),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_22),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_115),
.B(n_137),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_61),
.A2(n_41),
.B1(n_52),
.B2(n_38),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_129),
.B1(n_151),
.B2(n_56),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_43),
.B1(n_38),
.B2(n_30),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_82),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_20),
.B1(n_28),
.B2(n_31),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_126),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_59),
.B(n_36),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_143),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_41),
.B1(n_52),
.B2(n_38),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_43),
.B1(n_52),
.B2(n_41),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_69),
.B(n_50),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_57),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_63),
.B(n_35),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_66),
.B(n_35),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_66),
.B(n_36),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_67),
.B(n_31),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_155),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_86),
.A2(n_25),
.B1(n_30),
.B2(n_50),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_44),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_70),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_157),
.B(n_4),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_77),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_163),
.B(n_164),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_14),
.B(n_44),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_165),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_83),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_169),
.B(n_179),
.Y(n_258)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_42),
.B1(n_47),
.B2(n_37),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_70),
.C(n_103),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_174),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_108),
.A2(n_104),
.B(n_96),
.C(n_74),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_175),
.A2(n_219),
.B(n_160),
.C(n_154),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_122),
.B(n_55),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_113),
.B(n_37),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_99),
.B1(n_97),
.B2(n_92),
.Y(n_180)
);

AO22x1_ASAP7_75t_SL g260 ( 
.A1(n_180),
.A2(n_211),
.B1(n_154),
.B2(n_160),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_181),
.B(n_191),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_105),
.A2(n_91),
.B1(n_90),
.B2(n_81),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_136),
.B1(n_112),
.B2(n_123),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_75),
.B1(n_72),
.B2(n_64),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_183),
.A2(n_188),
.B1(n_200),
.B2(n_209),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_185),
.A2(n_152),
.B1(n_161),
.B2(n_154),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_195),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_187),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_135),
.A2(n_58),
.B1(n_30),
.B2(n_28),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_189),
.Y(n_265)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_47),
.C(n_42),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_111),
.B(n_30),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_148),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_193),
.B(n_194),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_14),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_127),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_201),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_203),
.Y(n_270)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_146),
.A2(n_30),
.B1(n_14),
.B2(n_2),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_109),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_210),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_109),
.B(n_0),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_149),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_159),
.B1(n_125),
.B2(n_138),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_1),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_107),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_213),
.Y(n_251)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_217),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_117),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_215),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_156),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_144),
.B1(n_107),
.B2(n_130),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_109),
.B(n_6),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_120),
.A2(n_6),
.B(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_158),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_222),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_185),
.A2(n_136),
.B1(n_112),
.B2(n_145),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_227),
.B1(n_238),
.B2(n_268),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g272 ( 
.A(n_231),
.B(n_249),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_130),
.B1(n_123),
.B2(n_145),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_166),
.B(n_144),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_247),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_245),
.B1(n_260),
.B2(n_266),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_188),
.A2(n_142),
.B1(n_121),
.B2(n_139),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_166),
.B(n_139),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_217),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_261),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_176),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_173),
.B(n_131),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_264),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_176),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_176),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_218),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_131),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_209),
.A2(n_125),
.B1(n_152),
.B2(n_118),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_200),
.A2(n_161),
.B1(n_133),
.B2(n_110),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_267),
.A2(n_164),
.B1(n_186),
.B2(n_215),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_178),
.A2(n_133),
.B1(n_10),
.B2(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_273),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_192),
.C(n_181),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_290),
.C(n_298),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_230),
.A2(n_177),
.B1(n_184),
.B2(n_180),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_275),
.A2(n_284),
.B1(n_303),
.B2(n_313),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_229),
.B(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_276),
.B(n_277),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_229),
.B(n_167),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_248),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_231),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_242),
.B(n_167),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_283),
.B(n_289),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_230),
.A2(n_177),
.B1(n_184),
.B2(n_180),
.Y(n_284)
);

BUFx8_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_288),
.B(n_292),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_252),
.B(n_179),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_198),
.C(n_201),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_291),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_248),
.B(n_191),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_247),
.B(n_174),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_295),
.B(n_300),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_222),
.A2(n_175),
.B1(n_216),
.B2(n_198),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_296),
.A2(n_245),
.B1(n_267),
.B2(n_266),
.Y(n_345)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_219),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_305),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_224),
.B(n_172),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_243),
.B(n_197),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_301),
.B(n_226),
.Y(n_330)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_211),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_226),
.B(n_211),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_205),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_309),
.A2(n_312),
.B(n_318),
.Y(n_358)
);

INVx4_ASAP7_75t_SL g310 ( 
.A(n_246),
.Y(n_310)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_233),
.B(n_220),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_250),
.A2(n_215),
.B(n_211),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_244),
.A2(n_214),
.B1(n_199),
.B2(n_204),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_196),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_316),
.Y(n_333)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_225),
.B(n_170),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_225),
.B(n_208),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_270),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_250),
.A2(n_213),
.B(n_190),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_272),
.A2(n_254),
.B(n_239),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_322),
.A2(n_324),
.B(n_318),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_254),
.B(n_239),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_309),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_306),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_225),
.C(n_270),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_356),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_330),
.B(n_342),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_302),
.A2(n_256),
.B1(n_223),
.B2(n_249),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_344),
.B1(n_312),
.B2(n_324),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_279),
.B(n_263),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_348),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_275),
.A2(n_222),
.B1(n_256),
.B2(n_227),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_345),
.A2(n_359),
.B1(n_287),
.B2(n_284),
.Y(n_363)
);

XOR2x1_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_316),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_222),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_279),
.B(n_222),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_353),
.Y(n_366)
);

CKINVDCx10_ASAP7_75t_R g350 ( 
.A(n_310),
.Y(n_350)
);

INVx3_ASAP7_75t_SL g378 ( 
.A(n_350),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_286),
.B(n_240),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_260),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_357),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_280),
.B(n_262),
.C(n_251),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_241),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_296),
.A2(n_260),
.B1(n_253),
.B2(n_238),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_280),
.B(n_268),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_281),
.Y(n_373)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_363),
.A2(n_368),
.B1(n_371),
.B2(n_339),
.Y(n_413)
);

XOR2x1_ASAP7_75t_L g421 ( 
.A(n_365),
.B(n_390),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_367),
.A2(n_376),
.B1(n_355),
.B2(n_360),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_288),
.B1(n_308),
.B2(n_305),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_350),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_369),
.B(n_372),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_345),
.A2(n_288),
.B1(n_299),
.B2(n_313),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_353),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_374),
.Y(n_398)
);

OAI32xp33_ASAP7_75t_L g374 ( 
.A1(n_323),
.A2(n_317),
.A3(n_273),
.B1(n_307),
.B2(n_297),
.Y(n_374)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_339),
.A2(n_281),
.B1(n_274),
.B2(n_290),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_326),
.B(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_381),
.B(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_357),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_384),
.A2(n_385),
.B(n_386),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_358),
.A2(n_294),
.B(n_255),
.Y(n_385)
);

A2O1A1O1Ixp25_ASAP7_75t_L g386 ( 
.A1(n_323),
.A2(n_293),
.B(n_310),
.C(n_315),
.D(n_285),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_285),
.Y(n_387)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_392),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_329),
.B(n_285),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_319),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_355),
.A2(n_322),
.B1(n_342),
.B2(n_327),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_291),
.B(n_241),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_391),
.Y(n_404)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_395),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_236),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_356),
.C(n_346),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_320),
.B(n_304),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_348),
.A2(n_253),
.B(n_236),
.Y(n_396)
);

OAI21xp33_ASAP7_75t_SL g416 ( 
.A1(n_396),
.A2(n_333),
.B(n_344),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_397),
.B(n_402),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_419),
.C(n_423),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_387),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_409),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_341),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_397),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_395),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_413),
.A2(n_416),
.B1(n_424),
.B2(n_366),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_414),
.A2(n_390),
.B1(n_384),
.B2(n_330),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_354),
.Y(n_415)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_321),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_325),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_355),
.C(n_320),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_341),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_420),
.A2(n_385),
.B1(n_396),
.B2(n_391),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_333),
.C(n_349),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_363),
.A2(n_371),
.B1(n_368),
.B2(n_373),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_362),
.B(n_347),
.Y(n_425)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_425),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_370),
.B(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_426),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_370),
.B(n_374),
.Y(n_427)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_376),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_435),
.C(n_437),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_430),
.A2(n_432),
.B1(n_439),
.B2(n_427),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_412),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_414),
.A2(n_366),
.B1(n_365),
.B2(n_340),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_433),
.A2(n_434),
.B1(n_436),
.B2(n_447),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_413),
.A2(n_393),
.B1(n_392),
.B2(n_361),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_388),
.B1(n_382),
.B2(n_377),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_389),
.C(n_328),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_443),
.C(n_444),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_398),
.A2(n_340),
.B1(n_328),
.B2(n_378),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_352),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_352),
.C(n_378),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_378),
.C(n_338),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_449),
.C(n_451),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_407),
.A2(n_404),
.B1(n_422),
.B2(n_398),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_332),
.C(n_351),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_401),
.Y(n_450)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_332),
.C(n_351),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_452),
.B(n_453),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_235),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_455),
.A2(n_462),
.B1(n_472),
.B2(n_334),
.Y(n_484)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_440),
.Y(n_456)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_456),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_434),
.Y(n_457)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_408),
.B(n_403),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_458),
.A2(n_438),
.B(n_428),
.Y(n_480)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_446),
.Y(n_460)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_444),
.A2(n_409),
.B1(n_420),
.B2(n_408),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_415),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_466),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_433),
.A2(n_426),
.B1(n_425),
.B2(n_410),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_465),
.B1(n_334),
.B2(n_435),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_L g465 ( 
.A1(n_448),
.A2(n_410),
.B(n_400),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_417),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_436),
.B(n_417),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_471),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_439),
.B(n_400),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_429),
.B(n_412),
.C(n_411),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_473),
.B(n_437),
.Y(n_481)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_432),
.B(n_351),
.CI(n_399),
.CON(n_474),
.SN(n_474)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_445),
.Y(n_479)
);

AO221x1_ASAP7_75t_L g477 ( 
.A1(n_461),
.A2(n_399),
.B1(n_411),
.B2(n_449),
.C(n_334),
.Y(n_477)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_477),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_429),
.C(n_443),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_478),
.B(n_481),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_479),
.A2(n_480),
.B(n_470),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_467),
.B1(n_463),
.B2(n_474),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_454),
.B1(n_464),
.B2(n_457),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_468),
.B(n_235),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_486),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_469),
.B(n_237),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_253),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_489),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_237),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_491),
.Y(n_506)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_460),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_478),
.B(n_469),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_494),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_497),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_470),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_483),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_462),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_458),
.B(n_455),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_499),
.A2(n_189),
.B(n_234),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_457),
.Y(n_500)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_500),
.Y(n_511)
);

AOI21x1_ASAP7_75t_L g502 ( 
.A1(n_475),
.A2(n_471),
.B(n_466),
.Y(n_502)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_502),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_503),
.A2(n_488),
.B1(n_475),
.B2(n_483),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_476),
.B(n_459),
.C(n_474),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_212),
.C(n_10),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_513),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_508),
.A2(n_510),
.B1(n_504),
.B2(n_500),
.Y(n_522)
);

AOI322xp5_ASAP7_75t_L g509 ( 
.A1(n_505),
.A2(n_491),
.A3(n_487),
.B1(n_489),
.B2(n_459),
.C1(n_265),
.C2(n_234),
.Y(n_509)
);

AOI31xp67_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_506),
.A3(n_501),
.B(n_495),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_496),
.A2(n_487),
.B1(n_189),
.B2(n_265),
.Y(n_510)
);

OAI211xp5_ASAP7_75t_L g523 ( 
.A1(n_512),
.A2(n_499),
.B(n_497),
.C(n_494),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_517)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_517),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_498),
.C(n_493),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_521),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_522),
.B(n_523),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_11),
.Y(n_524)
);

A2O1A1O1Ixp25_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_516),
.B(n_511),
.C(n_517),
.D(n_507),
.Y(n_528)
);

FAx1_ASAP7_75t_SL g526 ( 
.A(n_520),
.B(n_513),
.CI(n_514),
.CON(n_526),
.SN(n_526)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_528),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_527),
.C(n_508),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_527),
.B1(n_523),
.B2(n_512),
.Y(n_531)
);

AO21x1_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_532),
.B(n_13),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_529),
.A2(n_518),
.B(n_12),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_13),
.Y(n_534)
);


endmodule