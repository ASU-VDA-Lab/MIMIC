module fake_jpeg_14232_n_443 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_443);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_443;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_47),
.B(n_48),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_51),
.B(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx2_ASAP7_75t_SL g133 ( 
.A(n_56),
.Y(n_133)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_62),
.Y(n_95)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_15),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_15),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_68),
.B(n_82),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_83),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_88),
.Y(n_112)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_0),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_19),
.B(n_1),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_24),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_34),
.Y(n_94)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_91),
.Y(n_142)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_94),
.B(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_31),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_27),
.B1(n_25),
.B2(n_39),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_116),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_27),
.B1(n_25),
.B2(n_43),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_117),
.B1(n_122),
.B2(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_34),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_73),
.B1(n_86),
.B2(n_78),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_49),
.A2(n_27),
.B1(n_25),
.B2(n_43),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_77),
.A2(n_25),
.B1(n_43),
.B2(n_39),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_28),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_64),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_30),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_39),
.B1(n_43),
.B2(n_41),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_143),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_69),
.A2(n_42),
.B1(n_29),
.B2(n_41),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_144),
.B1(n_145),
.B2(n_7),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_71),
.A2(n_41),
.B1(n_32),
.B2(n_40),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_64),
.A2(n_41),
.B1(n_32),
.B2(n_40),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_42),
.B1(n_29),
.B2(n_40),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_106),
.B(n_56),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_155),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_32),
.B1(n_26),
.B2(n_30),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_147),
.A2(n_161),
.B1(n_131),
.B2(n_134),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_151),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_30),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_95),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_163),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_101),
.Y(n_158)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_1),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_159),
.B(n_171),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_84),
.C(n_70),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_174),
.C(n_182),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_92),
.A2(n_26),
.B1(n_44),
.B2(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_97),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_2),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_164),
.Y(n_218)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx6_ASAP7_75t_SL g167 ( 
.A(n_99),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_124),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_169),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_44),
.C(n_3),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_44),
.B1(n_4),
.B2(n_5),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_175),
.A2(n_184),
.B1(n_187),
.B2(n_113),
.Y(n_236)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_2),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_180),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_120),
.B(n_5),
.C(n_6),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_140),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_96),
.B(n_5),
.Y(n_182)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_112),
.A2(n_44),
.B1(n_8),
.B2(n_9),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_118),
.B(n_7),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_186),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_7),
.Y(n_186)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_111),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_123),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_96),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_104),
.B(n_10),
.Y(n_193)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_100),
.B(n_10),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_195),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_105),
.B(n_10),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_197),
.C(n_136),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_11),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_105),
.C(n_109),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_201),
.B(n_233),
.CI(n_160),
.CON(n_253),
.SN(n_253)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_154),
.B(n_109),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_205),
.B(n_189),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_162),
.A2(n_132),
.B1(n_113),
.B2(n_121),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_241),
.B1(n_187),
.B2(n_158),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_150),
.A2(n_132),
.B1(n_121),
.B2(n_131),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_194),
.B1(n_170),
.B2(n_178),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_216),
.B(n_11),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_150),
.A2(n_111),
.B(n_136),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_221),
.A2(n_231),
.B(n_110),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_166),
.A2(n_100),
.B(n_137),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_167),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_158),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_148),
.B(n_134),
.C(n_141),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_236),
.A2(n_239),
.B1(n_170),
.B2(n_188),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_166),
.A2(n_123),
.B1(n_141),
.B2(n_137),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_154),
.A2(n_110),
.B1(n_12),
.B2(n_13),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_164),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_244),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_243),
.B(n_245),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_164),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_157),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_155),
.B(n_197),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_249),
.B(n_275),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g247 ( 
.A1(n_202),
.A2(n_197),
.B(n_146),
.Y(n_247)
);

AO32x1_ASAP7_75t_L g291 ( 
.A1(n_247),
.A2(n_218),
.A3(n_241),
.B1(n_203),
.B2(n_237),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_248),
.A2(n_255),
.B1(n_259),
.B2(n_265),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_221),
.A2(n_184),
.B(n_175),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_257),
.B1(n_262),
.B2(n_266),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_253),
.B(n_276),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_149),
.B1(n_182),
.B2(n_174),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_211),
.A2(n_149),
.B1(n_172),
.B2(n_152),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_SL g301 ( 
.A1(n_256),
.A2(n_237),
.B(n_224),
.C(n_238),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_211),
.A2(n_159),
.B1(n_190),
.B2(n_173),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_198),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_258),
.B(n_261),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_235),
.A2(n_171),
.B1(n_191),
.B2(n_176),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_168),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_206),
.B(n_163),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_205),
.A2(n_183),
.B1(n_152),
.B2(n_178),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_209),
.A2(n_203),
.B1(n_226),
.B2(n_240),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_205),
.B(n_207),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_204),
.Y(n_269)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_207),
.A2(n_153),
.B1(n_165),
.B2(n_192),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_199),
.Y(n_272)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_202),
.A2(n_189),
.B1(n_110),
.B2(n_14),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_200),
.B1(n_227),
.B2(n_220),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_275),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_226),
.A2(n_13),
.B1(n_14),
.B2(n_206),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_200),
.B1(n_232),
.B2(n_222),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_13),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_227),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_234),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_225),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_210),
.B(n_233),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_309),
.B1(n_262),
.B2(n_267),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_230),
.B(n_234),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_284),
.A2(n_299),
.B(n_283),
.Y(n_325)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_287),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_201),
.C(n_216),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_300),
.C(n_307),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_276),
.C(n_261),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_295),
.A2(n_314),
.B1(n_278),
.B2(n_248),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_298),
.B(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_218),
.C(n_220),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_301),
.A2(n_274),
.B1(n_256),
.B2(n_271),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_311),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_228),
.C(n_214),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_238),
.C(n_225),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_310),
.C(n_300),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_254),
.A2(n_222),
.B1(n_215),
.B2(n_223),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_214),
.C(n_215),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_260),
.A3(n_250),
.B1(n_259),
.B2(n_244),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_263),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_267),
.A2(n_252),
.B1(n_257),
.B2(n_255),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_315),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_296),
.B(n_245),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_324),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_318),
.A2(n_329),
.B1(n_332),
.B2(n_334),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_319),
.A2(n_327),
.B(n_339),
.Y(n_354)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_326),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_253),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_330),
.C(n_336),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_292),
.B(n_258),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_328),
.B(n_302),
.Y(n_344)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_253),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_292),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_331),
.Y(n_355)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_243),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

AO32x1_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_246),
.A3(n_256),
.B1(n_274),
.B2(n_249),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_340),
.B1(n_342),
.B2(n_312),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_242),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_338),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_290),
.B(n_251),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_339),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_312),
.A2(n_273),
.B1(n_264),
.B2(n_270),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_269),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_298),
.C(n_301),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_344),
.A2(n_355),
.B(n_366),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_310),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_347),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_346),
.A2(n_359),
.B1(n_360),
.B2(n_320),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_293),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_293),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_358),
.C(n_364),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_322),
.A2(n_314),
.B1(n_282),
.B2(n_302),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_352),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_322),
.A2(n_302),
.B1(n_305),
.B2(n_284),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_333),
.A2(n_335),
.B1(n_328),
.B2(n_331),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_354),
.B(n_237),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_311),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_319),
.A2(n_308),
.B1(n_301),
.B2(n_307),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_301),
.B1(n_287),
.B2(n_289),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_337),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_278),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_342),
.A2(n_289),
.B1(n_272),
.B2(n_222),
.Y(n_365)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_365),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_368),
.B(n_371),
.Y(n_396)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_321),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_334),
.C(n_332),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_377),
.C(n_347),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_359),
.A2(n_315),
.B1(n_329),
.B2(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_381),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_376),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_348),
.B(n_237),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_337),
.C(n_223),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_378),
.A2(n_360),
.B(n_355),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_383),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_344),
.A2(n_229),
.B(n_199),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_SL g383 ( 
.A(n_352),
.B(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_384),
.Y(n_394)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_385),
.B(n_361),
.Y(n_398)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_364),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_373),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_398),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_363),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_392),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_349),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_401),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_379),
.A2(n_361),
.B1(n_362),
.B2(n_345),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_399),
.B(n_402),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_400),
.B(n_377),
.C(n_382),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_356),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_397),
.A2(n_374),
.B(n_367),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_395),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_407),
.C(n_412),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_370),
.C(n_382),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_396),
.B(n_370),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_408),
.B(n_413),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_401),
.A2(n_367),
.B(n_350),
.Y(n_411)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_411),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_392),
.C(n_391),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_399),
.Y(n_413)
);

AOI22x1_ASAP7_75t_L g427 ( 
.A1(n_415),
.A2(n_418),
.B1(n_423),
.B2(n_388),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_405),
.A2(n_394),
.B1(n_402),
.B2(n_390),
.Y(n_416)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_416),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_383),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_420),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_409),
.A2(n_375),
.B1(n_369),
.B2(n_390),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_414),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_356),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_419),
.A2(n_404),
.B(n_406),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_426),
.B(n_427),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_422),
.A2(n_407),
.B(n_403),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_429),
.B(n_417),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_415),
.A2(n_410),
.B(n_388),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_421),
.B(n_381),
.Y(n_434)
);

AND2x2_ASAP7_75t_SL g436 ( 
.A(n_431),
.B(n_410),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_428),
.A2(n_423),
.B(n_416),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_432),
.A2(n_434),
.B(n_424),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_435),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_436),
.B(n_437),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_389),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_438),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_440),
.A2(n_439),
.B(n_389),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_376),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_442),
.B(n_229),
.Y(n_443)
);


endmodule