module fake_jpeg_26520_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_51),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_0),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_48),
.B1(n_41),
.B2(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_69),
.B1(n_44),
.B2(n_73),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_53),
.B1(n_47),
.B2(n_52),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_52),
.B1(n_43),
.B2(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_1),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_1),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_89),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_43),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_86),
.B1(n_90),
.B2(n_3),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_85),
.Y(n_94)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_92),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_73),
.B1(n_21),
.B2(n_22),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_3),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_19),
.B1(n_38),
.B2(n_35),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_97),
.B1(n_81),
.B2(n_84),
.Y(n_110)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_80),
.CON(n_105),
.SN(n_105)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_15),
.B1(n_34),
.B2(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_7),
.Y(n_108)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_101),
.B1(n_81),
.B2(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_110),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_7),
.C(n_8),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_93),
.B1(n_97),
.B2(n_96),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_109),
.B1(n_107),
.B2(n_96),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_111),
.C(n_9),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_122),
.C(n_10),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_23),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_24),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_20),
.C(n_11),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_27),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_28),
.B1(n_12),
.B2(n_14),
.Y(n_131)
);


endmodule