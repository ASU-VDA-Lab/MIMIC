module fake_netlist_1_367_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
NOR2xp33_ASAP7_75t_L g10 ( .A(n_5), .B(n_4), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_9), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
BUFx8_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
NOR2x1p5_ASAP7_75t_L g18 ( .A(n_12), .B(n_1), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_10), .B(n_1), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_13), .B(n_2), .Y(n_22) );
OAI21x1_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_11), .B(n_16), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_17), .B1(n_15), .B2(n_14), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
OAI221xp5_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_16), .B1(n_4), .B2(n_5), .C(n_6), .Y(n_26) );
INVx4_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AOI31xp33_ASAP7_75t_L g29 ( .A1(n_24), .A2(n_21), .A3(n_20), .B(n_18), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_26), .B1(n_21), .B2(n_28), .C(n_27), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_27), .B1(n_28), .B2(n_23), .Y(n_36) );
AOI221xp5_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_27), .B1(n_23), .B2(n_6), .C(n_2), .Y(n_37) );
HB1xp67_ASAP7_75t_L g38 ( .A(n_34), .Y(n_38) );
XNOR2x1_ASAP7_75t_L g39 ( .A(n_38), .B(n_35), .Y(n_39) );
AOI22xp33_ASAP7_75t_SL g40 ( .A1(n_39), .A2(n_36), .B1(n_16), .B2(n_37), .Y(n_40) );
endmodule