module fake_jpeg_24083_n_131 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_14),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_21),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_46),
.B(n_48),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_27),
.C(n_19),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_55),
.C(n_7),
.Y(n_77)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.C(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_29),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_20),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_30),
.A2(n_23),
.B1(n_14),
.B2(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_24),
.B1(n_22),
.B2(n_17),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_76),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_24),
.B(n_17),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_78),
.B(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_70),
.A3(n_42),
.B1(n_53),
.B2(n_54),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_50),
.B(n_45),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_72),
.C(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_16),
.B1(n_25),
.B2(n_2),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_1),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_7),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_47),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_9),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_10),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_95),
.B1(n_71),
.B2(n_70),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_49),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_94),
.B(n_75),
.Y(n_101)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_63),
.B1(n_89),
.B2(n_64),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_69),
.C(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_102),
.C(n_105),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_105),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_69),
.C(n_74),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_74),
.C(n_71),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_76),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_110),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_102),
.C(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_95),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_99),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_120),
.C(n_109),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_96),
.B1(n_114),
.B2(n_101),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_122),
.B1(n_78),
.B2(n_123),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_107),
.B1(n_79),
.B2(n_91),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_124),
.B(n_52),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_107),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_79),
.B(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_127),
.B1(n_78),
.B2(n_43),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_118),
.C(n_51),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.C(n_111),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);


endmodule