module real_jpeg_33455_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g415 ( 
.A(n_0),
.Y(n_415)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_2),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_2),
.A2(n_81),
.B1(n_277),
.B2(n_281),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_2),
.A2(n_81),
.B1(n_567),
.B2(n_569),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_3),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_3),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_3),
.A2(n_168),
.B1(n_261),
.B2(n_264),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_3),
.A2(n_168),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_3),
.A2(n_168),
.B1(n_467),
.B2(n_471),
.Y(n_466)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_4),
.A2(n_291),
.B1(n_294),
.B2(n_297),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_4),
.Y(n_297)
);

AO22x1_ASAP7_75t_L g559 ( 
.A1(n_4),
.A2(n_297),
.B1(n_560),
.B2(n_563),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_196),
.B1(n_201),
.B2(n_202),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_5),
.A2(n_201),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_5),
.A2(n_201),
.B1(n_319),
.B2(n_323),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_5),
.A2(n_577),
.B(n_579),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_5),
.B(n_580),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_6),
.A2(n_146),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_6),
.A2(n_151),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_6),
.A2(n_65),
.B1(n_151),
.B2(n_382),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_6),
.A2(n_151),
.B1(n_535),
.B2(n_538),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_8),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_9),
.Y(n_377)
);

AOI22x1_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_118),
.B1(n_121),
.B2(n_126),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_10),
.A2(n_126),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_10),
.A2(n_126),
.B1(n_207),
.B2(n_388),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_10),
.A2(n_126),
.B1(n_403),
.B2(n_405),
.Y(n_402)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_11),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_12),
.A2(n_33),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_12),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_12),
.A2(n_93),
.B1(n_306),
.B2(n_309),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_12),
.A2(n_93),
.B1(n_349),
.B2(n_352),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_12),
.A2(n_93),
.B1(n_397),
.B2(n_401),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_13),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_13),
.A2(n_70),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_13),
.A2(n_70),
.B1(n_456),
.B2(n_460),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_14),
.A2(n_213),
.B1(n_215),
.B2(n_218),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_14),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_14),
.A2(n_207),
.B1(n_218),
.B2(n_520),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_16),
.A2(n_58),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_16),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_16),
.B(n_131),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_16),
.A2(n_72),
.B1(n_396),
.B2(n_414),
.Y(n_413)
);

OAI32xp33_ASAP7_75t_L g433 ( 
.A1(n_16),
.A2(n_155),
.A3(n_434),
.B1(n_438),
.B2(n_442),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_16),
.A2(n_327),
.B1(n_455),
.B2(n_459),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_17),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_17),
.Y(n_144)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_17),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_18),
.Y(n_464)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_546),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_505),
.B(n_543),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_332),
.B(n_502),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_298),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_248),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_29),
.B(n_248),
.C(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_172),
.C(n_223),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_30),
.B(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_88),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_31),
.B(n_251),
.C(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_62),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_32),
.A2(n_62),
.B1(n_63),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_32),
.Y(n_329)
);

OAI32xp33_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_37),
.A3(n_40),
.B1(n_46),
.B2(n_57),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g265 ( 
.A(n_35),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_36),
.Y(n_537)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_38),
.Y(n_156)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_39),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_52),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_56),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_56),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_56),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_56),
.Y(n_313)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_71),
.B1(n_78),
.B2(n_86),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_64),
.A2(n_71),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_66),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_68),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_71),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_71),
.A2(n_318),
.B1(n_381),
.B2(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_72),
.A2(n_79),
.B1(n_212),
.B2(n_219),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_72),
.A2(n_212),
.B(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_72),
.A2(n_396),
.B1(n_402),
.B2(n_409),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_72),
.B(n_527),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_75),
.Y(n_222)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_75),
.Y(n_317)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_77),
.Y(n_214)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_77),
.Y(n_372)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_85),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_129),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_90),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_98),
.B1(n_116),
.B2(n_127),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_92),
.A2(n_128),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_94),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_100),
.B1(n_103),
.B2(n_105),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_96),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_98),
.Y(n_236)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_98),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_98),
.A2(n_532),
.B1(n_533),
.B2(n_534),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_98),
.A2(n_127),
.B1(n_534),
.B2(n_576),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_107)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_109),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_110),
.Y(n_308)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_117),
.A2(n_128),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_124),
.Y(n_538)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2x1_ASAP7_75t_R g326 ( 
.A(n_128),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_128),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_129),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_145),
.B1(n_154),
.B2(n_163),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_130),
.A2(n_154),
.B1(n_163),
.B2(n_227),
.Y(n_226)
);

OAI22x1_ASAP7_75t_L g267 ( 
.A1(n_130),
.A2(n_145),
.B1(n_154),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_130),
.A2(n_154),
.B1(n_227),
.B2(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_130),
.A2(n_154),
.B1(n_305),
.B2(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22x1_ASAP7_75t_L g539 ( 
.A1(n_131),
.A2(n_540),
.B1(n_541),
.B2(n_542),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_131),
.A2(n_540),
.B1(n_542),
.B2(n_566),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_155),
.B(n_159),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_135),
.B1(n_138),
.B2(n_142),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_135),
.Y(n_352)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_136),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_137),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_137),
.Y(n_389)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_137),
.Y(n_441)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_137),
.Y(n_523)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_144),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_144),
.Y(n_562)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_149),
.Y(n_269)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_150),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_154),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_167),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_173),
.B(n_224),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_211),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_174),
.B(n_211),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_195),
.B1(n_205),
.B2(n_206),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_175),
.A2(n_195),
.B1(n_205),
.B2(n_241),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_175),
.A2(n_205),
.B1(n_206),
.B2(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_175),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_175),
.A2(n_205),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_175),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_175),
.A2(n_205),
.B1(n_276),
.B2(n_519),
.Y(n_518)
);

AO21x2_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_182),
.B(n_189),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_182),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_183),
.Y(n_280)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g470 ( 
.A(n_185),
.Y(n_470)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_189)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_190),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_190),
.Y(n_382)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_191),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_191),
.Y(n_322)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_191),
.Y(n_408)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_200),
.Y(n_283)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_205),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_205),
.B(n_327),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_217),
.Y(n_404)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_220),
.A2(n_422),
.B1(n_423),
.B2(n_424),
.Y(n_421)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.C(n_239),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_240),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_233),
.Y(n_570)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_235),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_241),
.Y(n_490)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_244),
.Y(n_445)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_244),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_250),
.B(n_274),
.C(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_274),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_255),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_256),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_266),
.B1(n_267),
.B2(n_273),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_260),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_263),
.Y(n_578)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_266),
.Y(n_514)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_268),
.Y(n_541)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_273),
.Y(n_513)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_275),
.B(n_284),
.Y(n_529)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_281),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

INVx3_ASAP7_75t_SL g527 ( 
.A(n_286),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_289),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_289),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_289),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_290),
.B(n_526),
.Y(n_525)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_330),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_300),
.B(n_330),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_303),
.C(n_328),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_301),
.B(n_499),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_303),
.B(n_328),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_314),
.C(n_326),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_304),
.B(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_314),
.A2(n_315),
.B1(n_326),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_326),
.Y(n_484)
);

OAI21xp33_ASAP7_75t_SL g341 ( 
.A1(n_327),
.A2(n_342),
.B(n_344),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_327),
.B(n_409),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_327),
.B(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_497),
.B(n_501),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_480),
.B(n_496),
.Y(n_334)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_429),
.B(n_479),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_392),
.B(n_428),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_368),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_338),
.B(n_368),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_354),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_339),
.A2(n_340),
.B1(n_354),
.B2(n_355),
.Y(n_420)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_347),
.B1(n_348),
.B2(n_353),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_347),
.A2(n_353),
.B1(n_466),
.B2(n_476),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_347),
.A2(n_353),
.B1(n_559),
.B2(n_564),
.Y(n_558)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_353),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_363),
.B1(n_364),
.B2(n_367),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_383),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_385),
.C(n_390),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_378),
.B2(n_380),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_390),
.B2(n_391),
.Y(n_383)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_384),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_385),
.Y(n_391)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

OAI31xp33_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_419),
.A3(n_425),
.B(n_427),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_412),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_411),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_395),
.B(n_411),
.Y(n_426)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_401),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

INVx8_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_421),
.Y(n_427)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_SL g479 ( 
.A(n_430),
.B(n_431),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_452),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_432),
.B(n_465),
.C(n_478),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_446),
.B1(n_450),
.B2(n_451),
.Y(n_432)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_433),
.B(n_451),
.Y(n_486)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_446),
.Y(n_451)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_465),
.B1(n_477),
.B2(n_478),
.Y(n_452)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_453),
.Y(n_478)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_495),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_495),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_485),
.B1(n_493),
.B2(n_494),
.Y(n_481)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_482),
.Y(n_494)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_485),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_487),
.B1(n_491),
.B2(n_492),
.Y(n_485)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_486),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_487),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_491),
.C(n_494),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_500),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_500),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_508),
.B(n_510),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_515),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_511),
.B(n_549),
.C(n_550),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.C(n_514),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_528),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

XNOR2x2_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_524),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_518),
.B(n_525),
.Y(n_573)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_519),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_521),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_525),
.B(n_575),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_528),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_529),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_539),
.Y(n_530)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_531),
.Y(n_554)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVxp33_ASAP7_75t_SL g555 ( 
.A(n_539),
.Y(n_555)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_583),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_551),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_548),
.B(n_551),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_556),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_554),
.C(n_555),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_557),
.A2(n_572),
.B1(n_581),
.B2(n_582),
.Y(n_556)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_557),
.Y(n_581)
);

OAI21xp33_ASAP7_75t_L g557 ( 
.A1(n_558),
.A2(n_565),
.B(n_571),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_565),
.Y(n_571)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_572),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_574),
.Y(n_572)
);

INVx8_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVxp33_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);


endmodule