module fake_aes_9858_n_629 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_629);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_629;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g74 ( .A(n_13), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_0), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_68), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_38), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_61), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_72), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_6), .Y(n_80) );
CKINVDCx14_ASAP7_75t_R g81 ( .A(n_40), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_53), .Y(n_82) );
NOR2xp67_ASAP7_75t_L g83 ( .A(n_30), .B(n_15), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_37), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_54), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_44), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_58), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_15), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_20), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_10), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_27), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_18), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_48), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_39), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_0), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_64), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_22), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_50), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_57), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_2), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_23), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_43), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_65), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_73), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_32), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_56), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_19), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_26), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_21), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_60), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_2), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_47), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_63), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_7), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_84), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_88), .Y(n_121) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_84), .A2(n_29), .B(n_69), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_85), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_96), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_75), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_119), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_119), .Y(n_127) );
INVx2_ASAP7_75t_SL g128 ( .A(n_85), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVxp67_ASAP7_75t_SL g130 ( .A(n_74), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_77), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_100), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_100), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_75), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_96), .Y(n_140) );
NOR2x1_ASAP7_75t_L g141 ( .A(n_83), .B(n_1), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_78), .Y(n_142) );
NOR2x1_ASAP7_75t_L g143 ( .A(n_79), .B(n_94), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_99), .B(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_107), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_108), .B(n_4), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_102), .B(n_5), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_110), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_104), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_81), .B(n_5), .Y(n_152) );
BUFx8_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_112), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_90), .B(n_6), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_90), .B(n_7), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_116), .B(n_8), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_117), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_93), .B(n_8), .Y(n_159) );
OR2x6_ASAP7_75t_L g160 ( .A(n_152), .B(n_80), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_120), .B(n_98), .Y(n_163) );
OAI21xp33_ASAP7_75t_L g164 ( .A1(n_120), .A2(n_82), .B(n_115), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_151), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_122), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_126), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_126), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_130), .B(n_118), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
AND2x4_ASAP7_75t_SL g176 ( .A(n_148), .B(n_140), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_143), .B(n_113), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_124), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_130), .B(n_118), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_143), .B(n_92), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
INVxp67_ASAP7_75t_SL g185 ( .A(n_140), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_124), .B(n_98), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_122), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_152), .A2(n_82), .B1(n_101), .B2(n_97), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_123), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_123), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_123), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_122), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_145), .B(n_97), .Y(n_194) );
AND2x6_ASAP7_75t_L g195 ( .A(n_152), .B(n_148), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g196 ( .A1(n_121), .A2(n_93), .B1(n_109), .B2(n_105), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_135), .Y(n_198) );
INVx5_ASAP7_75t_L g199 ( .A(n_126), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_122), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_121), .B(n_109), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_129), .A2(n_105), .B1(n_114), .B2(n_95), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_153), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_138), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_129), .B(n_106), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_127), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_127), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_128), .Y(n_211) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
INVx5_ASAP7_75t_L g213 ( .A(n_127), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_127), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_138), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_127), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_201), .B(n_148), .Y(n_217) );
INVx5_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_194), .B(n_137), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_170), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_165), .B(n_137), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_195), .A2(n_136), .B1(n_134), .B2(n_133), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_179), .B(n_155), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_179), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_165), .B(n_134), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_187), .Y(n_226) );
BUFx8_ASAP7_75t_L g227 ( .A(n_195), .Y(n_227) );
AO22x1_ASAP7_75t_L g228 ( .A1(n_195), .A2(n_141), .B1(n_76), .B2(n_91), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_212), .B(n_132), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_170), .Y(n_230) );
INVxp67_ASAP7_75t_L g231 ( .A(n_187), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_190), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_195), .B(n_136), .Y(n_233) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_176), .B(n_155), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_169), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_178), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_174), .B(n_146), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_195), .B(n_133), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_176), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_175), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_160), .B(n_141), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_191), .Y(n_243) );
AOI21xp33_ASAP7_75t_L g244 ( .A1(n_182), .A2(n_159), .B(n_157), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_210), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_212), .B(n_128), .Y(n_247) );
BUFx4f_ASAP7_75t_L g248 ( .A(n_195), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_185), .A2(n_144), .B1(n_131), .B2(n_147), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_197), .Y(n_250) );
INVx5_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
AOI22xp5_ASAP7_75t_SL g252 ( .A1(n_166), .A2(n_158), .B1(n_154), .B2(n_150), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_160), .B(n_158), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_210), .Y(n_255) );
INVx5_ASAP7_75t_L g256 ( .A(n_210), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_202), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_177), .B(n_154), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_166), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_206), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_208), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_196), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_210), .Y(n_263) );
BUFx4f_ASAP7_75t_L g264 ( .A(n_160), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_180), .B(n_150), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_215), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_212), .B(n_128), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_214), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_160), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_181), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_177), .B(n_146), .Y(n_272) );
INVx4_ASAP7_75t_L g273 ( .A(n_204), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_184), .B(n_145), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_204), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_221), .A2(n_211), .B(n_161), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_253), .B(n_205), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_224), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_220), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_253), .B(n_177), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_242), .A2(n_183), .B1(n_205), .B2(n_163), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_232), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_225), .A2(n_211), .B(n_161), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_253), .B(n_183), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_232), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_222), .A2(n_183), .B1(n_164), .B2(n_207), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_254), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_220), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_222), .A2(n_189), .B1(n_203), .B2(n_163), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_218), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_218), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_223), .B(n_207), .Y(n_293) );
OR2x6_ASAP7_75t_L g294 ( .A(n_269), .B(n_200), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_217), .B(n_142), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_254), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_242), .A2(n_200), .B1(n_168), .B2(n_188), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_242), .A2(n_200), .B1(n_168), .B2(n_188), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_264), .B(n_142), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_248), .B(n_188), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_264), .B(n_142), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_226), .A2(n_271), .B1(n_231), .B2(n_274), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_230), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_240), .B(n_125), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_259), .Y(n_306) );
INVx5_ASAP7_75t_L g307 ( .A(n_218), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_238), .A2(n_168), .B(n_161), .C(n_188), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_238), .B(n_125), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_218), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_227), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_230), .Y(n_312) );
INVx3_ASAP7_75t_SL g313 ( .A(n_259), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_227), .Y(n_314) );
AOI221xp5_ASAP7_75t_SL g315 ( .A1(n_219), .A2(n_188), .B1(n_161), .B2(n_168), .C(n_193), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_230), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_252), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_248), .A2(n_168), .B1(n_161), .B2(n_193), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_245), .A2(n_186), .B(n_172), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_234), .B(n_139), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_258), .A2(n_139), .B(n_125), .C(n_186), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
OAI21x1_ASAP7_75t_SL g323 ( .A1(n_286), .A2(n_233), .B(n_239), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_305), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_SL g325 ( .A1(n_308), .A2(n_247), .B(n_267), .C(n_229), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_280), .A2(n_234), .B1(n_274), .B2(n_250), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_305), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_313), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_285), .A2(n_274), .B1(n_246), .B2(n_257), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_278), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_287), .A2(n_261), .B1(n_243), .B2(n_260), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_SL g333 ( .A1(n_318), .A2(n_247), .B(n_267), .C(n_229), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_293), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_287), .A2(n_266), .B1(n_272), .B2(n_249), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_303), .A2(n_265), .B1(n_270), .B2(n_237), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_295), .A2(n_265), .B1(n_237), .B2(n_273), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_293), .A2(n_244), .B1(n_262), .B2(n_228), .C(n_241), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_307), .B(n_273), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_317), .A2(n_227), .B1(n_262), .B2(n_273), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_290), .B(n_236), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_313), .A2(n_235), .B1(n_230), .B2(n_275), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_313), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_307), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_309), .A2(n_125), .B1(n_193), .B2(n_127), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_SL g346 ( .A1(n_282), .A2(n_172), .B(n_162), .C(n_167), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_311), .A2(n_275), .B1(n_193), .B2(n_213), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_300), .B(n_275), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_321), .A2(n_193), .B(n_167), .C(n_171), .Y(n_349) );
NOR2xp67_ASAP7_75t_L g350 ( .A(n_306), .B(n_9), .Y(n_350) );
BUFx4f_ASAP7_75t_SL g351 ( .A(n_331), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_345), .A2(n_284), .B(n_276), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_332), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_326), .A2(n_320), .B1(n_300), .B2(n_302), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_338), .A2(n_302), .B1(n_314), .B2(n_311), .Y(n_356) );
CKINVDCx11_ASAP7_75t_R g357 ( .A(n_344), .Y(n_357) );
AOI22xp33_ASAP7_75t_SL g358 ( .A1(n_330), .A2(n_314), .B1(n_277), .B2(n_307), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_328), .A2(n_294), .B1(n_299), .B2(n_282), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_334), .A2(n_281), .B1(n_277), .B2(n_299), .C(n_288), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_294), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_345), .A2(n_325), .B(n_341), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_335), .A2(n_294), .B1(n_277), .B2(n_286), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_343), .Y(n_364) );
BUFx12f_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_336), .A2(n_277), .B1(n_307), .B2(n_294), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_337), .A2(n_319), .B(n_301), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_327), .A2(n_294), .B1(n_292), .B2(n_291), .Y(n_368) );
OAI222xp33_ASAP7_75t_L g369 ( .A1(n_340), .A2(n_283), .B1(n_288), .B2(n_296), .C1(n_301), .C2(n_310), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_348), .B(n_283), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_322), .A2(n_319), .B(n_301), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_322), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_350), .A2(n_296), .B1(n_289), .B2(n_279), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_329), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_370), .B(n_315), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_356), .A2(n_349), .B1(n_347), .B2(n_297), .C(n_298), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_354), .A2(n_349), .B1(n_342), .B2(n_325), .C(n_310), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_360), .B(n_333), .C(n_162), .D(n_171), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_355), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_362), .A2(n_333), .B(n_346), .Y(n_383) );
AO21x2_ASAP7_75t_L g384 ( .A1(n_362), .A2(n_346), .B(n_209), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_365), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_358), .A2(n_291), .B1(n_292), .B2(n_289), .C(n_279), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_353), .A2(n_292), .B1(n_291), .B2(n_209), .C(n_216), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_353), .B(n_316), .Y(n_389) );
OA222x2_ASAP7_75t_L g390 ( .A1(n_361), .A2(n_316), .B1(n_10), .B2(n_11), .C1(n_12), .C2(n_13), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_363), .A2(n_316), .B1(n_275), .B2(n_304), .Y(n_391) );
AOI21xp5_ASAP7_75t_SL g392 ( .A1(n_363), .A2(n_312), .B(n_304), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_372), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_312), .B1(n_304), .B2(n_216), .C(n_199), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_351), .B(n_9), .Y(n_395) );
AOI221xp5_ASAP7_75t_SL g396 ( .A1(n_360), .A2(n_214), .B1(n_304), .B2(n_312), .C(n_263), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_365), .A2(n_312), .B1(n_304), .B2(n_214), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_199), .B(n_213), .C(n_214), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_365), .A2(n_312), .B1(n_199), .B2(n_213), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_372), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g401 ( .A1(n_352), .A2(n_199), .B(n_213), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_369), .A2(n_214), .B1(n_199), .B2(n_213), .C(n_255), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_371), .A2(n_268), .B1(n_263), .B2(n_255), .C(n_245), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_370), .B(n_11), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_361), .A2(n_256), .B1(n_251), .B2(n_268), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_374), .B(n_12), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_374), .B(n_14), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_374), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_385), .B(n_359), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_385), .B(n_364), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
OAI33xp33_ASAP7_75t_L g415 ( .A1(n_395), .A2(n_373), .A3(n_371), .B1(n_376), .B2(n_14), .B3(n_16), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_381), .A2(n_368), .B1(n_373), .B2(n_376), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_386), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_396), .B(n_375), .C(n_376), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_393), .Y(n_420) );
OAI222xp33_ASAP7_75t_L g421 ( .A1(n_390), .A2(n_352), .B1(n_16), .B2(n_17), .C1(n_367), .C2(n_28), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_393), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_383), .A2(n_367), .B(n_17), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_398), .B(n_256), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_404), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_404), .B(n_24), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_410), .B(n_25), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_382), .Y(n_432) );
OAI321xp33_ASAP7_75t_L g433 ( .A1(n_381), .A2(n_31), .A3(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_410), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_380), .A2(n_256), .B1(n_251), .B2(n_46), .C(n_49), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_392), .B(n_42), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_389), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_377), .B(n_45), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_377), .Y(n_442) );
O2A1O1Ixp5_ASAP7_75t_L g443 ( .A1(n_401), .A2(n_51), .B(n_52), .C(n_55), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_408), .B(n_59), .Y(n_444) );
OAI33xp33_ASAP7_75t_L g445 ( .A1(n_390), .A2(n_62), .A3(n_66), .B1(n_70), .B2(n_251), .B3(n_256), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_400), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_408), .B(n_251), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_409), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_407), .B(n_406), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_407), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_384), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_392), .B(n_384), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_384), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_391), .B(n_396), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_391), .B(n_405), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_442), .B(n_402), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_442), .B(n_388), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_440), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_412), .B(n_417), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_412), .B(n_397), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_414), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_434), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_414), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_438), .B(n_399), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_438), .B(n_378), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_434), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_439), .B(n_403), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_413), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_439), .B(n_387), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_426), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_431), .B(n_394), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_424), .A2(n_457), .B(n_437), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_431), .B(n_432), .Y(n_477) );
OAI31xp33_ASAP7_75t_L g478 ( .A1(n_421), .A2(n_411), .A3(n_440), .B(n_444), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_448), .B(n_449), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_432), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_414), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_418), .B(n_425), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_418), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_418), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_448), .B(n_449), .Y(n_486) );
OR2x6_ASAP7_75t_L g487 ( .A(n_437), .B(n_455), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_450), .B(n_416), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_425), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_425), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_446), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_452), .B(n_454), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_452), .B(n_454), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_447), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_451), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_435), .A2(n_455), .B(n_444), .C(n_458), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_450), .B(n_430), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_436), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_436), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_420), .B(n_430), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_422), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_433), .B(n_429), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_429), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_422), .B(n_441), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_441), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_451), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_441), .B(n_451), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_419), .B(n_428), .C(n_456), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_423), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_495), .B(n_423), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_499), .B(n_423), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_478), .A2(n_419), .B(n_443), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_465), .B(n_447), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_466), .B(n_456), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_462), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_469), .B(n_415), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_469), .B(n_453), .Y(n_520) );
NOR2x1_ASAP7_75t_L g521 ( .A(n_472), .B(n_453), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_501), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_477), .Y(n_523) );
AOI211x1_ASAP7_75t_SL g524 ( .A1(n_511), .A2(n_445), .B(n_453), .C(n_505), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_499), .B(n_507), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_497), .B(n_509), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_479), .B(n_486), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_476), .A2(n_498), .B(n_461), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_510), .B(n_488), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_470), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_510), .B(n_494), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_483), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_492), .B(n_494), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_471), .B(n_460), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_477), .B(n_474), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g537 ( .A1(n_473), .A2(n_459), .A3(n_460), .B(n_471), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_492), .B(n_468), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_459), .B(n_463), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_500), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_483), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_506), .B(n_463), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_500), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_474), .B(n_480), .Y(n_544) );
NAND4xp25_ASAP7_75t_L g545 ( .A(n_468), .B(n_512), .C(n_504), .D(n_475), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_503), .B(n_497), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_509), .B(n_487), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_503), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_482), .B(n_491), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_481), .B(n_490), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_475), .A2(n_512), .B(n_487), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_487), .B(n_507), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_482), .B(n_493), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_516), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_536), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_527), .Y(n_557) );
XOR2x2_ASAP7_75t_L g558 ( .A(n_535), .B(n_493), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_526), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_523), .B(n_504), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_539), .B(n_481), .Y(n_561) );
BUFx6f_ASAP7_75t_SL g562 ( .A(n_547), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_542), .B(n_538), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_542), .B(n_489), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_519), .B(n_496), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_520), .B(n_489), .Y(n_566) );
NAND2xp33_ASAP7_75t_SL g567 ( .A(n_547), .B(n_496), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_521), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_549), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_525), .B(n_487), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g571 ( .A1(n_545), .A2(n_508), .B(n_496), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_519), .B(n_508), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_553), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_544), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_527), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_515), .B(n_484), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_531), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_548), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_525), .B(n_484), .Y(n_579) );
NAND2xp33_ASAP7_75t_SL g580 ( .A(n_547), .B(n_485), .Y(n_580) );
OAI332xp33_ASAP7_75t_L g581 ( .A1(n_537), .A2(n_464), .A3(n_467), .B1(n_485), .B2(n_490), .B3(n_502), .C1(n_513), .C2(n_528), .Y(n_581) );
NAND3xp33_ASAP7_75t_SL g582 ( .A(n_524), .B(n_502), .C(n_464), .Y(n_582) );
XNOR2x1_ASAP7_75t_L g583 ( .A(n_530), .B(n_467), .Y(n_583) );
OA22x2_ASAP7_75t_L g584 ( .A1(n_552), .A2(n_551), .B1(n_527), .B2(n_548), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g585 ( .A1(n_529), .A2(n_514), .B(n_552), .C(n_533), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_546), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_534), .B(n_532), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_550), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_533), .A2(n_541), .B(n_514), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
XOR2x2_ASAP7_75t_L g591 ( .A(n_552), .B(n_514), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_540), .A2(n_543), .B(n_522), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_537), .A2(n_519), .B1(n_535), .B2(n_529), .C(n_539), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_545), .A2(n_515), .B(n_529), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_515), .B(n_519), .C(n_421), .Y(n_596) );
XNOR2xp5_ASAP7_75t_L g597 ( .A(n_530), .B(n_472), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_578), .Y(n_598) );
A2O1A1Ixp33_ASAP7_75t_L g599 ( .A1(n_595), .A2(n_594), .B(n_585), .C(n_596), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_578), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_576), .B(n_557), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_594), .A2(n_565), .B1(n_584), .B2(n_572), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_584), .A2(n_565), .B(n_572), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g604 ( .A1(n_581), .A2(n_580), .B(n_571), .C(n_567), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_590), .Y(n_605) );
AOI311xp33_ASAP7_75t_L g606 ( .A1(n_589), .A2(n_555), .A3(n_569), .B(n_573), .C(n_592), .Y(n_606) );
AOI321xp33_ASAP7_75t_L g607 ( .A1(n_563), .A2(n_570), .A3(n_574), .B1(n_564), .B2(n_561), .C(n_588), .Y(n_607) );
O2A1O1Ixp5_ASAP7_75t_L g608 ( .A1(n_580), .A2(n_567), .B(n_559), .C(n_556), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_586), .Y(n_609) );
BUFx8_ASAP7_75t_L g610 ( .A(n_562), .Y(n_610) );
OAI211xp5_ASAP7_75t_SL g611 ( .A1(n_599), .A2(n_568), .B(n_575), .C(n_560), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_608), .A2(n_597), .B(n_558), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_605), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_602), .A2(n_554), .B1(n_582), .B2(n_568), .C(n_577), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_598), .Y(n_615) );
AOI211x1_ASAP7_75t_L g616 ( .A1(n_603), .A2(n_593), .B(n_579), .C(n_566), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_604), .A2(n_610), .B1(n_601), .B2(n_609), .Y(n_617) );
NOR2xp67_ASAP7_75t_SL g618 ( .A(n_612), .B(n_610), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_617), .Y(n_619) );
AOI211xp5_ASAP7_75t_SL g620 ( .A1(n_614), .A2(n_604), .B(n_606), .C(n_601), .Y(n_620) );
NOR4xp25_ASAP7_75t_L g621 ( .A(n_611), .B(n_607), .C(n_600), .D(n_593), .Y(n_621) );
NOR2x1p5_ASAP7_75t_L g622 ( .A(n_618), .B(n_613), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_619), .A2(n_615), .B1(n_562), .B2(n_591), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_622), .Y(n_624) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_623), .A2(n_621), .B(n_618), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_625), .A2(n_620), .B1(n_616), .B2(n_587), .Y(n_626) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_626), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_627), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_628), .A2(n_624), .B(n_583), .Y(n_629) );
endmodule