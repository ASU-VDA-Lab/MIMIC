module fake_jpeg_18863_n_324 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_10),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx6p67_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_12),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_16),
.Y(n_36)
);

AO22x2_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_16),
.B1(n_14),
.B2(n_17),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_32),
.B1(n_27),
.B2(n_31),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_62),
.Y(n_76)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_57),
.B1(n_38),
.B2(n_40),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_35),
.CI(n_26),
.CON(n_81),
.SN(n_81)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_13),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_78),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_26),
.C(n_46),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_77),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_26),
.C(n_30),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_36),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_59),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_40),
.B1(n_35),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_42),
.B1(n_39),
.B2(n_44),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_62),
.B1(n_51),
.B2(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_38),
.B1(n_66),
.B2(n_70),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_59),
.B(n_35),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_78),
.B(n_79),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_101),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_104),
.B1(n_108),
.B2(n_38),
.Y(n_109)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_19),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_22),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_35),
.B(n_50),
.C(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_38),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_58),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_79),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_42),
.B1(n_38),
.B2(n_51),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_109),
.A2(n_131),
.B1(n_53),
.B2(n_34),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_116),
.B(n_133),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_137),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_75),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_114),
.B(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_126),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_85),
.B(n_80),
.C(n_97),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_92),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_129),
.Y(n_172)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_103),
.B1(n_108),
.B2(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_102),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_69),
.B1(n_71),
.B2(n_34),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_120),
.B2(n_129),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_98),
.B1(n_66),
.B2(n_70),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_88),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_95),
.C(n_89),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_147),
.C(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_165),
.B1(n_113),
.B2(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_95),
.C(n_77),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_101),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_139),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_99),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_156),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_90),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_169),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_69),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_157),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_67),
.C(n_26),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_21),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_158),
.B(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_33),
.B1(n_58),
.B2(n_20),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_164),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_80),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_166),
.B1(n_165),
.B2(n_169),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_85),
.B(n_22),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_15),
.B(n_12),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_58),
.C(n_61),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_61),
.C(n_23),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_19),
.B1(n_85),
.B2(n_12),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_33),
.B1(n_85),
.B2(n_20),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_49),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_167),
.B(n_115),
.Y(n_179)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_110),
.B(n_33),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_183),
.B(n_14),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_14),
.B1(n_17),
.B2(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_109),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_15),
.B1(n_61),
.B2(n_24),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_15),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_191),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_14),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_148),
.B(n_8),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_149),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_23),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_14),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_170),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_202),
.A2(n_143),
.B(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_147),
.C(n_173),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_207),
.C(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_213),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_173),
.C(n_142),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_140),
.B1(n_157),
.B2(n_142),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_182),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_177),
.A2(n_140),
.B1(n_162),
.B2(n_23),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_9),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_140),
.C(n_23),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_224),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_24),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_192),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_225),
.B1(n_180),
.B2(n_196),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_17),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_188),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_178),
.B1(n_182),
.B2(n_181),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_249),
.B1(n_222),
.B2(n_219),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_233),
.B(n_226),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_217),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_178),
.B1(n_190),
.B2(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_224),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_174),
.B1(n_198),
.B2(n_175),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_175),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_174),
.B1(n_199),
.B2(n_191),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_216),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_232),
.B(n_240),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_204),
.C(n_207),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_230),
.C(n_236),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_261),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_223),
.B1(n_225),
.B2(n_245),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_218),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_197),
.B(n_195),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_265),
.B(n_230),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_234),
.B1(n_249),
.B2(n_228),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_277),
.B1(n_6),
.B2(n_2),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_273),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_241),
.C(n_244),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_201),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_252),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_6),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_284),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_290),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_255),
.B1(n_264),
.B2(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_7),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_254),
.C(n_266),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_274),
.B(n_266),
.Y(n_291)
);

FAx1_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_283),
.CI(n_288),
.CON(n_301),
.SN(n_301)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_274),
.Y(n_293)
);

OAI322xp33_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_268),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_300),
.B(n_304),
.Y(n_311)
);

INVx11_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_297),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_291),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_287),
.B(n_7),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_7),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_3),
.C(n_4),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_310),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_4),
.C(n_5),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_301),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_4),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_298),
.C(n_302),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_294),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_308),
.A3(n_311),
.B1(n_309),
.B2(n_312),
.C1(n_11),
.C2(n_10),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_316),
.B(n_315),
.Y(n_320)
);

AOI321xp33_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_318),
.A3(n_309),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_5),
.B(n_0),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_5),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_0),
.Y(n_324)
);


endmodule