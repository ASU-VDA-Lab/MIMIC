module real_jpeg_28808_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_60),
.Y(n_106)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_2),
.B(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_2),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_2),
.A2(n_24),
.B(n_76),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_96),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_51),
.B(n_64),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_2),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_2),
.A2(n_57),
.B1(n_88),
.B2(n_163),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_3),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_6),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_8),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_149)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_71),
.Y(n_79)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_14),
.A2(n_27),
.B1(n_94),
.B2(n_95),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_14),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_163)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_15),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_19),
.B(n_83),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.C(n_73),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_20),
.A2(n_21),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_22),
.B(n_39),
.C(n_45),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_23),
.A2(n_28),
.B1(n_33),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_42),
.Y(n_92)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_25),
.A2(n_34),
.A3(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_25),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_91)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_28),
.A2(n_33),
.B1(n_36),
.B2(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_30),
.B(n_35),
.Y(n_77)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_33),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_35),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_35),
.A2(n_65),
.B(n_96),
.C(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_41),
.A2(n_93),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_41),
.A2(n_42),
.B(n_94),
.C(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_94),
.Y(n_97)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_54),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_49),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_47),
.B(n_79),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_47),
.A2(n_55),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_56),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_51),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_50),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_57),
.A2(n_88),
.B1(n_155),
.B2(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_57),
.B(n_96),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_61),
.B(n_73),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B(n_69),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_66),
.B1(n_67),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_62),
.A2(n_66),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_62),
.A2(n_66),
.B1(n_127),
.B2(n_138),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_66),
.B(n_96),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_78),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_100),
.B1(n_101),
.B2(n_114),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_98),
.B2(n_99),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

HAxp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.CON(n_93),
.SN(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_131),
.B(n_177),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_119),
.B(n_128),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_125),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_121),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_171),
.B(n_176),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_151),
.B(n_170),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_147),
.C(n_148),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_159),
.B(n_169),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_153),
.B(n_157),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_164),
.B(n_168),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);


endmodule