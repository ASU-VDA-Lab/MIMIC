module fake_jpeg_17547_n_270 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx12f_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_25),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_21),
.B1(n_34),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_50),
.B1(n_55),
.B2(n_58),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_59),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_2),
.B(n_3),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_2),
.B(n_4),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_44),
.B1(n_36),
.B2(n_39),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_65),
.Y(n_84)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_72),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_42),
.Y(n_72)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_7),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_28),
.B1(n_24),
.B2(n_30),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_76),
.A2(n_77),
.B1(n_83),
.B2(n_6),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_28),
.B1(n_24),
.B2(n_30),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_32),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_17),
.B1(n_23),
.B2(n_29),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_45),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_7),
.Y(n_124)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_88),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_67),
.B1(n_63),
.B2(n_65),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_97),
.B1(n_32),
.B2(n_29),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_17),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_45),
.B(n_32),
.C(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_22),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_104),
.B1(n_68),
.B2(n_96),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_54),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_125),
.B(n_72),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_27),
.C(n_23),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_27),
.Y(n_106)
);

AO21x2_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_23),
.B(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_95),
.B1(n_79),
.B2(n_90),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_120),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_82),
.B(n_22),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_124),
.B(n_91),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_73),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_93),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_7),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_126),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_132),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_80),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_137),
.C(n_145),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_74),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_138),
.B(n_143),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_87),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_142),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_85),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_103),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_94),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_144),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_94),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_97),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_111),
.B1(n_116),
.B2(n_110),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_90),
.C(n_95),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_152),
.C(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_75),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_117),
.C(n_111),
.D(n_116),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_156),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_168),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_111),
.B(n_103),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_177),
.B(n_119),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_102),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_173),
.B1(n_177),
.B2(n_174),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_102),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_89),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_88),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_111),
.B(n_107),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_107),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_127),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_152),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_183),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_186),
.B1(n_169),
.B2(n_164),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_188),
.C(n_193),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_131),
.B1(n_111),
.B2(n_149),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_138),
.C(n_134),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_128),
.C(n_104),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_203),
.B(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_86),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_172),
.CI(n_168),
.CON(n_198),
.SN(n_198)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_191),
.CI(n_201),
.CON(n_210),
.SN(n_210)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_88),
.C(n_147),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_200),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_105),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_212),
.B1(n_215),
.B2(n_195),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_221),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_217),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_166),
.B1(n_203),
.B2(n_184),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_162),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_158),
.B(n_175),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_165),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_158),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_156),
.B(n_198),
.C(n_201),
.D(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_167),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_188),
.C(n_185),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_216),
.C(n_193),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_232),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_212),
.B1(n_220),
.B2(n_210),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_231),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_215),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_175),
.C(n_179),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_161),
.C(n_155),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_235),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_210),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_181),
.C(n_160),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_11),
.C(n_14),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_218),
.B(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_246),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_214),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_224),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_224),
.A2(n_206),
.B(n_181),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_249),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_12),
.B(n_16),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_238),
.C(n_237),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_11),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_14),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_8),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_240),
.B(n_239),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_237),
.B(n_93),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_254),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_9),
.A3(n_10),
.B1(n_255),
.B2(n_257),
.C1(n_258),
.C2(n_261),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_267),
.B1(n_9),
.B2(n_10),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g268 ( 
.A(n_266),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);


endmodule