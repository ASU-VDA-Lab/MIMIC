module real_aes_486_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_832, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_833, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_832;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_833;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_626;
wire n_400;
wire n_539;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g231 ( .A(n_0), .B(n_153), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_1), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g146 ( .A(n_2), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_3), .B(n_159), .Y(n_172) );
NAND2xp33_ASAP7_75t_SL g223 ( .A(n_4), .B(n_157), .Y(n_223) );
INVx1_ASAP7_75t_L g204 ( .A(n_5), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_6), .B(n_177), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_7), .A2(n_121), .B1(n_122), .B2(n_124), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_7), .Y(n_121) );
INVx1_ASAP7_75t_L g530 ( .A(n_8), .Y(n_530) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_9), .Y(n_111) );
AND2x2_ASAP7_75t_L g170 ( .A(n_10), .B(n_163), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_11), .Y(n_497) );
INVx2_ASAP7_75t_L g164 ( .A(n_12), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_13), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_14), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_14), .B(n_27), .Y(n_726) );
INVx1_ASAP7_75t_L g558 ( .A(n_15), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g815 ( .A1(n_16), .A2(n_27), .B1(n_780), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_16), .Y(n_816) );
AOI221x1_ASAP7_75t_L g217 ( .A1(n_17), .A2(n_141), .B1(n_218), .B2(n_220), .C(n_222), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_18), .B(n_159), .Y(n_192) );
INVx1_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
INVx1_ASAP7_75t_L g556 ( .A(n_20), .Y(n_556) );
INVx1_ASAP7_75t_SL g479 ( .A(n_21), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_22), .B(n_160), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_23), .A2(n_141), .B(n_174), .Y(n_173) );
AOI221xp5_ASAP7_75t_SL g184 ( .A1(n_24), .A2(n_40), .B1(n_141), .B2(n_159), .C(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_25), .B(n_153), .Y(n_175) );
AOI33xp33_ASAP7_75t_L g516 ( .A1(n_26), .A2(n_53), .A3(n_207), .B1(n_213), .B2(n_517), .B3(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g780 ( .A(n_27), .Y(n_780) );
INVx1_ASAP7_75t_L g490 ( .A(n_28), .Y(n_490) );
OR2x2_ASAP7_75t_L g165 ( .A(n_29), .B(n_93), .Y(n_165) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_29), .A2(n_93), .B(n_164), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_30), .B(n_149), .Y(n_196) );
INVxp67_ASAP7_75t_L g216 ( .A(n_31), .Y(n_216) );
AND2x2_ASAP7_75t_L g247 ( .A(n_32), .B(n_162), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_33), .B(n_205), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_34), .A2(n_141), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_35), .B(n_149), .Y(n_186) );
AND2x2_ASAP7_75t_L g142 ( .A(n_36), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g157 ( .A(n_36), .B(n_146), .Y(n_157) );
INVx1_ASAP7_75t_L g212 ( .A(n_36), .Y(n_212) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_37), .B(n_110), .C(n_112), .Y(n_109) );
OR2x6_ASAP7_75t_L g789 ( .A(n_37), .B(n_790), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_38), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_39), .B(n_205), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_41), .A2(n_177), .B1(n_221), .B2(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_42), .B(n_548), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_43), .A2(n_83), .B1(n_141), .B2(n_210), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_44), .B(n_160), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_45), .B(n_153), .Y(n_245) );
INVx1_ASAP7_75t_L g787 ( .A(n_46), .Y(n_787) );
XNOR2xp5_ASAP7_75t_L g818 ( .A(n_47), .B(n_87), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_48), .B(n_197), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_49), .B(n_160), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_50), .Y(n_543) );
AND2x2_ASAP7_75t_L g234 ( .A(n_51), .B(n_162), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_52), .B(n_162), .Y(n_188) );
XOR2xp5_ASAP7_75t_L g810 ( .A(n_52), .B(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_54), .B(n_160), .Y(n_508) );
INVx1_ASAP7_75t_L g145 ( .A(n_55), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_55), .Y(n_155) );
AND2x2_ASAP7_75t_L g509 ( .A(n_56), .B(n_162), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_57), .A2(n_76), .B1(n_205), .B2(n_210), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_58), .B(n_205), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_59), .B(n_159), .Y(n_246) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_60), .A2(n_120), .B1(n_125), .B2(n_126), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_60), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_61), .B(n_221), .Y(n_499) );
AOI21xp5_ASAP7_75t_SL g468 ( .A1(n_62), .A2(n_210), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g166 ( .A(n_63), .B(n_162), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_64), .B(n_149), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_65), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_66), .B(n_163), .Y(n_199) );
INVx1_ASAP7_75t_L g553 ( .A(n_67), .Y(n_553) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_68), .B(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_69), .A2(n_141), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g507 ( .A(n_70), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_71), .B(n_149), .Y(n_176) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_72), .B(n_197), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_73), .A2(n_210), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g143 ( .A(n_74), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_74), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_75), .B(n_205), .Y(n_519) );
AND2x2_ASAP7_75t_L g481 ( .A(n_77), .B(n_220), .Y(n_481) );
INVx1_ASAP7_75t_L g554 ( .A(n_78), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_79), .A2(n_210), .B(n_478), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_80), .A2(n_210), .B(n_280), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_81), .B(n_159), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_82), .A2(n_86), .B1(n_159), .B2(n_205), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_84), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g791 ( .A(n_84), .Y(n_791) );
AND2x2_ASAP7_75t_SL g466 ( .A(n_85), .B(n_220), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_88), .A2(n_210), .B1(n_514), .B2(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_89), .B(n_153), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_90), .B(n_153), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g792 ( .A(n_91), .B(n_793), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_92), .A2(n_141), .B(n_147), .Y(n_140) );
INVx1_ASAP7_75t_L g470 ( .A(n_94), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_95), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g520 ( .A(n_96), .B(n_220), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_97), .Y(n_828) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_98), .A2(n_488), .B(n_489), .C(n_491), .Y(n_487) );
INVxp67_ASAP7_75t_L g219 ( .A(n_99), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_100), .B(n_159), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_101), .B(n_149), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_102), .A2(n_141), .B(n_194), .Y(n_193) );
BUFx2_ASAP7_75t_SL g785 ( .A(n_103), .Y(n_785) );
BUFx2_ASAP7_75t_L g802 ( .A(n_103), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_104), .B(n_160), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_116), .B(n_827), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx4f_ASAP7_75t_SL g830 ( .A(n_108), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_109), .B(n_114), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_112), .B(n_780), .Y(n_779) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_113), .Y(n_129) );
OR2x2_ASAP7_75t_L g788 ( .A(n_113), .B(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_113), .B(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_115), .B(n_791), .Y(n_790) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_803), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_781), .B(n_797), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_127), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g826 ( .A(n_119), .Y(n_826) );
INVxp33_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
INVx1_ASAP7_75t_L g124 ( .A(n_122), .Y(n_124) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_128), .Y(n_825) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_456), .Y(n_128) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_395), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_288), .C(n_339), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_178), .B(n_235), .C(n_266), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_167), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_137), .B(n_240), .Y(n_403) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g248 ( .A(n_138), .B(n_169), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_138), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g265 ( .A(n_138), .B(n_255), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_138), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g302 ( .A(n_138), .B(n_278), .Y(n_302) );
INVx2_ASAP7_75t_L g328 ( .A(n_138), .Y(n_328) );
AND2x4_ASAP7_75t_L g337 ( .A(n_138), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g442 ( .A(n_138), .B(n_309), .Y(n_442) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_161), .B(n_166), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_158), .Y(n_139) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
BUFx3_ASAP7_75t_L g209 ( .A(n_142), .Y(n_209) );
AND2x6_ASAP7_75t_L g153 ( .A(n_143), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g214 ( .A(n_143), .Y(n_214) );
AND2x4_ASAP7_75t_L g210 ( .A(n_144), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g149 ( .A(n_145), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_156), .Y(n_147) );
INVxp67_ASAP7_75t_L g559 ( .A(n_149), .Y(n_559) );
AND2x4_ASAP7_75t_L g160 ( .A(n_150), .B(n_154), .Y(n_160) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVxp67_ASAP7_75t_L g557 ( .A(n_153), .Y(n_557) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_156), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_156), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_156), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_156), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_156), .A2(n_244), .B(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_156), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_156), .A2(n_471), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_156), .A2(n_471), .B(n_507), .C(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g514 ( .A(n_156), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_156), .A2(n_471), .B(n_530), .C(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_156), .A2(n_546), .B(n_547), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_156), .B(n_177), .Y(n_560) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g159 ( .A(n_157), .B(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_157), .Y(n_491) );
INVx1_ASAP7_75t_L g224 ( .A(n_160), .Y(n_224) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_161), .A2(n_241), .B(n_247), .Y(n_240) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_161), .A2(n_241), .B(n_247), .Y(n_255) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_161), .A2(n_475), .B(n_481), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_162), .Y(n_161) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_162), .A2(n_184), .B(n_188), .Y(n_183) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_164), .B(n_165), .Y(n_163) );
AND2x4_ASAP7_75t_L g177 ( .A(n_164), .B(n_165), .Y(n_177) );
AND2x2_ASAP7_75t_L g326 ( .A(n_167), .B(n_327), .Y(n_326) );
OAI32xp33_ASAP7_75t_L g409 ( .A1(n_167), .A2(n_331), .A3(n_335), .B1(n_342), .B2(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_167), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g263 ( .A(n_168), .B(n_264), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_168), .B(n_258), .C(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g362 ( .A(n_168), .B(n_265), .Y(n_362) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_169), .Y(n_252) );
INVx5_ASAP7_75t_L g287 ( .A(n_169), .Y(n_287) );
AND2x4_ASAP7_75t_L g343 ( .A(n_169), .B(n_255), .Y(n_343) );
OR2x2_ASAP7_75t_L g358 ( .A(n_169), .B(n_278), .Y(n_358) );
OR2x2_ASAP7_75t_L g384 ( .A(n_169), .B(n_240), .Y(n_384) );
AND2x2_ASAP7_75t_L g392 ( .A(n_169), .B(n_338), .Y(n_392) );
AND2x4_ASAP7_75t_SL g417 ( .A(n_169), .B(n_337), .Y(n_417) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_177), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_177), .B(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_177), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_177), .B(n_219), .Y(n_218) );
NOR3xp33_ASAP7_75t_L g222 ( .A(n_177), .B(n_223), .C(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_177), .A2(n_468), .B(n_473), .Y(n_467) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_179), .B(n_337), .Y(n_413) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_189), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_180), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OR2x6_ASAP7_75t_SL g237 ( .A(n_181), .B(n_238), .Y(n_237) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g262 ( .A(n_182), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_182), .B(n_297), .Y(n_315) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_182), .Y(n_453) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g270 ( .A(n_183), .Y(n_270) );
AND2x2_ASAP7_75t_L g295 ( .A(n_183), .B(n_226), .Y(n_295) );
INVx2_ASAP7_75t_L g323 ( .A(n_183), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_183), .B(n_190), .Y(n_364) );
BUFx3_ASAP7_75t_L g388 ( .A(n_183), .Y(n_388) );
OR2x2_ASAP7_75t_L g400 ( .A(n_183), .B(n_190), .Y(n_400) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_183), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_189), .A2(n_431), .B1(n_434), .B2(n_435), .Y(n_430) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_200), .Y(n_189) );
INVx1_ASAP7_75t_L g258 ( .A(n_190), .Y(n_258) );
OR2x2_ASAP7_75t_L g269 ( .A(n_190), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g276 ( .A(n_190), .Y(n_276) );
AND2x4_ASAP7_75t_SL g293 ( .A(n_190), .B(n_201), .Y(n_293) );
AND2x4_ASAP7_75t_L g298 ( .A(n_190), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g307 ( .A(n_190), .Y(n_307) );
OR2x2_ASAP7_75t_L g313 ( .A(n_190), .B(n_201), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_190), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_190), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_190), .B(n_295), .Y(n_429) );
OR2x2_ASAP7_75t_L g445 ( .A(n_190), .B(n_348), .Y(n_445) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_199), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_197), .Y(n_191) );
INVx2_ASAP7_75t_SL g280 ( .A(n_197), .Y(n_280) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_197), .A2(n_528), .B(n_532), .Y(n_527) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g221 ( .A(n_198), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_200), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g271 ( .A(n_200), .Y(n_271) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_200), .B(n_262), .Y(n_378) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_225), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_201), .B(n_226), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_201), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_201), .B(n_270), .Y(n_274) );
INVx3_ASAP7_75t_L g299 ( .A(n_201), .Y(n_299) );
INVx1_ASAP7_75t_L g332 ( .A(n_201), .Y(n_332) );
AND2x2_ASAP7_75t_L g412 ( .A(n_201), .B(n_276), .Y(n_412) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_217), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B1(n_210), .B2(n_215), .Y(n_202) );
INVx1_ASAP7_75t_L g500 ( .A(n_205), .Y(n_500) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_209), .Y(n_205) );
INVx1_ASAP7_75t_L g541 ( .A(n_206), .Y(n_541) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
OR2x6_ASAP7_75t_L g471 ( .A(n_207), .B(n_214), .Y(n_471) );
INVxp33_ASAP7_75t_L g517 ( .A(n_207), .Y(n_517) );
INVx1_ASAP7_75t_L g542 ( .A(n_209), .Y(n_542) );
INVxp67_ASAP7_75t_L g498 ( .A(n_210), .Y(n_498) );
NOR2x1p5_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx1_ASAP7_75t_L g518 ( .A(n_213), .Y(n_518) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_220), .A2(n_487), .B1(n_492), .B2(n_493), .Y(n_486) );
INVx3_ASAP7_75t_L g493 ( .A(n_220), .Y(n_493) );
INVx4_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AOI21x1_ASAP7_75t_L g227 ( .A1(n_221), .A2(n_228), .B(n_234), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_221), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_224), .B(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_224), .A2(n_471), .B1(n_553), .B2(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_226), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g297 ( .A(n_226), .Y(n_297) );
AND2x2_ASAP7_75t_L g322 ( .A(n_226), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g348 ( .A(n_226), .B(n_270), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_226), .B(n_299), .Y(n_365) );
INVx1_ASAP7_75t_L g371 ( .A(n_226), .Y(n_371) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
AOI222xp33_ASAP7_75t_SL g235 ( .A1(n_236), .A2(n_239), .B1(n_249), .B2(n_256), .C1(n_259), .C2(n_263), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_248), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_240), .B(n_309), .Y(n_360) );
AND2x4_ASAP7_75t_L g376 ( .A(n_240), .B(n_287), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_246), .Y(n_241) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_251), .B(n_253), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g301 ( .A(n_252), .B(n_302), .Y(n_301) );
AOI222xp33_ASAP7_75t_L g266 ( .A1(n_253), .A2(n_267), .B1(n_272), .B2(n_277), .C1(n_285), .C2(n_832), .Y(n_266) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g405 ( .A(n_254), .B(n_309), .Y(n_405) );
OR2x2_ASAP7_75t_L g448 ( .A(n_254), .B(n_354), .Y(n_448) );
AND2x2_ASAP7_75t_L g277 ( .A(n_255), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g338 ( .A(n_255), .Y(n_338) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_255), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g366 ( .A1(n_256), .A2(n_367), .B(n_372), .C(n_373), .Y(n_366) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g394 ( .A(n_258), .Y(n_394) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g324 ( .A(n_263), .Y(n_324) );
AND2x2_ASAP7_75t_L g308 ( .A(n_264), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g317 ( .A(n_264), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI31xp33_ASAP7_75t_L g359 ( .A1(n_267), .A2(n_285), .A3(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_268), .A2(n_318), .B(n_362), .C(n_363), .Y(n_361) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
OR2x2_ASAP7_75t_L g350 ( .A(n_269), .B(n_299), .Y(n_350) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
BUFx2_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
AND2x2_ASAP7_75t_L g327 ( .A(n_278), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_279), .Y(n_309) );
AOI21x1_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_284), .Y(n_279) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_280), .A2(n_512), .B(n_520), .Y(n_511) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_280), .A2(n_512), .B(n_520), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_287), .B(n_344), .Y(n_436) );
OAI211xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_300), .B(n_303), .C(n_325), .Y(n_288) );
INVxp33_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_291), .B(n_296), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g329 ( .A(n_293), .B(n_322), .Y(n_329) );
OR2x2_ASAP7_75t_L g305 ( .A(n_294), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g335 ( .A(n_294), .B(n_309), .Y(n_335) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g411 ( .A(n_295), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g434 ( .A(n_296), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_298), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_298), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g446 ( .A(n_298), .B(n_322), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_298), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g389 ( .A(n_299), .B(n_371), .Y(n_389) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AOI322xp5_ASAP7_75t_L g443 ( .A1(n_302), .A2(n_322), .A3(n_376), .B1(n_401), .B2(n_444), .C1(n_446), .C2(n_447), .Y(n_443) );
AOI211xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_308), .B(n_310), .C(n_319), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_306), .B(n_334), .Y(n_356) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g321 ( .A(n_307), .B(n_322), .Y(n_321) );
NOR2x1p5_ASAP7_75t_L g387 ( .A(n_307), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_307), .Y(n_420) );
O2A1O1Ixp33_ASAP7_75t_L g325 ( .A1(n_308), .A2(n_326), .B(n_329), .C(n_330), .Y(n_325) );
AND2x4_ASAP7_75t_L g344 ( .A(n_309), .B(n_328), .Y(n_344) );
INVx2_ASAP7_75t_L g354 ( .A(n_309), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_309), .B(n_343), .Y(n_374) );
AND2x2_ASAP7_75t_L g416 ( .A(n_309), .B(n_417), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_309), .B(n_433), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_309), .B(n_337), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B(n_316), .Y(n_310) );
AND2x2_ASAP7_75t_L g406 ( .A(n_312), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g334 ( .A(n_315), .Y(n_334) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_327), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g421 ( .A(n_327), .Y(n_421) );
O2A1O1Ixp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_333), .B(n_335), .C(n_336), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_334), .Y(n_418) );
INVx3_ASAP7_75t_SL g433 ( .A(n_337), .Y(n_433) );
NAND5xp2_ASAP7_75t_L g339 ( .A(n_340), .B(n_359), .C(n_366), .D(n_379), .E(n_390), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B1(n_349), .B2(n_351), .C1(n_355), .C2(n_357), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_342), .A2(n_423), .B1(n_427), .B2(n_428), .Y(n_422) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g372 ( .A(n_343), .B(n_344), .Y(n_372) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_353), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_354), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g391 ( .A(n_354), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g402 ( .A(n_354), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g432 ( .A(n_358), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_377), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_376), .A2(n_380), .B1(n_381), .B2(n_385), .Y(n_379) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g393 ( .A(n_378), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g398 ( .A(n_380), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_SL g426 ( .A(n_389), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_414), .C(n_437), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_413), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .B1(n_404), .B2(n_406), .C(n_409), .Y(n_397) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g438 ( .A(n_400), .B(n_426), .Y(n_438) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
OAI321xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_418), .A3(n_419), .B1(n_421), .B2(n_422), .C(n_430), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_428), .A2(n_450), .B1(n_454), .B2(n_455), .Y(n_449) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_439), .B(n_443), .C(n_449), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_777), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_727), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_667), .B(n_726), .Y(n_458) );
NOR3xp33_ASAP7_75t_L g777 ( .A(n_459), .B(n_728), .C(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g821 ( .A(n_459), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_631), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_572), .C(n_601), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_462), .B(n_561), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_482), .B1(n_521), .B2(n_533), .Y(n_462) );
NAND2x1_ASAP7_75t_L g763 ( .A(n_463), .B(n_562), .Y(n_763) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_474), .Y(n_464) );
INVx2_ASAP7_75t_L g535 ( .A(n_465), .Y(n_535) );
INVx4_ASAP7_75t_L g577 ( .A(n_465), .Y(n_577) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_465), .Y(n_597) );
AND2x4_ASAP7_75t_L g608 ( .A(n_465), .B(n_576), .Y(n_608) );
AND2x2_ASAP7_75t_L g614 ( .A(n_465), .B(n_538), .Y(n_614) );
NOR2x1_ASAP7_75t_SL g687 ( .A(n_465), .B(n_549), .Y(n_687) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVxp67_ASAP7_75t_L g488 ( .A(n_471), .Y(n_488) );
INVx2_ASAP7_75t_L g548 ( .A(n_471), .Y(n_548) );
INVx2_ASAP7_75t_L g580 ( .A(n_474), .Y(n_580) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_474), .Y(n_594) );
INVx1_ASAP7_75t_L g605 ( .A(n_474), .Y(n_605) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_474), .Y(n_617) );
AND2x2_ASAP7_75t_L g649 ( .A(n_474), .B(n_549), .Y(n_649) );
INVx1_ASAP7_75t_L g675 ( .A(n_474), .Y(n_675) );
AND2x2_ASAP7_75t_L g737 ( .A(n_474), .B(n_565), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_501), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g630 ( .A(n_484), .B(n_569), .Y(n_630) );
INVx2_ASAP7_75t_L g672 ( .A(n_484), .Y(n_672) );
AND2x2_ASAP7_75t_L g774 ( .A(n_484), .B(n_501), .Y(n_774) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_485), .B(n_524), .Y(n_568) );
INVx2_ASAP7_75t_L g589 ( .A(n_485), .Y(n_589) );
AND2x4_ASAP7_75t_L g611 ( .A(n_485), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g646 ( .A(n_485), .Y(n_646) );
AND2x2_ASAP7_75t_L g770 ( .A(n_485), .B(n_527), .Y(n_770) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_493), .A2(n_503), .B(n_509), .Y(n_502) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_493), .A2(n_503), .B(n_509), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g744 ( .A(n_501), .Y(n_744) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
NOR2xp67_ASAP7_75t_L g619 ( .A(n_502), .B(n_589), .Y(n_619) );
AND2x2_ASAP7_75t_L g624 ( .A(n_502), .B(n_589), .Y(n_624) );
INVx2_ASAP7_75t_L g637 ( .A(n_502), .Y(n_637) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_502), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AND2x4_ASAP7_75t_L g610 ( .A(n_510), .B(n_523), .Y(n_610) );
AND2x2_ASAP7_75t_L g625 ( .A(n_510), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g680 ( .A(n_510), .Y(n_680) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_511), .B(n_527), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_511), .B(n_524), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVxp33_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx3_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
AND2x2_ASAP7_75t_L g698 ( .A(n_524), .B(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g641 ( .A(n_525), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_525), .B(n_680), .Y(n_721) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g588 ( .A(n_526), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g569 ( .A(n_527), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g612 ( .A(n_527), .Y(n_612) );
INVxp67_ASAP7_75t_L g626 ( .A(n_527), .Y(n_626) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_527), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_527), .Y(n_703) );
INVx1_ASAP7_75t_L g681 ( .A(n_533), .Y(n_681) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_534), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g723 ( .A(n_535), .B(n_564), .Y(n_723) );
OR2x2_ASAP7_75t_L g775 ( .A(n_536), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g674 ( .A(n_537), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g710 ( .A(n_537), .B(n_597), .Y(n_710) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_549), .Y(n_537) );
AND2x4_ASAP7_75t_L g564 ( .A(n_538), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g576 ( .A(n_538), .Y(n_576) );
INVx2_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_538), .Y(n_719) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .C(n_543), .Y(n_540) );
INVx3_ASAP7_75t_L g565 ( .A(n_549), .Y(n_565) );
INVx2_ASAP7_75t_L g659 ( .A(n_549), .Y(n_659) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .B(n_560), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_566), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_563), .B(n_639), .Y(n_656) );
NOR2x1_ASAP7_75t_L g748 ( .A(n_563), .B(n_577), .Y(n_748) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_564), .B(n_639), .Y(n_725) );
AND2x2_ASAP7_75t_L g592 ( .A(n_565), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g606 ( .A(n_565), .Y(n_606) );
AOI22xp5_ASAP7_75t_SL g654 ( .A1(n_566), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_567), .B(n_625), .Y(n_651) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g759 ( .A(n_568), .B(n_600), .Y(n_759) );
AND2x2_ASAP7_75t_L g582 ( .A(n_569), .B(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g618 ( .A(n_569), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g761 ( .A(n_569), .B(n_672), .Y(n_761) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g636 ( .A(n_571), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g662 ( .A(n_571), .Y(n_662) );
AND2x2_ASAP7_75t_L g697 ( .A(n_571), .B(n_589), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_581), .B1(n_585), .B2(n_590), .C(n_595), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
INVx1_ASAP7_75t_L g653 ( .A(n_575), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_575), .B(n_649), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_575), .B(n_737), .Y(n_736) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2xp67_ASAP7_75t_SL g621 ( .A(n_577), .B(n_622), .Y(n_621) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_577), .Y(n_634) );
AND2x4_ASAP7_75t_SL g718 ( .A(n_577), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g765 ( .A(n_577), .B(n_766), .Y(n_765) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_580), .Y(n_776) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI221x1_ASAP7_75t_L g729 ( .A1(n_582), .A2(n_730), .B1(n_732), .B2(n_733), .C(n_735), .Y(n_729) );
AND2x2_ASAP7_75t_L g655 ( .A(n_583), .B(n_611), .Y(n_655) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AND2x2_ASAP7_75t_L g598 ( .A(n_586), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_586), .B(n_588), .Y(n_772) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_592), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_592), .B(n_605), .Y(n_622) );
INVx2_ASAP7_75t_L g629 ( .A(n_592), .Y(n_629) );
INVx1_ASAP7_75t_L g691 ( .A(n_593), .Y(n_691) );
BUFx2_ASAP7_75t_L g711 ( .A(n_594), .Y(n_711) );
NAND2xp33_ASAP7_75t_SL g595 ( .A(n_596), .B(n_598), .Y(n_595) );
OR2x6_ASAP7_75t_L g628 ( .A(n_597), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g757 ( .A(n_597), .B(n_649), .Y(n_757) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_620), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_609), .B1(n_613), .B2(n_618), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
AND2x2_ASAP7_75t_SL g666 ( .A(n_604), .B(n_608), .Y(n_666) );
AND2x4_ASAP7_75t_L g732 ( .A(n_604), .B(n_690), .Y(n_732) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_605), .B(n_606), .Y(n_604) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_605), .Y(n_747) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_608), .B(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_608), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_608), .B(n_639), .Y(n_731) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g752 ( .A(n_610), .B(n_671), .Y(n_752) );
INVx3_ASAP7_75t_L g663 ( .A(n_611), .Y(n_663) );
AND2x2_ASAP7_75t_L g684 ( .A(n_611), .B(n_636), .Y(n_684) );
NAND2x1_ASAP7_75t_SL g755 ( .A(n_611), .B(n_662), .Y(n_755) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B1(n_627), .B2(n_630), .Y(n_620) );
BUFx2_ASAP7_75t_L g676 ( .A(n_622), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_623), .A2(n_714), .B1(n_723), .B2(n_724), .Y(n_722) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g679 ( .A(n_624), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g644 ( .A(n_625), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_629), .B(n_709), .C(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g664 ( .A(n_630), .Y(n_664) );
AOI211x1_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_640), .B(n_642), .C(n_660), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_635), .B(n_723), .Y(n_742) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_636), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g714 ( .A(n_636), .B(n_672), .Y(n_714) );
AND2x2_ASAP7_75t_L g769 ( .A(n_636), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g692 ( .A(n_639), .Y(n_692) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g734 ( .A(n_641), .B(n_679), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_654), .Y(n_642) );
AOI22xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_647), .B1(n_650), .B2(n_652), .Y(n_643) );
BUFx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g707 ( .A(n_646), .B(n_702), .Y(n_707) );
INVx1_ASAP7_75t_SL g749 ( .A(n_646), .Y(n_749) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_SL g717 ( .A(n_649), .B(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g753 ( .A(n_658), .B(n_675), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_665), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_662), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g677 ( .A(n_663), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_667), .Y(n_823) );
NAND3x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_704), .C(n_712), .Y(n_667) );
NAND4xp25_ASAP7_75t_L g778 ( .A(n_668), .B(n_704), .C(n_712), .D(n_779), .Y(n_778) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_682), .Y(n_668) );
OAI222xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_673), .B1(n_676), .B2(n_677), .C1(n_679), .C2(n_681), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g756 ( .A1(n_674), .A2(n_757), .B(n_758), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_675), .B(n_690), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_678), .A2(n_736), .B1(n_738), .B2(n_739), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_693), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_686), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_690), .B(n_692), .Y(n_695) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_700), .B2(n_701), .Y(n_693) );
AND2x4_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
AND2x2_ASAP7_75t_L g701 ( .A(n_697), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_708), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g738 ( .A(n_707), .Y(n_738) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_722), .Y(n_712) );
AOI22xp5_ASAP7_75t_SL g713 ( .A1(n_714), .A2(n_715), .B1(n_717), .B2(n_720), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp33_ASAP7_75t_L g727 ( .A(n_726), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g822 ( .A(n_728), .Y(n_822) );
NAND3x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_740), .C(n_760), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_732), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g766 ( .A(n_737), .Y(n_766) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_750), .Y(n_740) );
AOI21xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_743), .B(n_749), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_756), .Y(n_750) );
INVx2_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_755), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_764), .B2(n_767), .C(n_771), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVxp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B(n_775), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVxp67_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g824 ( .A(n_782), .B(n_825), .C(n_826), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_792), .Y(n_782) );
INVxp33_ASAP7_75t_L g799 ( .A(n_783), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
CKINVDCx8_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_789), .Y(n_796) );
OAI32xp33_ASAP7_75t_L g797 ( .A1(n_789), .A2(n_798), .A3(n_799), .B1(n_800), .B2(n_833), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_792), .Y(n_798) );
INVx1_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2x1_ASAP7_75t_R g801 ( .A(n_795), .B(n_802), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_798), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_802), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_810), .B(n_824), .Y(n_803) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
BUFx3_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_812), .A2(n_813), .B1(n_819), .B2(n_820), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
AND3x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .C(n_823), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
endmodule