module fake_jpeg_29933_n_193 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_19),
.B1(n_21),
.B2(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_59),
.B1(n_63),
.B2(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_0),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_21),
.B1(n_33),
.B2(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_0),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_36),
.A2(n_23),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_16),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_56),
.B(n_44),
.C(n_61),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_55),
.B(n_61),
.C(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_46),
.B1(n_18),
.B2(n_23),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_67),
.B1(n_57),
.B2(n_55),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_17),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_64),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_89),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_29),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_12),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_13),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_11),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_100),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_1),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_9),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_103),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_57),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_89),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_94),
.B(n_84),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_78),
.B1(n_83),
.B2(n_95),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_67),
.B1(n_65),
.B2(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_129),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_118),
.B(n_107),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_78),
.B(n_88),
.C(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_138),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_133),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_78),
.B1(n_99),
.B2(n_79),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_137),
.B1(n_121),
.B2(n_123),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_87),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_141),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_99),
.B1(n_78),
.B2(n_97),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_65),
.B1(n_62),
.B2(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_104),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_3),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_10),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_116),
.B(n_110),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_147),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_104),
.B(n_105),
.C(n_110),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_138),
.B(n_136),
.C(n_132),
.D(n_139),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_118),
.C(n_13),
.Y(n_148)
);

OA21x2_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_152),
.B(n_3),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_125),
.B1(n_137),
.B2(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_119),
.C(n_121),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_133),
.C(n_124),
.Y(n_159)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_162),
.B(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_152),
.B1(n_140),
.B2(n_5),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_164),
.C(n_165),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_125),
.C(n_103),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_65),
.C(n_122),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_122),
.B(n_140),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_147),
.B(n_143),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_173),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_172),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_149),
.B1(n_146),
.B2(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_145),
.B1(n_146),
.B2(n_140),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_160),
.B(n_159),
.C(n_158),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_166),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_SL g175 ( 
.A(n_167),
.B(n_156),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_160),
.B(n_165),
.C(n_164),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_167),
.B1(n_170),
.B2(n_173),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_184),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_185),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_4),
.C(n_7),
.Y(n_185)
);

OAI31xp33_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_176),
.A3(n_179),
.B(n_181),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_187),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_190),
.Y(n_193)
);


endmodule