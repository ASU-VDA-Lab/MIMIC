module fake_jpeg_15567_n_182 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_8),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_21),
.A2(n_31),
.B1(n_17),
.B2(n_32),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_28),
.B(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_56),
.B1(n_26),
.B2(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_18),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_52),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_25),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_61),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_33),
.B1(n_28),
.B2(n_29),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_61),
.B1(n_77),
.B2(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_33),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_19),
.B(n_22),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_76),
.B(n_59),
.C(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_89),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_57),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_12),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_12),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_80),
.B1(n_75),
.B2(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_49),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_104),
.B1(n_93),
.B2(n_107),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_103),
.B(n_84),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_111),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_74),
.B(n_73),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_78),
.B1(n_65),
.B2(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_84),
.Y(n_122)
);

NAND2x1p5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_64),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_88),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_80),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_116),
.C(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_116),
.B1(n_97),
.B2(n_92),
.Y(n_138)
);

OAI21x1_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_90),
.B(n_97),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_117),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_87),
.B1(n_61),
.B2(n_67),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_125),
.B(n_128),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_98),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_94),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_137),
.B1(n_139),
.B2(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_94),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_95),
.B1(n_96),
.B2(n_137),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_140),
.B1(n_122),
.B2(n_130),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_99),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_106),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_149),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_144),
.B1(n_153),
.B2(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_127),
.B1(n_125),
.B2(n_119),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_150),
.B1(n_152),
.B2(n_157),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_129),
.C(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_128),
.B1(n_131),
.B2(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_145),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_121),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_132),
.C(n_133),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_155),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_127),
.B1(n_124),
.B2(n_136),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_147),
.B(n_151),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_143),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_157),
.B(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_158),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_164),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_172),
.B1(n_173),
.B2(n_171),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.C(n_161),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_161),
.C(n_167),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_178),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_179),
.B(n_171),
.Y(n_182)
);


endmodule