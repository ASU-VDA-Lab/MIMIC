module real_jpeg_16667_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_493;
wire n_93;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_1),
.B(n_132),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_1),
.B(n_288),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_1),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_1),
.B(n_437),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_SL g474 ( 
.A(n_1),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_1),
.B(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_1),
.B(n_507),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_2),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_2),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_2),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_2),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_2),
.B(n_135),
.Y(n_134)
);

NAND2x1p5_ASAP7_75t_L g222 ( 
.A(n_2),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_3),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g478 ( 
.A(n_3),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_4),
.Y(n_349)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_4),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_5),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_5),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_5),
.B(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_5),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_5),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_5),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_7),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_7),
.Y(n_461)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_8),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_8),
.Y(n_352)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_8),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_9),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_9),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_9),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_9),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_9),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_9),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_9),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_9),
.B(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_10),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_10),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_10),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_10),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_10),
.B(n_432),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_10),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_10),
.B(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_10),
.B(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

BUFx8_ASAP7_75t_L g214 ( 
.A(n_11),
.Y(n_214)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_12),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_12),
.B(n_55),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_12),
.A2(n_17),
.B1(n_309),
.B2(n_313),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_12),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_12),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_12),
.B(n_493),
.Y(n_492)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_13),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_13),
.Y(n_290)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_14),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_14),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_14),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_14),
.B(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g212 ( 
.A(n_16),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_16),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_16),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_17),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_17),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_17),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_17),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_17),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_131),
.Y(n_236)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_256),
.B(n_529),
.C(n_536),
.D(n_538),
.Y(n_21)
);

NOR3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_226),
.C(n_244),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_179),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21x1_ASAP7_75t_SL g531 ( 
.A1(n_25),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_147),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_26),
.B(n_147),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_111),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_27),
.B(n_112),
.C(n_124),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_77),
.C(n_93),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_28),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.C(n_62),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_29),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_40),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_38),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_31),
.B(n_39),
.C(n_40),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_31),
.B(n_297),
.C(n_298),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_31),
.A2(n_38),
.B1(n_297),
.B2(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_33),
.Y(n_444)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_34),
.B(n_96),
.C(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_34),
.A2(n_39),
.B1(n_96),
.B2(n_97),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_34),
.B(n_215),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_SL g408 ( 
.A(n_34),
.B(n_306),
.Y(n_408)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_36),
.Y(n_163)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_36),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_37),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_38),
.B(n_115),
.C(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_41),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_41),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_46),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_46),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_47),
.B(n_62),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.C(n_57),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_165)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_57),
.A2(n_58),
.B1(n_115),
.B2(n_117),
.Y(n_318)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_58),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_58),
.B(n_115),
.C(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_61),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_71),
.C(n_75),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_63),
.B(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_63),
.B(n_138),
.C(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_71),
.A2(n_76),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_76),
.B(n_138),
.C(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_77),
.B(n_93),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_87),
.B2(n_92),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_82),
.C(n_87),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_81),
.B(n_168),
.C(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_81),
.B(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_86),
.Y(n_315)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_87),
.A2(n_92),
.B1(n_250),
.B2(n_253),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_87),
.B(n_251),
.C(n_252),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_107),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_94),
.A2(n_95),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_158),
.C(n_161),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_96),
.A2(n_97),
.B1(n_161),
.B2(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_96),
.B(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_97),
.B(n_416),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_98),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_99),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_99),
.Y(n_251)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_103),
.A2(n_247),
.B(n_537),
.Y(n_538)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_104),
.B(n_107),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_107),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_107),
.A2(n_143),
.B1(n_173),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_110),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_124),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_123),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_117),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_117),
.B(n_134),
.C(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_123),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_139),
.B2(n_140),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_127),
.B(n_128),
.C(n_139),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_134),
.A2(n_138),
.B1(n_221),
.B2(n_222),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_134),
.A2(n_138),
.B1(n_195),
.B2(n_266),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_141),
.B(n_143),
.C(n_145),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_167),
.C(n_173),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_152),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_150),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_166),
.C(n_176),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_154),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_164),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_155),
.B(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_157),
.B(n_164),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_159),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_159),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_161),
.A2(n_162),
.B1(n_293),
.B2(n_294),
.Y(n_344)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_162),
.B(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_176),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_193),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_170),
.Y(n_299)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

OR2x2_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_180),
.B(n_182),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_189),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_183),
.B(n_187),
.Y(n_393)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_189),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_202),
.C(n_206),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_190),
.A2(n_191),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_199),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g378 ( 
.A(n_192),
.B(n_379),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_194),
.B(n_200),
.Y(n_379)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.C(n_221),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_208),
.A2(n_209),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_210),
.A2(n_215),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_210),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_213),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_215),
.Y(n_306)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_217),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

BUFx2_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g530 ( 
.A1(n_227),
.A2(n_245),
.B(n_531),
.C(n_534),
.D(n_535),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_243),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_228),
.B(n_243),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_231),
.C(n_242),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_241),
.B2(n_242),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_237),
.C(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_255),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_246),
.B(n_255),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_246),
.Y(n_540)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.CI(n_254),
.CON(n_246),
.SN(n_246)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_248),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

NAND2x1_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_523),
.Y(n_256)
);

NAND4xp25_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_380),
.C(n_394),
.D(n_399),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_357),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_333),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_260),
.B(n_333),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_300),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_261),
.B(n_301),
.C(n_316),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_278),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_263),
.Y(n_361)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_267),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_276),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_268)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_269),
.A2(n_272),
.B(n_276),
.C(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_271),
.B(n_275),
.Y(n_374)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_274),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_278),
.B(n_361),
.C(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_291),
.C(n_296),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_279),
.B(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_283),
.C(n_287),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_291),
.A2(n_292),
.B1(n_296),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g516 ( 
.A(n_295),
.Y(n_516)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_297),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_316),
.Y(n_300)
);

XOR2x2_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_303),
.B(n_367),
.C(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_320),
.B(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_SL g494 ( 
.A(n_311),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.C(n_326),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_319),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_326),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.C(n_331),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_406)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.C(n_340),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_334),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_336),
.A2(n_337),
.B1(n_340),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.C(n_345),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_341),
.B(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_344),
.B(n_345),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_350),
.C(n_353),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_346),
.B(n_353),
.Y(n_446)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_350),
.B(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

OAI21x1_ASAP7_75t_SL g524 ( 
.A1(n_357),
.A2(n_525),
.B(n_526),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_358),
.B(n_359),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_364),
.C(n_378),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_377),
.B2(n_378),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_373),
.B1(n_375),
.B2(n_376),
.Y(n_369)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_370),
.Y(n_375)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_373),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_388),
.C(n_389),
.Y(n_387)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

A2O1A1O1Ixp25_ASAP7_75t_L g523 ( 
.A1(n_380),
.A2(n_394),
.B(n_524),
.C(n_527),
.D(n_528),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_392),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_381),
.B(n_392),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_386),
.C(n_390),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_382),
.A2(n_383),
.B1(n_390),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_384),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_395),
.B(n_396),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_424),
.B(n_522),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_421),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_401),
.B(n_421),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_405),
.C(n_407),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_402),
.A2(n_403),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_405),
.B(n_407),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.C(n_415),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_408),
.A2(n_409),
.B1(n_410),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_408),
.Y(n_429)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_415),
.B(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

AOI21x1_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_450),
.B(n_521),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_447),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_426),
.B(n_447),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.C(n_445),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_445),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_436),
.C(n_442),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_455),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_435),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_442),
.Y(n_455)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_469),
.B(n_520),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_467),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_452),
.B(n_467),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_456),
.C(n_465),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_453),
.A2(n_454),
.B1(n_480),
.B2(n_482),
.Y(n_479)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_456),
.A2(n_465),
.B1(n_466),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_456),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_462),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_457),
.A2(n_458),
.B1(n_462),
.B2(n_463),
.Y(n_472)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_483),
.B(n_519),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_479),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_471),
.B(n_479),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.C(n_477),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_496),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_477),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_480),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_484),
.A2(n_498),
.B(n_518),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_495),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_485),
.B(n_495),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_492),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_492),
.Y(n_504)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_505),
.B(n_517),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_504),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_500),
.B(n_504),
.Y(n_517)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_513),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_537),
.Y(n_536)
);


endmodule