module fake_jpeg_12462_n_570 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_570);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_570;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_11),
.B(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_7),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_61),
.B(n_77),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_62),
.Y(n_183)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_78),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_84),
.Y(n_187)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_87),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_32),
.B(n_7),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_90),
.B(n_97),
.Y(n_157)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_22),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_32),
.B(n_8),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_27),
.B(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_124),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_8),
.B(n_17),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_33),
.B(n_6),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_33),
.B(n_18),
.Y(n_124)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_19),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_54),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_132),
.B(n_135),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_66),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_77),
.B(n_54),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_149),
.B(n_152),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_80),
.A2(n_24),
.B1(n_58),
.B2(n_23),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_150),
.A2(n_186),
.B1(n_198),
.B2(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_46),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_46),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_96),
.B(n_45),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_62),
.A2(n_24),
.B1(n_35),
.B2(n_59),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_178),
.A2(n_58),
.B1(n_35),
.B2(n_111),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_98),
.B(n_45),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_191),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_103),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_199),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_60),
.A2(n_24),
.B1(n_52),
.B2(n_59),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_70),
.A2(n_52),
.B1(n_57),
.B2(n_28),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_190),
.B1(n_202),
.B2(n_20),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_73),
.A2(n_57),
.B1(n_51),
.B2(n_50),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_105),
.B(n_40),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_40),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_195),
.B(n_206),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_71),
.A2(n_39),
.B1(n_51),
.B2(n_50),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_114),
.B(n_49),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_74),
.A2(n_35),
.B(n_58),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_20),
.C(n_1),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_85),
.A2(n_58),
.B1(n_35),
.B2(n_39),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_75),
.A2(n_38),
.B1(n_37),
.B2(n_49),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_76),
.A2(n_58),
.B1(n_35),
.B2(n_37),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_122),
.B(n_38),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_208),
.Y(n_302)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_210),
.B(n_229),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_211),
.Y(n_324)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_212),
.Y(n_325)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_213),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_215),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_110),
.B1(n_102),
.B2(n_95),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_216),
.Y(n_306)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_217),
.Y(n_316)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_219),
.Y(n_301)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_224),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_146),
.B(n_0),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_225),
.B(n_238),
.Y(n_314)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_154),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_226),
.B(n_234),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_227),
.Y(n_328)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_162),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_127),
.A2(n_93),
.B1(n_88),
.B2(n_84),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_230),
.A2(n_236),
.B1(n_256),
.B2(n_258),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_186),
.A2(n_79),
.B1(n_78),
.B2(n_20),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_231),
.A2(n_232),
.B1(n_261),
.B2(n_145),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_20),
.B1(n_9),
.B2(n_2),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_233),
.A2(n_247),
.B(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_144),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_20),
.B1(n_9),
.B2(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_146),
.A2(n_6),
.B1(n_17),
.B2(n_3),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_241),
.A2(n_187),
.B(n_197),
.Y(n_297)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

BUFx2_ASAP7_75t_SL g243 ( 
.A(n_151),
.Y(n_243)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_246),
.A2(n_265),
.B1(n_272),
.B2(n_219),
.Y(n_299)
);

NAND2x1_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_4),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_248),
.B(n_249),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_198),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_183),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_251),
.B(n_259),
.Y(n_290)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_143),
.Y(n_253)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_131),
.Y(n_254)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_190),
.A2(n_4),
.B1(n_5),
.B2(n_14),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_266),
.B1(n_171),
.B2(n_175),
.Y(n_288)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_134),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_128),
.A2(n_4),
.B(n_5),
.C(n_15),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_257),
.A2(n_276),
.B(n_269),
.C(n_253),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_167),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_157),
.B(n_5),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_263),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_201),
.A2(n_1),
.B1(n_15),
.B2(n_16),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_161),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_262),
.B(n_267),
.Y(n_292)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_126),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_172),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_264),
.B(n_258),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_189),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_130),
.B(n_196),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_177),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_268),
.B(n_270),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g269 ( 
.A1(n_126),
.A2(n_207),
.B1(n_171),
.B2(n_137),
.Y(n_269)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_269),
.A2(n_277),
.B1(n_263),
.B2(n_242),
.Y(n_320)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_145),
.A2(n_142),
.B1(n_140),
.B2(n_203),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_204),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_159),
.B(n_165),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_139),
.B(n_141),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_276),
.B(n_275),
.Y(n_311)
);

AO22x2_ASAP7_75t_SL g277 ( 
.A1(n_168),
.A2(n_153),
.B1(n_175),
.B2(n_137),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_233),
.A2(n_168),
.B1(n_153),
.B2(n_207),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_279),
.A2(n_283),
.B1(n_288),
.B2(n_289),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_248),
.A2(n_238),
.B1(n_215),
.B2(n_277),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_129),
.B1(n_136),
.B2(n_156),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_223),
.A2(n_136),
.B1(n_156),
.B2(n_192),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_291),
.A2(n_304),
.B1(n_326),
.B2(n_332),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_311),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_231),
.A2(n_197),
.B1(n_187),
.B2(n_148),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_294),
.A2(n_299),
.B1(n_301),
.B2(n_322),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_299),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_266),
.A2(n_239),
.B1(n_241),
.B2(n_273),
.Y(n_304)
);

AOI32xp33_ASAP7_75t_L g310 ( 
.A1(n_245),
.A2(n_225),
.A3(n_240),
.B1(n_247),
.B2(n_214),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_310),
.B(n_290),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_225),
.A2(n_235),
.B(n_261),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_232),
.A2(n_257),
.B(n_275),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_320),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_331),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_269),
.A2(n_209),
.B1(n_213),
.B2(n_228),
.Y(n_326)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_276),
.A2(n_264),
.B(n_221),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_269),
.A2(n_252),
.B1(n_254),
.B2(n_208),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_303),
.A2(n_211),
.B1(n_265),
.B2(n_272),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_335),
.A2(n_340),
.B1(n_343),
.B2(n_345),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_296),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_354),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_220),
.C(n_224),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_352),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_283),
.A2(n_250),
.B1(n_256),
.B2(n_260),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_339),
.A2(n_325),
.B(n_348),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_303),
.A2(n_218),
.B1(n_222),
.B2(n_327),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_303),
.A2(n_327),
.B1(n_293),
.B2(n_308),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_310),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_367),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_318),
.A2(n_313),
.B1(n_306),
.B2(n_321),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_346),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_355),
.B1(n_323),
.B2(n_312),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_291),
.A2(n_279),
.B1(n_289),
.B2(n_326),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_350),
.A2(n_349),
.B1(n_339),
.B2(n_370),
.Y(n_406)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_286),
.C(n_311),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_285),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_320),
.A2(n_297),
.B1(n_304),
.B2(n_280),
.Y(n_355)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_292),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_320),
.A2(n_288),
.B1(n_280),
.B2(n_292),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_357),
.A2(n_365),
.B1(n_369),
.B2(n_374),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_285),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_360),
.Y(n_381)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_329),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_316),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_366),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_364),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_290),
.B1(n_301),
.B2(n_332),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_316),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_298),
.B(n_309),
.C(n_331),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_371),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_320),
.A2(n_317),
.B1(n_328),
.B2(n_282),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_325),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_298),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_372),
.B(n_284),
.Y(n_389)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_278),
.Y(n_373)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_282),
.A2(n_319),
.B1(n_324),
.B2(n_309),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_342),
.A2(n_319),
.B1(n_287),
.B2(n_324),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_375),
.A2(n_394),
.B1(n_401),
.B2(n_406),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_360),
.B(n_278),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_398),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_323),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_383),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_389),
.B(n_358),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_390),
.A2(n_396),
.B1(n_397),
.B2(n_361),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_342),
.A2(n_287),
.B1(n_284),
.B2(n_330),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_362),
.A2(n_312),
.B1(n_305),
.B2(n_281),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_335),
.A2(n_330),
.B1(n_300),
.B2(n_281),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_399),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_368),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_405),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_349),
.A2(n_300),
.B1(n_315),
.B2(n_302),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_353),
.A2(n_305),
.B(n_315),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_403),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_336),
.B(n_354),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_334),
.B(n_333),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_407),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_334),
.Y(n_409)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_409),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_387),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_388),
.A2(n_350),
.B1(n_355),
.B2(n_334),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_412),
.A2(n_419),
.B1(n_426),
.B2(n_438),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_344),
.C(n_352),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_415),
.C(n_421),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_380),
.B(n_344),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_388),
.A2(n_334),
.B1(n_357),
.B2(n_333),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_338),
.C(n_345),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_406),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_343),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_431),
.C(n_437),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_382),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_434),
.Y(n_442)
);

OAI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_408),
.A2(n_365),
.B1(n_369),
.B2(n_340),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_429),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_SL g430 ( 
.A1(n_378),
.A2(n_333),
.B(n_367),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_430),
.A2(n_383),
.B1(n_409),
.B2(n_407),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_380),
.B(n_333),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_379),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_432),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_393),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_378),
.Y(n_435)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_435),
.Y(n_447)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_436),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_392),
.B(n_363),
.C(n_337),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_386),
.A2(n_347),
.B1(n_346),
.B2(n_341),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_439),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_457),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_445),
.A2(n_412),
.B1(n_419),
.B2(n_417),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_446),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_381),
.B(n_389),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_448),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_429),
.A2(n_391),
.B1(n_400),
.B2(n_409),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_450),
.A2(n_466),
.B1(n_394),
.B2(n_401),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_415),
.B(n_381),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_451),
.B(n_452),
.Y(n_489)
);

XNOR2x1_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_383),
.Y(n_452)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_454),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_433),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_440),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_398),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_414),
.A2(n_391),
.B1(n_405),
.B2(n_386),
.Y(n_460)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_460),
.Y(n_475)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_416),
.Y(n_461)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_413),
.B(n_407),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_465),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_377),
.C(n_403),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_410),
.C(n_440),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_404),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_414),
.A2(n_439),
.B1(n_436),
.B2(n_425),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_467),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_420),
.B(n_384),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_416),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_464),
.A2(n_410),
.B1(n_427),
.B2(n_418),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_469),
.A2(n_476),
.B1(n_450),
.B2(n_445),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_418),
.Y(n_471)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_434),
.Y(n_474)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_464),
.A2(n_441),
.B1(n_453),
.B2(n_449),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_484),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_458),
.Y(n_505)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_481),
.Y(n_496)
);

AOI21xp33_ASAP7_75t_L g483 ( 
.A1(n_465),
.A2(n_427),
.B(n_422),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_483),
.B(n_487),
.Y(n_494)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_442),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_485),
.A2(n_459),
.B(n_456),
.Y(n_500)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_447),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_399),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_445),
.A2(n_417),
.B1(n_422),
.B2(n_375),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_488),
.A2(n_490),
.B1(n_454),
.B2(n_376),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_371),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_491),
.B(n_463),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_495),
.Y(n_517)
);

XOR2x1_ASAP7_75t_SL g497 ( 
.A(n_489),
.B(n_444),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_500),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_498),
.A2(n_511),
.B1(n_485),
.B2(n_488),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_471),
.B(n_459),
.CI(n_452),
.CON(n_502),
.SN(n_502)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_479),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_503),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_458),
.C(n_462),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_505),
.C(n_507),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_482),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_474),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_451),
.C(n_456),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_443),
.C(n_387),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_509),
.C(n_486),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_432),
.C(n_393),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_510),
.A2(n_469),
.B1(n_475),
.B2(n_476),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_475),
.A2(n_402),
.B1(n_376),
.B2(n_374),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_526),
.Y(n_539)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_503),
.Y(n_515)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_515),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_516),
.A2(n_510),
.B1(n_496),
.B2(n_509),
.Y(n_534)
);

OAI22x1_ASAP7_75t_L g530 ( 
.A1(n_518),
.A2(n_498),
.B1(n_490),
.B2(n_501),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_493),
.B(n_470),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_525),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_523),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_499),
.Y(n_521)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_521),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_484),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_494),
.B(n_487),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_508),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_499),
.A2(n_470),
.B(n_481),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_477),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_529),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_519),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_518),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_531),
.B(n_532),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_526),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_534),
.A2(n_500),
.B1(n_511),
.B2(n_513),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_477),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_537),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_492),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_535),
.A2(n_516),
.B(n_515),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_541),
.A2(n_548),
.B(n_539),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_520),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_542),
.B(n_544),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_543),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_528),
.A2(n_496),
.B1(n_513),
.B2(n_523),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_547),
.Y(n_555)
);

FAx1_ASAP7_75t_SL g547 ( 
.A(n_535),
.B(n_497),
.CI(n_502),
.CON(n_547),
.SN(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_539),
.A2(n_522),
.B(n_505),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_550),
.B(n_541),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_549),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_551),
.B(n_553),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_546),
.A2(n_534),
.B(n_533),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_552),
.A2(n_540),
.B(n_547),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_522),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_558),
.B(n_547),
.C(n_530),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_554),
.B(n_544),
.C(n_543),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_560),
.B(n_561),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_555),
.A2(n_556),
.B(n_552),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_562),
.B(n_564),
.C(n_506),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_557),
.A2(n_559),
.B(n_504),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_565),
.B(n_566),
.C(n_472),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_472),
.C(n_492),
.Y(n_566)
);

A2O1A1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_567),
.A2(n_502),
.B(n_376),
.C(n_366),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_402),
.C(n_351),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_364),
.C(n_557),
.Y(n_570)
);


endmodule