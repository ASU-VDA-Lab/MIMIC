module fake_jpeg_12837_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_5),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

BUFx12f_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_82),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_24),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_65),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_67),
.Y(n_147)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_29),
.B(n_0),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_25),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_83),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_34),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_30),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_45),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

BUFx4f_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_31),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_45),
.B1(n_38),
.B2(n_32),
.Y(n_144)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_32),
.Y(n_141)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_31),
.B1(n_26),
.B2(n_37),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_117),
.A2(n_129),
.B1(n_144),
.B2(n_155),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_120),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_83),
.B1(n_54),
.B2(n_60),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_121),
.A2(n_77),
.B1(n_104),
.B2(n_106),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_126),
.B(n_87),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_68),
.A2(n_45),
.B1(n_51),
.B2(n_50),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_128),
.A2(n_156),
.B(n_171),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_53),
.A2(n_26),
.B1(n_37),
.B2(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_65),
.B(n_38),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_141),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_78),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_52),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_55),
.B(n_52),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_160),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_62),
.A2(n_37),
.B1(n_40),
.B2(n_46),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_72),
.A2(n_51),
.B1(n_50),
.B2(n_46),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_81),
.B(n_39),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_34),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_93),
.A2(n_50),
.B1(n_51),
.B2(n_34),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_116),
.B(n_110),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_173),
.B(n_176),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_109),
.B(n_22),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_121),
.A2(n_64),
.B1(n_75),
.B2(n_97),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_177),
.A2(n_196),
.B1(n_42),
.B2(n_2),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_113),
.A2(n_67),
.B(n_39),
.C(n_20),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_178),
.A2(n_42),
.B(n_124),
.C(n_3),
.Y(n_262)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_179),
.Y(n_271)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g258 ( 
.A(n_182),
.Y(n_258)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_36),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_189),
.Y(n_264)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_191),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_220),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_118),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_203),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_199),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_132),
.A2(n_91),
.B1(n_80),
.B2(n_86),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_206),
.A2(n_210),
.B1(n_221),
.B2(n_164),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_138),
.B(n_36),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_136),
.Y(n_208)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_208),
.Y(n_285)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_136),
.A2(n_85),
.B1(n_35),
.B2(n_28),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_212),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_213),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_114),
.Y(n_256)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_156),
.A2(n_171),
.B1(n_128),
.B2(n_135),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_216),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_288)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_112),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_162),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_218),
.B(n_225),
.Y(n_283)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_229),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_137),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_135),
.A2(n_35),
.B1(n_28),
.B2(n_22),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_222),
.B(n_66),
.Y(n_265)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_139),
.B(n_0),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_233),
.Y(n_260)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_230),
.Y(n_279)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_134),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_234),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_139),
.B(n_158),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_153),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_161),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_183),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_239),
.B(n_252),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_173),
.B(n_145),
.CI(n_152),
.CON(n_242),
.SN(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_242),
.A2(n_225),
.B(n_215),
.C(n_218),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_223),
.A2(n_114),
.B1(n_130),
.B2(n_133),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_185),
.A2(n_133),
.B1(n_164),
.B2(n_142),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_247),
.A2(n_243),
.B1(n_258),
.B2(n_193),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_154),
.B(n_130),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_255),
.A2(n_11),
.B(n_14),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_256),
.B(n_261),
.Y(n_335)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_186),
.B(n_124),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_262),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_265),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_176),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_280),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_177),
.A2(n_124),
.B1(n_153),
.B2(n_134),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_275),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_142),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_212),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_192),
.B(n_87),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_66),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_211),
.C(n_179),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_190),
.B1(n_178),
.B2(n_208),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_210),
.B1(n_231),
.B2(n_182),
.Y(n_300)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_253),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_292),
.B(n_306),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_254),
.B(n_204),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_293),
.B(n_302),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_255),
.A2(n_185),
.B1(n_204),
.B2(n_224),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_295),
.A2(n_297),
.B1(n_300),
.B2(n_301),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_224),
.B1(n_206),
.B2(n_228),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_299),
.A2(n_320),
.B1(n_334),
.B2(n_269),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_214),
.B1(n_205),
.B2(n_229),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_256),
.B(n_180),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_304),
.A2(n_330),
.B1(n_339),
.B2(n_269),
.Y(n_341)
);

AO21x2_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_201),
.B(n_174),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_309),
.B1(n_258),
.B2(n_278),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_283),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_332),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_250),
.B(n_175),
.Y(n_308)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_313),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_247),
.A2(n_188),
.B1(n_181),
.B2(n_219),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_260),
.A2(n_197),
.B1(n_200),
.B2(n_232),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_310),
.A2(n_319),
.B1(n_327),
.B2(n_333),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_312),
.A2(n_315),
.B(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_SL g315 ( 
.A1(n_262),
.A2(n_230),
.B(n_213),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_317),
.B(n_322),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_260),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_246),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_284),
.B(n_250),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_261),
.B(n_242),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_323),
.B(n_326),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_324),
.A2(n_338),
.B1(n_238),
.B2(n_282),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_261),
.B(n_8),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_288),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_242),
.B(n_17),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_290),
.Y(n_372)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_264),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_236),
.B(n_238),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_251),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_263),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_264),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_237),
.A2(n_16),
.B1(n_263),
.B2(n_283),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_337),
.Y(n_380)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_272),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_237),
.A2(n_258),
.B1(n_268),
.B2(n_271),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_357),
.B1(n_359),
.B2(n_329),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_341),
.A2(n_345),
.B(n_369),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_335),
.C(n_302),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_355),
.C(n_364),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_346),
.A2(n_348),
.B1(n_349),
.B2(n_359),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_316),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_356),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_311),
.A2(n_323),
.B1(n_328),
.B2(n_305),
.Y(n_348)
);

OAI22x1_ASAP7_75t_SL g349 ( 
.A1(n_305),
.A2(n_245),
.B1(n_271),
.B2(n_282),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_322),
.B(n_268),
.C(n_257),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_317),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_278),
.B1(n_241),
.B2(n_272),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_305),
.A2(n_241),
.B1(n_285),
.B2(n_245),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_295),
.A2(n_285),
.B1(n_248),
.B2(n_287),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_360),
.A2(n_362),
.B1(n_371),
.B2(n_370),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_305),
.A2(n_294),
.B1(n_299),
.B2(n_293),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_373),
.B1(n_374),
.B2(n_377),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_297),
.A2(n_248),
.B1(n_287),
.B2(n_240),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_363),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_286),
.C(n_259),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_296),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_365),
.B(n_372),
.Y(n_404)
);

AO22x1_ASAP7_75t_L g369 ( 
.A1(n_312),
.A2(n_281),
.B1(n_249),
.B2(n_259),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_301),
.A2(n_240),
.B1(n_281),
.B2(n_279),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_305),
.A2(n_249),
.B1(n_290),
.B2(n_294),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_296),
.A2(n_309),
.B1(n_307),
.B2(n_306),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_302),
.C(n_313),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_336),
.C(n_314),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_292),
.A2(n_300),
.B1(n_302),
.B2(n_298),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_310),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_350),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_380),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_335),
.B(n_331),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_382),
.A2(n_390),
.B(n_410),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_350),
.A2(n_291),
.B1(n_303),
.B2(n_332),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_379),
.B1(n_349),
.B2(n_369),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_342),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_384),
.B(n_387),
.C(n_393),
.Y(n_435)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_385),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_326),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_374),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_391),
.Y(n_425)
);

AOI22x1_ASAP7_75t_L g390 ( 
.A1(n_361),
.A2(n_318),
.B1(n_327),
.B2(n_319),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_392),
.Y(n_434)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_399),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_308),
.C(n_321),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_405),
.C(n_412),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_344),
.A2(n_333),
.B(n_338),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_398),
.A2(n_354),
.B(n_370),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_375),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_346),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_402),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_406),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_325),
.C(n_368),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_408),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_356),
.B(n_365),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_347),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_411),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_369),
.A2(n_378),
.B(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_368),
.C(n_355),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_343),
.B(n_366),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_414),
.B(n_366),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_377),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_348),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_416),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_426),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_421),
.A2(n_422),
.B1(n_438),
.B2(n_423),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_402),
.B1(n_415),
.B2(n_401),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_423),
.A2(n_438),
.B1(n_388),
.B2(n_385),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_417),
.A2(n_341),
.B1(n_358),
.B2(n_343),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_424),
.A2(n_433),
.B1(n_440),
.B2(n_442),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_372),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_362),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_428),
.B(n_429),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_354),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_413),
.B(n_345),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_436),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_395),
.A2(n_410),
.B(n_417),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_383),
.A2(n_358),
.B1(n_381),
.B2(n_371),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_387),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_446),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_400),
.A2(n_408),
.B1(n_398),
.B2(n_382),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_400),
.A2(n_381),
.B1(n_405),
.B2(n_395),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_404),
.Y(n_445)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_445),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_386),
.B(n_393),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_396),
.B(n_412),
.C(n_414),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_394),
.C(n_403),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_390),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_411),
.Y(n_465)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_441),
.Y(n_449)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_441),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_450),
.B(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_455),
.A2(n_470),
.B1(n_434),
.B2(n_419),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_459),
.Y(n_480)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_390),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_406),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_465),
.Y(n_479)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_420),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_466),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_392),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_463),
.Y(n_478)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_388),
.C(n_435),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_468),
.A2(n_418),
.B1(n_448),
.B2(n_430),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_436),
.A2(n_437),
.B1(n_430),
.B2(n_422),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_435),
.C(n_447),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_472),
.Y(n_482)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_432),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_424),
.A2(n_425),
.B1(n_440),
.B2(n_442),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_473),
.A2(n_464),
.B1(n_449),
.B2(n_454),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_431),
.B(n_443),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_474),
.B(n_453),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_477),
.A2(n_484),
.B1(n_492),
.B2(n_457),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_464),
.A2(n_425),
.B1(n_418),
.B2(n_433),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_481),
.A2(n_491),
.B1(n_451),
.B2(n_452),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_483),
.B(n_471),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_439),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_485),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_434),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_495),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_455),
.A2(n_470),
.B1(n_461),
.B2(n_462),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_469),
.A2(n_459),
.B(n_465),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_493),
.A2(n_484),
.B(n_476),
.Y(n_511)
);

XOR2x1_ASAP7_75t_SL g494 ( 
.A(n_463),
.B(n_458),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_466),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_452),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_482),
.B(n_456),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g519 ( 
.A(n_496),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_511),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_500),
.B(n_504),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_501),
.B(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_503),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_492),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_476),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_505),
.A2(n_475),
.B1(n_490),
.B2(n_478),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_495),
.C(n_488),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_479),
.C(n_481),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_480),
.B(n_489),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_507),
.Y(n_513)
);

INVx6_ASAP7_75t_L g508 ( 
.A(n_494),
.Y(n_508)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_508),
.Y(n_521)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_509),
.Y(n_522)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_477),
.A2(n_493),
.B(n_475),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_512),
.A2(n_490),
.B(n_479),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_526),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_499),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_517),
.B(n_499),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_497),
.A2(n_508),
.B1(n_505),
.B2(n_503),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_524),
.B(n_521),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_512),
.A2(n_502),
.B(n_498),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_509),
.B1(n_510),
.B2(n_501),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_528),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_518),
.B(n_506),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_511),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_529),
.B(n_530),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_535),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_523),
.C(n_514),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_SL g541 ( 
.A(n_532),
.B(n_534),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_513),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_533),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_540),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_532),
.A2(n_516),
.B(n_514),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_534),
.C(n_530),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_539),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g543 ( 
.A(n_537),
.B(n_521),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_542),
.C(n_544),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_SL g547 ( 
.A(n_545),
.B(n_546),
.C(n_541),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_547),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_520),
.C(n_522),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_520),
.B(n_522),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_525),
.C(n_549),
.Y(n_551)
);


endmodule