module real_aes_13318_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_102;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx2_ASAP7_75t_SL g133 ( .A(n_0), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_1), .Y(n_286) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_2), .A2(n_45), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g139 ( .A(n_2), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_3), .B(n_129), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_4), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g717 ( .A(n_5), .Y(n_717) );
INVx1_ASAP7_75t_L g555 ( .A(n_6), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_6), .A2(n_32), .B1(n_659), .B2(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g645 ( .A(n_7), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_7), .A2(n_37), .B1(n_659), .B2(n_661), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_8), .A2(n_26), .B1(n_527), .B2(n_535), .Y(n_526) );
INVx1_ASAP7_75t_L g594 ( .A(n_8), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_9), .Y(n_649) );
AND2x2_ASAP7_75t_L g225 ( .A(n_10), .B(n_146), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_11), .B(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g534 ( .A(n_12), .Y(n_534) );
INVx3_ASAP7_75t_L g579 ( .A(n_13), .Y(n_579) );
INVx1_ASAP7_75t_L g538 ( .A(n_14), .Y(n_538) );
INVx2_ASAP7_75t_L g552 ( .A(n_14), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_15), .B(n_237), .Y(n_259) );
INVx1_ASAP7_75t_L g96 ( .A(n_16), .Y(n_96) );
BUFx3_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_17), .B(n_145), .Y(n_269) );
BUFx10_ASAP7_75t_L g702 ( .A(n_18), .Y(n_702) );
XNOR2xp5_ASAP7_75t_L g522 ( .A(n_19), .B(n_523), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_20), .Y(n_250) );
NAND3xp33_ASAP7_75t_L g203 ( .A(n_21), .B(n_201), .C(n_204), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_22), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_23), .B(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_24), .Y(n_620) );
INVx1_ASAP7_75t_L g670 ( .A(n_24), .Y(n_670) );
OAI33xp33_ASAP7_75t_L g595 ( .A1(n_25), .A2(n_59), .A3(n_596), .B1(n_599), .B2(n_600), .B3(n_602), .Y(n_595) );
INVx1_ASAP7_75t_L g640 ( .A(n_25), .Y(n_640) );
INVx1_ASAP7_75t_L g657 ( .A(n_26), .Y(n_657) );
INVx1_ASAP7_75t_L g87 ( .A(n_27), .Y(n_87) );
INVx2_ASAP7_75t_L g586 ( .A(n_28), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_29), .B(n_115), .Y(n_114) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_30), .A2(n_612), .B(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g646 ( .A(n_30), .Y(n_646) );
INVx1_ASAP7_75t_L g559 ( .A(n_31), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_31), .A2(n_582), .B(n_590), .Y(n_581) );
OAI21xp5_ASAP7_75t_SL g539 ( .A1(n_32), .A2(n_540), .B(n_545), .Y(n_539) );
INVx1_ASAP7_75t_L g642 ( .A(n_33), .Y(n_642) );
AOI21xp5_ASAP7_75t_SL g673 ( .A1(n_33), .A2(n_674), .B(n_675), .Y(n_673) );
INVx2_ASAP7_75t_L g589 ( .A(n_34), .Y(n_589) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_34), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_34), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_35), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_36), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g629 ( .A(n_37), .Y(n_629) );
AND2x4_ASAP7_75t_L g86 ( .A(n_38), .B(n_87), .Y(n_86) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_38), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_39), .B(n_145), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_40), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_41), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g532 ( .A(n_42), .Y(n_532) );
INVx1_ASAP7_75t_L g544 ( .A(n_42), .Y(n_544) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_43), .Y(n_723) );
INVx1_ASAP7_75t_L g719 ( .A(n_44), .Y(n_719) );
INVx1_ASAP7_75t_L g138 ( .A(n_45), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_46), .Y(n_222) );
INVx1_ASAP7_75t_L g564 ( .A(n_47), .Y(n_564) );
AOI21xp33_ASAP7_75t_L g663 ( .A1(n_47), .A2(n_664), .B(n_668), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g127 ( .A1(n_48), .A2(n_128), .B(n_130), .C(n_134), .Y(n_127) );
INVx1_ASAP7_75t_L g126 ( .A(n_49), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_50), .B(n_145), .Y(n_292) );
INVx3_ASAP7_75t_L g247 ( .A(n_51), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_52), .B(n_151), .Y(n_158) );
INVx1_ASAP7_75t_L g262 ( .A(n_53), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_54), .B(n_196), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_55), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_56), .B(n_204), .Y(n_283) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_57), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_58), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_59), .B(n_631), .Y(n_650) );
INVx1_ASAP7_75t_L g113 ( .A(n_60), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_61), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_62), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_63), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g91 ( .A(n_64), .Y(n_91) );
INVx1_ASAP7_75t_L g121 ( .A(n_64), .Y(n_121) );
BUFx3_ASAP7_75t_L g237 ( .A(n_64), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_65), .B(n_196), .Y(n_284) );
INVx1_ASAP7_75t_L g245 ( .A(n_66), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_67), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g632 ( .A(n_67), .Y(n_632) );
INVx2_ASAP7_75t_L g585 ( .A(n_68), .Y(n_585) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_68), .Y(n_604) );
AND2x2_ASAP7_75t_L g660 ( .A(n_68), .B(n_586), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_69), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_70), .B(n_146), .Y(n_187) );
INVx2_ASAP7_75t_L g576 ( .A(n_71), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_72), .B(n_93), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_73), .Y(n_240) );
INVx1_ASAP7_75t_L g235 ( .A(n_74), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_75), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_75), .A2(n_692), .B1(n_715), .B2(n_726), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g733 ( .A1(n_75), .A2(n_715), .B1(n_734), .B2(n_736), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_76), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_97), .B(n_521), .Y(n_77) );
CKINVDCx6p67_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx11_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
BUFx6f_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_88), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_83), .A2(n_211), .A3(n_224), .B(n_225), .Y(n_210) );
AO31x2_ASAP7_75t_L g386 ( .A1(n_83), .A2(n_211), .A3(n_224), .B(n_225), .Y(n_386) );
BUFx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
OAI21xp33_ASAP7_75t_L g135 ( .A1(n_85), .A2(n_123), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx2_ASAP7_75t_L g165 ( .A(n_86), .Y(n_165) );
BUFx6f_ASAP7_75t_SL g186 ( .A(n_86), .Y(n_186) );
INVx3_ASAP7_75t_L g238 ( .A(n_86), .Y(n_238) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_87), .Y(n_688) );
AO21x2_ASAP7_75t_L g741 ( .A1(n_88), .A2(n_687), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
AOI21x1_ASAP7_75t_L g194 ( .A1(n_90), .A2(n_195), .B(n_197), .Y(n_194) );
AOI22x1_ASAP7_75t_L g212 ( .A1(n_90), .A2(n_118), .B1(n_213), .B2(n_219), .Y(n_212) );
BUFx3_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g185 ( .A(n_91), .Y(n_185) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
INVx2_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
INVx2_ASAP7_75t_L g290 ( .A(n_95), .Y(n_290) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g117 ( .A(n_96), .Y(n_117) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND3x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_425), .C(n_471), .Y(n_98) );
NOR2xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_369), .Y(n_99) );
NAND3xp33_ASAP7_75t_SL g100 ( .A(n_101), .B(n_306), .C(n_341), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_166), .B1(n_293), .B2(n_300), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_141), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g421 ( .A(n_105), .B(n_169), .Y(n_421) );
AND2x4_ASAP7_75t_L g434 ( .A(n_105), .B(n_329), .Y(n_434) );
AND2x2_ASAP7_75t_L g465 ( .A(n_105), .B(n_350), .Y(n_465) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_105), .Y(n_498) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x6_ASAP7_75t_L g318 ( .A(n_106), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_SL g330 ( .A(n_106), .B(n_297), .Y(n_330) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g296 ( .A(n_107), .Y(n_296) );
OAI21x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_122), .B(n_135), .Y(n_107) );
AOI21x1_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_114), .B(n_118), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_113), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g175 ( .A(n_111), .Y(n_175) );
INVx2_ASAP7_75t_L g196 ( .A(n_111), .Y(n_196) );
INVx3_ASAP7_75t_L g215 ( .A(n_111), .Y(n_215) );
INVx2_ASAP7_75t_L g221 ( .A(n_111), .Y(n_221) );
INVx2_ASAP7_75t_L g288 ( .A(n_111), .Y(n_288) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_112), .Y(n_132) );
INVx2_ASAP7_75t_L g205 ( .A(n_112), .Y(n_205) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g177 ( .A(n_116), .Y(n_177) );
INVx2_ASAP7_75t_L g180 ( .A(n_116), .Y(n_180) );
INVx2_ASAP7_75t_L g198 ( .A(n_116), .Y(n_198) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_117), .Y(n_183) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_119), .A2(n_150), .B(n_153), .Y(n_149) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g242 ( .A(n_120), .Y(n_242) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx3_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_127), .Y(n_122) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
INVx1_ASAP7_75t_L g299 ( .A(n_124), .Y(n_299) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g147 ( .A(n_125), .Y(n_147) );
BUFx2_ASAP7_75t_L g255 ( .A(n_125), .Y(n_255) );
INVx1_ASAP7_75t_L g140 ( .A(n_126), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_128), .A2(n_220), .B1(n_222), .B2(n_223), .Y(n_219) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
INVx1_ASAP7_75t_L g268 ( .A(n_132), .Y(n_268) );
INVxp67_ASAP7_75t_L g224 ( .A(n_136), .Y(n_224) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_140), .Y(n_137) );
AOI21x1_ASAP7_75t_L g231 ( .A1(n_138), .A2(n_139), .B(n_140), .Y(n_231) );
OR2x2_ASAP7_75t_L g410 ( .A(n_141), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g431 ( .A(n_141), .B(n_318), .Y(n_431) );
BUFx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g338 ( .A(n_142), .Y(n_338) );
AND2x2_ASAP7_75t_L g345 ( .A(n_142), .B(n_297), .Y(n_345) );
INVx2_ASAP7_75t_L g350 ( .A(n_142), .Y(n_350) );
AND2x2_ASAP7_75t_L g365 ( .A(n_142), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g375 ( .A(n_142), .B(n_189), .Y(n_375) );
OR2x2_ASAP7_75t_L g391 ( .A(n_142), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g420 ( .A(n_142), .Y(n_420) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2x1_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI21x1_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_156), .B(n_161), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_151), .A2(n_244), .B1(n_246), .B2(n_248), .Y(n_243) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_152), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_159), .Y(n_156) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_160), .A2(n_174), .B(n_176), .Y(n_173) );
NOR2x1_ASAP7_75t_SL g161 ( .A(n_162), .B(n_163), .Y(n_161) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_162), .Y(n_171) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_208), .B1(n_270), .B2(n_274), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g458 ( .A(n_168), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_188), .Y(n_168) );
BUFx3_ASAP7_75t_L g272 ( .A(n_169), .Y(n_272) );
AND2x2_ASAP7_75t_L g363 ( .A(n_169), .B(n_338), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_169), .Y(n_366) );
AND2x2_ASAP7_75t_L g480 ( .A(n_169), .B(n_296), .Y(n_480) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_170), .Y(n_402) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_187), .Y(n_170) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_171), .A2(n_212), .B(n_304), .Y(n_303) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_171), .A2(n_172), .B(n_187), .Y(n_329) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_178), .B(n_186), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_181), .B(n_184), .Y(n_178) );
INVx2_ASAP7_75t_L g217 ( .A(n_180), .Y(n_217) );
INVxp67_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_183), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_184), .A2(n_266), .B(n_267), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_184), .A2(n_283), .B(n_284), .Y(n_282) );
BUFx10_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g201 ( .A(n_185), .Y(n_201) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_186), .A2(n_257), .B(n_265), .Y(n_256) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_188), .Y(n_378) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_189), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_189), .B(n_296), .Y(n_411) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g319 ( .A(n_190), .Y(n_319) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_190), .Y(n_392) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_207), .Y(n_191) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_193), .A2(n_207), .B(n_298), .Y(n_297) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_199), .B(n_206), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_202), .B(n_203), .Y(n_199) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_206), .A2(n_282), .B(n_285), .Y(n_281) );
INVx2_ASAP7_75t_L g371 ( .A(n_208), .Y(n_371) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_226), .Y(n_208) );
INVx1_ASAP7_75t_L g336 ( .A(n_209), .Y(n_336) );
INVx1_ASAP7_75t_L g368 ( .A(n_209), .Y(n_368) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g354 ( .A(n_210), .Y(n_354) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OAI22x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_216), .B1(n_217), .B2(n_218), .Y(n_213) );
INVxp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVxp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVxp67_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_222), .Y(n_738) );
INVx1_ASAP7_75t_L g304 ( .A(n_225), .Y(n_304) );
INVx1_ASAP7_75t_L g504 ( .A(n_226), .Y(n_504) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_226), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_251), .Y(n_226) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_227), .B(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g340 ( .A(n_227), .Y(n_340) );
INVx1_ASAP7_75t_L g382 ( .A(n_227), .Y(n_382) );
AND2x2_ASAP7_75t_L g441 ( .A(n_227), .B(n_252), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_227), .B(n_305), .Y(n_463) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g301 ( .A(n_228), .B(n_252), .Y(n_301) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_232), .B(n_249), .Y(n_228) );
AO21x1_ASAP7_75t_L g314 ( .A1(n_229), .A2(n_232), .B(n_249), .Y(n_314) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g249 ( .A(n_230), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_243), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_236), .B1(n_239), .B2(n_241), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NOR3xp33_ASAP7_75t_L g244 ( .A(n_237), .B(n_238), .C(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g263 ( .A(n_237), .Y(n_263) );
INVx2_ASAP7_75t_L g291 ( .A(n_237), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_238), .B(n_242), .Y(n_241) );
NOR3xp33_ASAP7_75t_L g246 ( .A(n_238), .B(n_242), .C(n_247), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_245), .A2(n_721), .B1(n_722), .B2(n_725), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_245), .Y(n_725) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_252), .Y(n_276) );
INVx3_ASAP7_75t_L g310 ( .A(n_252), .Y(n_310) );
INVx2_ASAP7_75t_L g323 ( .A(n_252), .Y(n_323) );
AND2x2_ASAP7_75t_L g327 ( .A(n_252), .B(n_303), .Y(n_327) );
INVx1_ASAP7_75t_L g351 ( .A(n_252), .Y(n_351) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_256), .B(n_269), .Y(n_253) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_254), .A2(n_281), .B(n_292), .Y(n_280) );
BUFx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_260), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_272), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g389 ( .A(n_272), .Y(n_389) );
OR2x2_ASAP7_75t_L g430 ( .A(n_272), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
OR2x2_ASAP7_75t_L g510 ( .A(n_275), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g326 ( .A(n_278), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_278), .B(n_310), .Y(n_359) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_278), .B(n_309), .Y(n_469) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
AND2x2_ASAP7_75t_L g312 ( .A(n_279), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g424 ( .A(n_279), .B(n_303), .Y(n_424) );
INVx1_ASAP7_75t_L g447 ( .A(n_279), .Y(n_447) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
O2A1O1Ixp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_289), .C(n_291), .Y(n_285) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI211xp5_ASAP7_75t_L g306 ( .A1(n_295), .A2(n_307), .B(n_315), .C(n_331), .Y(n_306) );
AND2x2_ASAP7_75t_L g455 ( .A(n_295), .B(n_419), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_295), .B(n_350), .Y(n_508) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
AND2x4_ASAP7_75t_L g344 ( .A(n_296), .B(n_329), .Y(n_344) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AOI32xp33_ASAP7_75t_L g432 ( .A1(n_300), .A2(n_374), .A3(n_433), .B1(n_435), .B2(n_437), .Y(n_432) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g423 ( .A(n_301), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_302), .B(n_382), .Y(n_398) );
AND2x2_ASAP7_75t_L g451 ( .A(n_302), .B(n_340), .Y(n_451) );
AND2x2_ASAP7_75t_L g514 ( .A(n_302), .B(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
OR2x2_ASAP7_75t_L g385 ( .A(n_305), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AOI21xp33_ASAP7_75t_SL g404 ( .A1(n_308), .A2(n_362), .B(n_403), .Y(n_404) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
BUFx2_ASAP7_75t_L g449 ( .A(n_309), .Y(n_449) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_310), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g414 ( .A(n_310), .B(n_386), .Y(n_414) );
INVx1_ASAP7_75t_L g348 ( .A(n_311), .Y(n_348) );
OR2x2_ASAP7_75t_L g394 ( .A(n_311), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_312), .Y(n_415) );
AND2x2_ASAP7_75t_L g456 ( .A(n_312), .B(n_354), .Y(n_456) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g322 ( .A(n_314), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_314), .B(n_361), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B1(n_325), .B2(n_328), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_317), .B(n_365), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_317), .A2(n_487), .B1(n_489), .B2(n_491), .Y(n_486) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g407 ( .A(n_318), .B(n_350), .Y(n_407) );
AND2x2_ASAP7_75t_L g335 ( .A(n_319), .B(n_329), .Y(n_335) );
INVx2_ASAP7_75t_L g520 ( .A(n_320), .Y(n_520) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g428 ( .A(n_322), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g437 ( .A(n_322), .B(n_424), .Y(n_437) );
AND2x2_ASAP7_75t_L g476 ( .A(n_322), .B(n_368), .Y(n_476) );
AND2x2_ASAP7_75t_L g495 ( .A(n_322), .B(n_459), .Y(n_495) );
INVx1_ASAP7_75t_L g342 ( .A(n_324), .Y(n_342) );
OAI321xp33_ASAP7_75t_L g512 ( .A1(n_325), .A2(n_401), .A3(n_435), .B1(n_513), .B2(n_516), .C(n_519), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_326), .B(n_468), .Y(n_511) );
INVx1_ASAP7_75t_L g395 ( .A(n_327), .Y(n_395) );
AND2x4_ASAP7_75t_L g461 ( .A(n_327), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g482 ( .A(n_328), .Y(n_482) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g374 ( .A(n_329), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
NOR4xp25_ASAP7_75t_L g331 ( .A(n_332), .B(n_336), .C(n_337), .D(n_339), .Y(n_331) );
NAND2x1_ASAP7_75t_L g372 ( .A(n_332), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_333), .A2(n_408), .B1(n_455), .B2(n_456), .Y(n_454) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OAI322xp33_ASAP7_75t_L g493 ( .A1(n_336), .A2(n_494), .A3(n_496), .B1(n_502), .B2(n_505), .C1(n_506), .C2(n_510), .Y(n_493) );
AND2x2_ASAP7_75t_L g453 ( .A(n_337), .B(n_421), .Y(n_453) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g436 ( .A(n_338), .B(n_392), .Y(n_436) );
INVx1_ASAP7_75t_L g459 ( .A(n_338), .Y(n_459) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2x1_ASAP7_75t_L g408 ( .A(n_340), .B(n_385), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_346), .C(n_357), .Y(n_341) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g417 ( .A(n_344), .Y(n_417) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_344), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g403 ( .A(n_345), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_349), .B(n_352), .C(n_355), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g509 ( .A(n_350), .B(n_480), .Y(n_509) );
INVx2_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
OR2x6_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx2_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_354), .B(n_441), .Y(n_440) );
NAND2xp33_ASAP7_75t_SL g491 ( .A(n_355), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OAI32xp33_ASAP7_75t_L g357 ( .A1(n_356), .A2(n_358), .A3(n_362), .B1(n_364), .B2(n_367), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_356), .B(n_459), .Y(n_505) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g468 ( .A(n_360), .Y(n_468) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g439 ( .A(n_366), .B(n_411), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_387), .C(n_405), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_376), .B2(n_379), .Y(n_370) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
O2A1O1Ixp5_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_417), .B(n_418), .C(n_422), .Y(n_416) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_375), .Y(n_474) );
INVx1_ASAP7_75t_L g518 ( .A(n_375), .Y(n_518) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g485 ( .A(n_381), .Y(n_485) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g490 ( .A(n_382), .B(n_447), .Y(n_490) );
INVx1_ASAP7_75t_L g397 ( .A(n_383), .Y(n_397) );
NOR2x1p5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g448 ( .A(n_386), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .B1(n_396), .B2(n_399), .C(n_404), .Y(n_387) );
INVx1_ASAP7_75t_L g443 ( .A(n_388), .Y(n_443) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g478 ( .A(n_391), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_393), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g470 ( .A(n_402), .B(n_436), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_409), .B2(n_412), .C(n_416), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
AND2x4_ASAP7_75t_L g489 ( .A(n_413), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g488 ( .A(n_414), .B(n_463), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_R g492 ( .A(n_421), .Y(n_492) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_438), .C(n_442), .D(n_457), .Y(n_425) );
OAI21xp33_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_430), .B(n_432), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_SL g438 ( .A1(n_430), .A2(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_434), .A2(n_470), .B(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI221xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_444), .B1(n_450), .B2(n_452), .C(n_454), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_444), .A2(n_458), .B1(n_460), .B2(n_464), .C(n_466), .Y(n_457) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g484 ( .A(n_446), .Y(n_484) );
AND2x4_ASAP7_75t_L g503 ( .A(n_446), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g500 ( .A(n_447), .Y(n_500) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_459), .B(n_482), .C(n_483), .D(n_485), .Y(n_481) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_493), .C(n_512), .Y(n_471) );
NAND4xp25_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .C(n_481), .D(n_486), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_480), .Y(n_501) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_SL g496 ( .A(n_497), .B(n_501), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_680), .B2(n_691), .C(n_732), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_523), .A2(n_733), .B1(n_737), .B2(n_739), .Y(n_732) );
INVxp33_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_580), .C(n_622), .Y(n_524) );
OAI31xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_539), .A3(n_553), .B(n_572), .Y(n_525) );
CKINVDCx8_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g550 ( .A(n_531), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g558 ( .A(n_531), .B(n_552), .Y(n_558) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g567 ( .A(n_532), .B(n_552), .Y(n_567) );
AND2x4_ASAP7_75t_L g536 ( .A(n_533), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g541 ( .A(n_533), .Y(n_541) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_533), .A2(n_554), .B(n_563), .Y(n_553) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g548 ( .A(n_534), .Y(n_548) );
AND2x4_ASAP7_75t_L g654 ( .A(n_534), .B(n_575), .Y(n_654) );
OR2x2_ASAP7_75t_L g704 ( .A(n_534), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g714 ( .A(n_534), .B(n_705), .Y(n_714) );
CKINVDCx14_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_537), .B(n_701), .C(n_703), .Y(n_700) );
AND2x4_ASAP7_75t_L g711 ( .A(n_537), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x4_ASAP7_75t_L g543 ( .A(n_538), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g627 ( .A(n_538), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx8_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
CKINVDCx8_ASAP7_75t_R g641 ( .A(n_543), .Y(n_641) );
AND2x4_ASAP7_75t_L g562 ( .A(n_544), .B(n_551), .Y(n_562) );
INVx1_ASAP7_75t_L g628 ( .A(n_544), .Y(n_628) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g636 ( .A(n_548), .B(n_575), .Y(n_636) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_549), .Y(n_639) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_550), .Y(n_570) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B1(n_559), .B2(n_560), .Y(n_554) );
INVx5_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx12f_ASAP7_75t_L g631 ( .A(n_562), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_568), .B2(n_571), .Y(n_563) );
BUFx4f_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_569), .A2(n_641), .B1(n_645), .B2(n_646), .Y(n_644) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g590 ( .A1(n_571), .A2(n_591), .B1(n_594), .B2(n_595), .C1(n_605), .C2(n_608), .Y(n_590) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_577), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g705 ( .A(n_576), .Y(n_705) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g621 ( .A(n_578), .Y(n_621) );
BUFx3_ASAP7_75t_L g679 ( .A(n_578), .Y(n_679) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g635 ( .A(n_579), .Y(n_635) );
INVx1_ASAP7_75t_L g653 ( .A(n_579), .Y(n_653) );
OAI31xp33_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_609), .A3(n_611), .B(n_619), .Y(n_580) );
OR2x6_ASAP7_75t_L g582 ( .A(n_583), .B(n_587), .Y(n_582) );
OR2x2_ASAP7_75t_SL g610 ( .A(n_583), .B(n_606), .Y(n_610) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx2_ASAP7_75t_L g598 ( .A(n_585), .Y(n_598) );
AND2x4_ASAP7_75t_L g662 ( .A(n_585), .B(n_593), .Y(n_662) );
INVx2_ASAP7_75t_L g593 ( .A(n_586), .Y(n_593) );
INVx2_ASAP7_75t_L g601 ( .A(n_586), .Y(n_601) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g591 ( .A(n_588), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_SL g608 ( .A(n_588), .B(n_603), .Y(n_608) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g676 ( .A(n_589), .B(n_670), .Y(n_676) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g667 ( .A(n_593), .Y(n_667) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_598), .B(n_601), .Y(n_615) );
AND2x4_ASAP7_75t_L g618 ( .A(n_598), .B(n_601), .Y(n_618) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g666 ( .A(n_604), .B(n_667), .Y(n_666) );
INVx3_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g617 ( .A(n_606), .B(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_614), .A2(n_657), .B(n_658), .C(n_663), .Y(n_656) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_614), .A2(n_649), .B(n_672), .C(n_673), .Y(n_671) );
BUFx12f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
CKINVDCx8_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_643), .C(n_655), .Y(n_622) );
NOR3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_633), .C(n_637), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_629), .B1(n_630), .B2(n_632), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g648 ( .A(n_626), .Y(n_648) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
AND2x6_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .C(n_651), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B(n_650), .Y(n_647) );
CKINVDCx8_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
AND2x6_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_671), .B(n_677), .Y(n_655) );
BUFx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx4_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g674 ( .A(n_665), .Y(n_674) );
INVx5_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx4_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
INVx3_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g698 ( .A(n_688), .Y(n_698) );
AND2x2_ASAP7_75t_L g742 ( .A(n_689), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_690), .B(n_698), .Y(n_697) );
INVx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g735 ( .A(n_694), .Y(n_735) );
INVx5_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x6_ASAP7_75t_L g695 ( .A(n_696), .B(n_706), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVxp67_ASAP7_75t_L g730 ( .A(n_697), .Y(n_730) );
INVx1_ASAP7_75t_L g743 ( .A(n_698), .Y(n_743) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_700), .B(n_710), .Y(n_731) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
CKINVDCx11_ASAP7_75t_R g708 ( .A(n_702), .Y(n_708) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
XOR2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_720), .Y(n_715) );
XNOR2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
XOR2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx4f_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
BUFx6f_ASAP7_75t_SL g736 ( .A(n_728), .Y(n_736) );
INVx4_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
endmodule