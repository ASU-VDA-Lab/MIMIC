module fake_jpeg_27267_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_1),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_61),
.Y(n_82)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_59),
.Y(n_80)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_66),
.B1(n_60),
.B2(n_58),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_63),
.B1(n_64),
.B2(n_55),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_76),
.B1(n_84),
.B2(n_54),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_52),
.B1(n_51),
.B2(n_62),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_43),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_71),
.B1(n_65),
.B2(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_94),
.Y(n_107)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_93),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_98),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_56),
.B1(n_46),
.B2(n_49),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_3),
.Y(n_118)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_118),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_99),
.B1(n_92),
.B2(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_115),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_44),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_117),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_109),
.B1(n_101),
.B2(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_90),
.C(n_86),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_26),
.C(n_12),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_2),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_3),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_50),
.B(n_108),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_123),
.B(n_132),
.Y(n_139)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_124),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_90),
.B(n_22),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_19),
.B(n_24),
.C(n_25),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_130),
.C(n_27),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_8),
.B(n_13),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_135),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_14),
.C(n_17),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_136),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_139),
.C(n_140),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_141),
.B(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_127),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_137),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_137),
.Y(n_154)
);


endmodule