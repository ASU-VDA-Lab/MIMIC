module fake_jpeg_31255_n_83 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_83);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_83;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_5),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_28),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_10),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_20),
.B(n_19),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_47),
.B1(n_41),
.B2(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_19),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_56),
.C(n_34),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_59),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_18),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_66),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_50),
.B1(n_41),
.B2(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_21),
.B1(n_34),
.B2(n_12),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_55),
.C(n_60),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_61),
.C(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_72),
.B(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_68),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_77),
.A2(n_71),
.B(n_64),
.Y(n_79)
);

OAI31xp33_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_76),
.A3(n_5),
.B(n_9),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_3),
.B(n_9),
.C(n_34),
.Y(n_82)
);

OAI21x1_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_80),
.B(n_12),
.Y(n_83)
);


endmodule