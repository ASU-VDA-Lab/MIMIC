module fake_jpeg_12124_n_585 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_585);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_585;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_60),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_62),
.Y(n_195)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_63),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_66),
.Y(n_173)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_70),
.Y(n_199)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_75),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_80),
.B(n_85),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_109),
.Y(n_123)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_18),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_86),
.Y(n_197)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_18),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_95),
.B(n_99),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_18),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_104),
.Y(n_139)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_105),
.B(n_107),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_31),
.B(n_15),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_106),
.B(n_29),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_108),
.B(n_110),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_33),
.B1(n_48),
.B2(n_20),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_117),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_34),
.B(n_13),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_26),
.C(n_24),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_20),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_20),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_146),
.B1(n_192),
.B2(n_10),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_33),
.B1(n_56),
.B2(n_26),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_128),
.A2(n_129),
.B1(n_135),
.B2(n_156),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_61),
.A2(n_49),
.B1(n_46),
.B2(n_37),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_48),
.B1(n_49),
.B2(n_46),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_133),
.A2(n_140),
.B1(n_187),
.B2(n_134),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_56),
.B1(n_36),
.B2(n_35),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_138),
.B(n_142),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_48),
.B1(n_37),
.B2(n_30),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_106),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_68),
.A2(n_19),
.B1(n_36),
.B2(n_35),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_27),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_148),
.B(n_159),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_23),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_165),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_70),
.A2(n_27),
.B1(n_24),
.B2(n_29),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_28),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_161),
.B(n_164),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_28),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_97),
.B(n_30),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_8),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_103),
.B(n_19),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_168),
.B(n_176),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_74),
.A2(n_48),
.B1(n_1),
.B2(n_3),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_170),
.A2(n_184),
.B1(n_193),
.B2(n_181),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_0),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_79),
.B(n_0),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_186),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_104),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_195),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_89),
.A2(n_13),
.B1(n_1),
.B2(n_3),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_0),
.C(n_4),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_198),
.C(n_150),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_114),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_117),
.B(n_5),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_188),
.B(n_158),
.Y(n_261)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

BUFx4f_ASAP7_75t_SL g252 ( 
.A(n_190),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_92),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_100),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_200),
.A2(n_261),
.B(n_271),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_152),
.B(n_165),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_201),
.B(n_242),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_160),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_202),
.B(n_251),
.C(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_205),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_207),
.B(n_210),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_130),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_96),
.B1(n_98),
.B2(n_10),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g296 ( 
.A1(n_211),
.A2(n_246),
.B1(n_215),
.B2(n_217),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_126),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_212),
.B(n_214),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_213),
.A2(n_200),
.B1(n_201),
.B2(n_228),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_215),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_216),
.Y(n_328)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_217),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_12),
.B1(n_166),
.B2(n_193),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_218),
.A2(n_220),
.B(n_259),
.Y(n_318)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_222),
.B(n_245),
.Y(n_321)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_139),
.A2(n_147),
.B1(n_149),
.B2(n_174),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_224),
.A2(n_240),
.B1(n_249),
.B2(n_255),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_226),
.Y(n_295)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_227),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_132),
.B(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_231),
.Y(n_312)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_232),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_145),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_234),
.B(n_239),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_124),
.A2(n_150),
.B1(n_189),
.B2(n_131),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_123),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_238),
.B(n_244),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_127),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_139),
.A2(n_147),
.B1(n_149),
.B2(n_183),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

OR2x2_ASAP7_75t_SL g243 ( 
.A(n_157),
.B(n_172),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_243),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_139),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_178),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_122),
.A2(n_183),
.B1(n_198),
.B2(n_167),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_247),
.A2(n_262),
.B1(n_266),
.B2(n_269),
.Y(n_300)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_248),
.B(n_250),
.Y(n_279)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_131),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_253),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_181),
.B(n_137),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_189),
.A2(n_199),
.B1(n_163),
.B2(n_197),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_137),
.B(n_197),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_256),
.B(n_260),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_163),
.B(n_199),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_268),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_194),
.B(n_179),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_153),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_134),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

INVx11_ASAP7_75t_SL g305 ( 
.A(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_153),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_265),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_124),
.A2(n_173),
.B1(n_134),
.B2(n_151),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_153),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_169),
.B(n_173),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_169),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_169),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_151),
.B(n_158),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_209),
.B(n_158),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_272),
.B(n_290),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_249),
.A2(n_219),
.B1(n_218),
.B2(n_222),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_280),
.A2(n_293),
.B1(n_329),
.B2(n_294),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_281),
.A2(n_309),
.B1(n_275),
.B2(n_321),
.Y(n_336)
);

OR2x2_ASAP7_75t_SL g284 ( 
.A(n_243),
.B(n_201),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_284),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_209),
.B(n_225),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_200),
.A2(n_251),
.B(n_202),
.C(n_203),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_308),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_219),
.A2(n_211),
.B1(n_246),
.B2(n_258),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_296),
.B(n_318),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_202),
.A2(n_246),
.B1(n_211),
.B2(n_259),
.Y(n_301)
);

AO21x2_ASAP7_75t_L g349 ( 
.A1(n_301),
.A2(n_296),
.B(n_278),
.Y(n_349)
);

OR2x4_ASAP7_75t_L g306 ( 
.A(n_237),
.B(n_206),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_273),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_229),
.B(n_230),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_211),
.A2(n_246),
.B1(n_257),
.B2(n_254),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_226),
.B(n_231),
.C(n_268),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_331),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_205),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_291),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_252),
.A2(n_264),
.B(n_242),
.C(n_241),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_323),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_204),
.B(n_227),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_312),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_260),
.A2(n_248),
.B1(n_250),
.B2(n_216),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_208),
.A2(n_232),
.B1(n_269),
.B2(n_270),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_330),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_252),
.B(n_262),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_304),
.Y(n_332)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_309),
.A2(n_236),
.B1(n_247),
.B2(n_252),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_333),
.A2(n_336),
.B1(n_352),
.B2(n_354),
.Y(n_398)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_287),
.Y(n_334)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_325),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_337),
.B(n_346),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_275),
.B(n_290),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_355),
.Y(n_382)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_341),
.Y(n_384)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_343),
.B(n_344),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_285),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_349),
.A2(n_356),
.B1(n_313),
.B2(n_315),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_322),
.B(n_307),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_350),
.B(n_353),
.Y(n_409)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_311),
.Y(n_351)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_281),
.A2(n_278),
.B1(n_276),
.B2(n_274),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_277),
.B(n_326),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_276),
.A2(n_293),
.B1(n_280),
.B2(n_274),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_308),
.A2(n_289),
.B1(n_296),
.B2(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_359),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_289),
.A2(n_292),
.B1(n_317),
.B2(n_284),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_303),
.B(n_272),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_364),
.Y(n_396)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_288),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_372),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_327),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_302),
.A2(n_286),
.B1(n_294),
.B2(n_300),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_373),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_294),
.B(n_331),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_305),
.C(n_328),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_282),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_370),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_297),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_371),
.B(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_279),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_316),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_324),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_283),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_319),
.B(n_310),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_SL g380 ( 
.A(n_335),
.B(n_286),
.C(n_324),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_394),
.Y(n_423)
);

O2A1O1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_323),
.B(n_319),
.C(n_324),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_383),
.A2(n_345),
.B(n_351),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_386),
.A2(n_333),
.B1(n_367),
.B2(n_334),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_358),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_404),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_366),
.A2(n_315),
.B1(n_283),
.B2(n_313),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_347),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_392),
.B(n_393),
.C(n_377),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_374),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_339),
.B(n_299),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_411),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_344),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_413),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_375),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_408),
.B(n_415),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_337),
.B(n_299),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_343),
.B(n_328),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_376),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_354),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_416),
.B(n_352),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_415),
.A2(n_376),
.B(n_348),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_418),
.A2(n_419),
.B(n_446),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_372),
.B(n_335),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_377),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_430),
.C(n_439),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_414),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_436),
.Y(n_451)
);

AOI22x1_ASAP7_75t_L g425 ( 
.A1(n_386),
.A2(n_365),
.B1(n_349),
.B2(n_355),
.Y(n_425)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_407),
.B(n_332),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_426),
.B(n_397),
.Y(n_463)
);

XNOR2x1_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_405),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_429),
.A2(n_435),
.B1(n_437),
.B2(n_412),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_347),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_395),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_433),
.B(n_396),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_449),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_391),
.A2(n_336),
.B1(n_349),
.B2(n_367),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_381),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_388),
.A2(n_349),
.B1(n_368),
.B2(n_361),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_382),
.B(n_346),
.C(n_357),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_394),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_441),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_408),
.B(n_349),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_443),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_410),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_349),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_444),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_385),
.A2(n_350),
.B(n_340),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_385),
.B(n_342),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_406),
.C(n_379),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_448),
.A2(n_383),
.B(n_379),
.Y(n_467)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_363),
.C(n_359),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_387),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_402),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_393),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_454),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_430),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_455),
.B(n_459),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_402),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_398),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_400),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_463),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_398),
.C(n_411),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_468),
.C(n_470),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_443),
.B(n_409),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_466),
.B(n_401),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_467),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_379),
.C(n_397),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_416),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_444),
.A2(n_441),
.B1(n_448),
.B2(n_423),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_473),
.A2(n_429),
.B1(n_417),
.B2(n_436),
.Y(n_494)
);

OAI21xp33_ASAP7_75t_L g475 ( 
.A1(n_422),
.A2(n_390),
.B(n_409),
.Y(n_475)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_476),
.A2(n_427),
.B1(n_440),
.B2(n_425),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_412),
.C(n_387),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_478),
.C(n_468),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_419),
.B(n_432),
.Y(n_478)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_452),
.B(n_456),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_488),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_469),
.A2(n_423),
.B(n_445),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_484),
.A2(n_460),
.B(n_470),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_460),
.B(n_434),
.CI(n_427),
.CON(n_485),
.SN(n_485)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_478),
.Y(n_507)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_487),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_456),
.B(n_455),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_476),
.A2(n_425),
.B1(n_417),
.B2(n_438),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_489),
.B(n_491),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_490),
.B(n_493),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_454),
.B(n_400),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_494),
.A2(n_503),
.B1(n_467),
.B2(n_464),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_451),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_496),
.B(n_499),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_451),
.B(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_498),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_462),
.A2(n_413),
.B1(n_442),
.B2(n_420),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_500),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_502),
.B(n_472),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_453),
.A2(n_431),
.B1(n_401),
.B2(n_403),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_457),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_465),
.C(n_477),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_517),
.C(n_522),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_507),
.A2(n_506),
.B(n_522),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_508),
.A2(n_521),
.B1(n_492),
.B2(n_489),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_497),
.Y(n_509)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_509),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_384),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_480),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_514),
.B(n_524),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_459),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_482),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_473),
.C(n_453),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_484),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_518),
.B(n_523),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_494),
.A2(n_458),
.B1(n_474),
.B2(n_471),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_490),
.B(n_458),
.C(n_474),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_487),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_481),
.B(n_384),
.Y(n_524)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_526),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_536),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_505),
.A2(n_486),
.B1(n_485),
.B2(n_493),
.Y(n_528)
);

OAI21xp33_ASAP7_75t_L g548 ( 
.A1(n_528),
.A2(n_520),
.B(n_519),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_508),
.A2(n_499),
.B1(n_485),
.B2(n_495),
.Y(n_530)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_525),
.C(n_399),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_521),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_532),
.A2(n_528),
.B1(n_530),
.B2(n_526),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_535),
.B(n_537),
.Y(n_553)
);

FAx1_ASAP7_75t_SL g536 ( 
.A(n_517),
.B(n_486),
.CI(n_483),
.CON(n_536),
.SN(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_488),
.C(n_483),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_510),
.A2(n_503),
.B(n_403),
.Y(n_539)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_539),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_515),
.C(n_520),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_513),
.B(n_399),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_541),
.B(n_542),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_516),
.B(n_399),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_545),
.Y(n_566)
);

MAJx2_ASAP7_75t_L g557 ( 
.A(n_548),
.B(n_554),
.C(n_527),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_529),
.B(n_535),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_549),
.B(n_550),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_529),
.B(n_509),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_534),
.B(n_519),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_551),
.B(n_552),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_534),
.B(n_362),
.C(n_341),
.Y(n_552)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_557),
.Y(n_571)
);

OAI21xp33_ASAP7_75t_L g558 ( 
.A1(n_556),
.A2(n_532),
.B(n_533),
.Y(n_558)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_558),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_553),
.B(n_538),
.C(n_537),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_560),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_533),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_546),
.A2(n_540),
.B(n_539),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_561),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_556),
.B(n_536),
.C(n_555),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_563),
.B(n_567),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_555),
.A2(n_536),
.B1(n_547),
.B2(n_543),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_564),
.Y(n_573)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_548),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_565),
.B(n_544),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_566),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_575),
.B(n_579),
.Y(n_581)
);

NAND2x1_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_567),
.Y(n_576)
);

MAJx2_ASAP7_75t_L g582 ( 
.A(n_576),
.B(n_558),
.C(n_557),
.Y(n_582)
);

AO21x1_ASAP7_75t_L g577 ( 
.A1(n_572),
.A2(n_564),
.B(n_562),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_577),
.A2(n_578),
.B(n_568),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_570),
.A2(n_573),
.B(n_571),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_568),
.Y(n_579)
);

BUFx24_ASAP7_75t_SL g583 ( 
.A(n_580),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_583),
.B(n_581),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_582),
.Y(n_585)
);


endmodule