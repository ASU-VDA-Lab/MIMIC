module fake_netlist_5_388_n_323 (n_91, n_82, n_122, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_323);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_323;

wire n_137;
wire n_294;
wire n_318;
wire n_194;
wire n_316;
wire n_248;
wire n_124;
wire n_146;
wire n_136;
wire n_315;
wire n_268;
wire n_127;
wire n_235;
wire n_226;
wire n_155;
wire n_284;
wire n_245;
wire n_139;
wire n_280;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_321;
wire n_292;
wire n_212;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_147;
wire n_307;
wire n_150;
wire n_209;
wire n_259;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_204;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_282;
wire n_132;
wire n_281;
wire n_240;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_152;
wire n_317;
wire n_195;
wire n_227;
wire n_271;
wire n_123;
wire n_167;
wire n_234;
wire n_308;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_158;
wire n_138;
wire n_264;
wire n_276;
wire n_163;
wire n_183;
wire n_185;
wire n_243;
wire n_169;
wire n_255;
wire n_215;
wire n_196;
wire n_211;
wire n_218;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_287;
wire n_141;
wire n_145;
wire n_313;
wire n_216;
wire n_168;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_140;
wire n_299;
wire n_303;
wire n_296;
wire n_241;
wire n_184;
wire n_144;
wire n_165;
wire n_213;
wire n_129;
wire n_197;
wire n_236;
wire n_249;
wire n_304;
wire n_203;
wire n_274;
wire n_277;
wire n_149;
wire n_309;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_239;
wire n_310;
wire n_170;
wire n_161;
wire n_273;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_312;
wire n_210;
wire n_176;
wire n_182;
wire n_143;
wire n_237;
wire n_180;
wire n_207;
wire n_229;
wire n_177;
wire n_233;
wire n_205;
wire n_246;
wire n_179;
wire n_125;
wire n_269;
wire n_128;
wire n_285;
wire n_232;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_193;
wire n_251;
wire n_160;
wire n_154;
wire n_148;
wire n_300;
wire n_159;
wire n_175;
wire n_262;
wire n_238;
wire n_319;
wire n_242;
wire n_200;
wire n_162;
wire n_222;
wire n_199;
wire n_187;
wire n_166;
wire n_256;
wire n_305;
wire n_278;

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_29),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_43),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_45),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_49),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_17),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_36),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_14),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_R g138 ( 
.A(n_6),
.B(n_104),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_38),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_55),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_26),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_105),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_SL g146 ( 
.A(n_56),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_46),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_71),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_47),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_51),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_68),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_R g156 ( 
.A(n_52),
.B(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_48),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_97),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_53),
.Y(n_160)
);

INVxp33_ASAP7_75t_SL g161 ( 
.A(n_74),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_30),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_35),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_21),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_31),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_76),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_2),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_79),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_42),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_32),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_25),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_59),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVxp33_ASAP7_75t_SL g179 ( 
.A(n_41),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_111),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_57),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_13),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_34),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_90),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_66),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_28),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_61),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_60),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_11),
.B(n_44),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_82),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_80),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_101),
.B(n_87),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

INVxp33_ASAP7_75t_SL g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_33),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_40),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_10),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_83),
.B(n_73),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_58),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_118),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_4),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_88),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_50),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_133),
.A2(n_0),
.B1(n_1),
.B2(n_8),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_127),
.B(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_0),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_141),
.B(n_12),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_123),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_161),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_22),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_23),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_24),
.Y(n_228)
);

OR2x2_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_37),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_39),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_65),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_135),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_144),
.A2(n_67),
.B1(n_72),
.B2(n_78),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_147),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_151),
.B(n_84),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_152),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_L g241 ( 
.A(n_138),
.B(n_156),
.Y(n_241)
);

NOR2x1p5_ASAP7_75t_L g242 ( 
.A(n_154),
.B(n_89),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_125),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_140),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_179),
.B(n_95),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_162),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_132),
.B(n_148),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_166),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_149),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_167),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_197),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_184),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_222),
.B(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_249),
.B(n_182),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_218),
.B(n_215),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_209),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_242),
.B(n_183),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_231),
.B(n_181),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_219),
.B(n_206),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_203),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_225),
.B(n_168),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_227),
.B(n_165),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_239),
.B(n_185),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_224),
.B(n_164),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_200),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_SL g271 ( 
.A(n_232),
.B(n_202),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_246),
.B(n_155),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_177),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_237),
.B(n_194),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_223),
.B(n_192),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_234),
.B(n_236),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_233),
.B(n_241),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_233),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_229),
.B1(n_158),
.B2(n_189),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_275),
.B1(n_261),
.B2(n_273),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

AO21x2_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_266),
.B(n_267),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_233),
.B1(n_252),
.B2(n_250),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_257),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_128),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_R g294 ( 
.A(n_278),
.B(n_190),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_286),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_193),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_R g298 ( 
.A(n_281),
.B(n_274),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_262),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_R g300 ( 
.A(n_282),
.B(n_163),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_256),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

AO31x2_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_195),
.A3(n_186),
.B(n_153),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_288),
.B1(n_290),
.B2(n_286),
.Y(n_304)
);

NAND2x1_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_196),
.Y(n_305)
);

OAI33xp33_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_226),
.A3(n_221),
.B1(n_254),
.B2(n_247),
.B3(n_243),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_269),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

AO221x2_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_198),
.B1(n_207),
.B2(n_180),
.C(n_204),
.Y(n_309)
);

AO221x2_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_175),
.B1(n_201),
.B2(n_199),
.C(n_230),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_SL g311 ( 
.A(n_308),
.B(n_298),
.Y(n_311)
);

AO221x2_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_238),
.B1(n_240),
.B2(n_220),
.C(n_294),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_301),
.B1(n_300),
.B2(n_188),
.C(n_136),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_296),
.B(n_305),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_311),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_312),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_309),
.B1(n_315),
.B2(n_172),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_143),
.B1(n_142),
.B2(n_159),
.Y(n_321)
);

AOI222xp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_139),
.B1(n_191),
.B2(n_126),
.C1(n_306),
.C2(n_130),
.Y(n_322)
);

OAI221xp5_ASAP7_75t_R g323 ( 
.A1(n_322),
.A2(n_170),
.B1(n_150),
.B2(n_145),
.C(n_314),
.Y(n_323)
);


endmodule