module real_jpeg_10899_n_12 (n_290, n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_289, n_3, n_10, n_9, n_12);

input n_290;
input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_289;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_181;
wire n_85;
wire n_102;
wire n_274;
wire n_256;
wire n_101;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_11),
.B1(n_18),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_1),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_1),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_66),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_10),
.B(n_26),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_11),
.B1(n_18),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_29),
.B1(n_71),
.B2(n_72),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_70)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_6),
.A2(n_46),
.B(n_70),
.C(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_6),
.B(n_46),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_10),
.B(n_72),
.Y(n_106)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_11),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_9),
.A2(n_19),
.B1(n_71),
.B2(n_72),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_9),
.A2(n_19),
.B1(n_46),
.B2(n_47),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_11),
.B1(n_18),
.B2(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_43),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_10),
.A2(n_25),
.B(n_45),
.C(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_27),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_22),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_11),
.A2(n_22),
.B(n_58),
.C(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_35),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_33),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_30),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_15),
.B(n_37),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_27),
.B2(n_28),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_17),
.A2(n_24),
.B(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_21),
.A2(n_24),
.B1(n_57),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_25),
.A2(n_44),
.B(n_45),
.C(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_27),
.A2(n_56),
.B(n_65),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_32),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_79),
.B(n_287),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_38),
.B(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_38),
.B(n_285),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_54),
.CI(n_59),
.CON(n_38),
.SN(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_43),
.B1(n_51),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_42),
.B(n_137),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_43),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_43),
.A2(n_51),
.B1(n_135),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_44),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_46),
.A2(n_50),
.B(n_58),
.Y(n_141)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_58),
.B(n_75),
.C(n_106),
.Y(n_105)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_52),
.B(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_57),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_58),
.B(n_70),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.C(n_67),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_60),
.A2(n_67),
.B1(n_265),
.B2(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_61),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_62),
.A2(n_63),
.B1(n_151),
.B2(n_157),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_62),
.B(n_151),
.C(n_194),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_62),
.A2(n_63),
.B1(n_134),
.B2(n_138),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_62),
.B(n_134),
.C(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_62),
.A2(n_63),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_67),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_67),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_78),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_69),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_70),
.A2(n_76),
.B1(n_100),
.B2(n_103),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_70),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_229),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_284),
.B(n_286),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_257),
.A3(n_277),
.B1(n_282),
.B2(n_283),
.C(n_289),
.Y(n_80)
);

AOI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_213),
.A3(n_233),
.B1(n_251),
.B2(n_256),
.C(n_290),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_182),
.C(n_210),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_162),
.B(n_181),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_147),
.B(n_161),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_129),
.B(n_146),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_118),
.B(n_128),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_108),
.B(n_117),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_97),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_97),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_89),
.A2(n_110),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_89),
.B(n_151),
.C(n_156),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B(n_93),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_92),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_92),
.A2(n_144),
.B1(n_189),
.B2(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_94),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_95),
.A2(n_188),
.B(n_190),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_105),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_107),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_134),
.C(n_145),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_98),
.A2(n_107),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B(n_102),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_102),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_103),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_107),
.B(n_187),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B(n_116),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_123),
.C(n_126),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_115),
.A2(n_127),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_115),
.B(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_120),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_126),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_125),
.A2(n_126),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_125),
.B(n_201),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_150),
.C(n_160),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_139),
.B2(n_145),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_138),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_168),
.C(n_172),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_136),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_139),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_143),
.B(n_203),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_148),
.B(n_149),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_157),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_157),
.B(n_239),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_173),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_174),
.C(n_180),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_171),
.B2(n_172),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_168),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_172),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_171),
.A2(n_172),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_171),
.A2(n_172),
.B1(n_271),
.B2(n_275),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_171),
.B(n_265),
.C(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_171),
.B(n_275),
.C(n_276),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_205),
.C(n_207),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_174),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_178),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_183),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_195),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_184),
.B(n_195),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_191),
.CI(n_192),
.CON(n_184),
.SN(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_209),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_204),
.C(n_209),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_214),
.A2(n_252),
.B(n_255),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_215),
.B(n_216),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_232),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_224),
.B2(n_225),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_225),
.C(n_232),
.Y(n_234)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_220),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_231),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_227),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_228),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_242),
.B(n_244),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_235),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_249),
.B2(n_250),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_241),
.B1(n_247),
.B2(n_248),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_238),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_248),
.C(n_250),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_259),
.C(n_267),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_259),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_244),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_269),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_269),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_262),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_268),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.Y(n_269)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);


endmodule