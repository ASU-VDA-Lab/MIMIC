module real_jpeg_14372_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_162)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_6),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_6),
.A2(n_38),
.B1(n_75),
.B2(n_76),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_8),
.A2(n_75),
.B1(n_76),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_133),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_133),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_75),
.B1(n_76),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_10),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_147),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_147),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_11),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_55),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_75),
.B1(n_76),
.B2(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_13),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_72),
.B(n_75),
.C(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_13),
.B(n_82),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_13),
.B(n_61),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_SL g214 ( 
.A1(n_13),
.A2(n_61),
.B(n_200),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_13),
.B(n_30),
.C(n_49),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_144),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_13),
.B(n_88),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_14),
.A2(n_75),
.B1(n_76),
.B2(n_80),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_14),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_80),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_80),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_15),
.A2(n_33),
.B1(n_75),
.B2(n_76),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_15),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_15),
.A2(n_33),
.B1(n_61),
.B2(n_62),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_136),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_19),
.B(n_112),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_84),
.B2(n_111),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.C(n_69),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_22),
.A2(n_23),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_266)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_27),
.A2(n_35),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_122),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_28),
.A2(n_34),
.B(n_162),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_28),
.A2(n_161),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_29),
.A2(n_124),
.B(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_31),
.B1(n_49),
.B2(n_50),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_31),
.B(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_35),
.A2(n_36),
.B(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_35),
.A2(n_121),
.B(n_123),
.Y(n_120)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_35),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_35),
.A2(n_36),
.B1(n_229),
.B2(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_36),
.B(n_37),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_36),
.B(n_144),
.Y(n_235)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_42),
.A2(n_52),
.B(n_93),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_SL g201 ( 
.A(n_43),
.B(n_58),
.C(n_62),
.Y(n_201)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_44),
.A2(n_59),
.B(n_199),
.C(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_44),
.B(n_223),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_94),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_54),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_47),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_47),
.A2(n_53),
.B1(n_195),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_47),
.A2(n_53),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_47),
.A2(n_53),
.B1(n_216),
.B2(n_226),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_52),
.B(n_144),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_94),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_69),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_64),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_57),
.A2(n_66),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_57),
.A2(n_66),
.B1(n_150),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_57),
.A2(n_66),
.B1(n_172),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_62),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_73),
.B(n_144),
.Y(n_165)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_66),
.A2(n_151),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_68),
.B(n_88),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_79),
.B(n_81),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_71),
.B1(n_79),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_70),
.A2(n_71),
.B1(n_132),
.B2(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_82),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_96),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B(n_95),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_88),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_91),
.A2(n_154),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_103),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_118),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_117),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_118),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.C(n_130),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_119),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_125),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_268)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_271),
.B(n_276),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_184),
.B(n_262),
.C(n_270),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_173),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_139),
.B(n_173),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_157),
.C(n_166),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_152),
.C(n_156),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_158),
.B1(n_166),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_174),
.B(n_182),
.C(n_183),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_176),
.B(n_177),
.C(n_180),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_260),
.B(n_261),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_204),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_187),
.B(n_190),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_196),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_196),
.B1(n_197),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_202),
.B1(n_203),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_217),
.B(n_259),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_215),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_253),
.B(n_258),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_243),
.B(n_252),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_232),
.B(n_242),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_227),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_224),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_241),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_248),
.C(n_251),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_266),
.C(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);


endmodule