module fake_jpeg_31010_n_140 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_SL g37 ( 
.A(n_2),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_1),
.Y(n_58)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_49),
.Y(n_80)
);

BUFx2_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_66),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_32),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_15),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_82),
.Y(n_93)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_34),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_39),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_38),
.B(n_48),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_99),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_96),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_16),
.B(n_30),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_8),
.B(n_9),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_21),
.Y(n_111)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_5),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_5),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_109),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_19),
.C(n_7),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_115),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_14),
.C(n_18),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_25),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_94),
.B1(n_100),
.B2(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_112),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_129),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_130),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

OAI31xp33_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_85),
.A3(n_121),
.B(n_113),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_129),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_132),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_105),
.C(n_122),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_120),
.C(n_123),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_125),
.Y(n_140)
);


endmodule