module fake_jpeg_11381_n_48 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_48);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_48;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_26),
.Y(n_27)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_20),
.B(n_4),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_4),
.B(n_5),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_2),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_17),
.B1(n_21),
.B2(n_5),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_37),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_31),
.B(n_10),
.Y(n_43)
);

AND2x6_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_27),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_30),
.CI(n_41),
.CON(n_42),
.SN(n_42)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_6),
.C(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_44),
.Y(n_46)
);

OAI21x1_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_12),
.B(n_13),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_14),
.Y(n_48)
);


endmodule