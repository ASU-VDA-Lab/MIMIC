module fake_netlist_5_848_n_47 (n_8, n_10, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_11, n_6, n_1, n_47);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_11;
input n_6;
input n_1;

output n_47;

wire n_29;
wire n_16;
wire n_43;
wire n_12;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_42;
wire n_22;
wire n_45;
wire n_24;
wire n_28;
wire n_46;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_38;
wire n_35;
wire n_32;
wire n_41;
wire n_17;
wire n_19;
wire n_37;
wire n_15;
wire n_26;
wire n_30;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_20;
wire n_39;

CKINVDCx6p67_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_5),
.B1(n_9),
.B2(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_10),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_4),
.A2(n_5),
.B(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

OAI22x1_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_2),
.B1(n_21),
.B2(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

AOI211x1_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_13),
.B(n_16),
.C(n_17),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B(n_23),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_19),
.C(n_12),
.Y(n_29)
);

OAI21x1_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_17),
.B(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OR2x6_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_30),
.Y(n_32)
);

OAI21x1_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_17),
.B(n_14),
.Y(n_33)
);

OAI21x1_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_17),
.B(n_14),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_14),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_31),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_35),
.B(n_32),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_35),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_41),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_37),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_32),
.B1(n_20),
.B2(n_18),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_18),
.B(n_20),
.Y(n_45)
);

AOI221xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_18),
.B1(n_20),
.B2(n_33),
.C(n_32),
.Y(n_46)
);

OR2x6_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_45),
.Y(n_47)
);


endmodule