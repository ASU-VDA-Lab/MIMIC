module fake_jpeg_30968_n_453 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_59),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_49),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_15),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_50),
.B(n_52),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_87),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_19),
.B1(n_33),
.B2(n_20),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_23),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_24),
.B(n_14),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_66),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_12),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_93),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_78),
.Y(n_109)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_11),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_47),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_39),
.B(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_98),
.B(n_33),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_35),
.B1(n_16),
.B2(n_45),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_100),
.A2(n_113),
.B1(n_120),
.B2(n_20),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_26),
.B1(n_16),
.B2(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_122),
.B1(n_33),
.B2(n_20),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_52),
.A2(n_27),
.B(n_23),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_105),
.A2(n_18),
.A3(n_17),
.B1(n_37),
.B2(n_41),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_143),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_49),
.A2(n_35),
.B1(n_16),
.B2(n_42),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_61),
.B(n_19),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_116),
.B(n_140),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_51),
.B(n_16),
.C(n_41),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_46),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_53),
.A2(n_46),
.B1(n_36),
.B2(n_47),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_61),
.B(n_19),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_55),
.B(n_47),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_26),
.B1(n_71),
.B2(n_78),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_147),
.A2(n_165),
.B1(n_182),
.B2(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_123),
.B1(n_108),
.B2(n_133),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_102),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_153),
.B(n_157),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_154),
.A2(n_163),
.B(n_167),
.Y(n_235)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_156),
.B(n_189),
.Y(n_206)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_96),
.A2(n_18),
.B1(n_93),
.B2(n_90),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g204 ( 
.A(n_166),
.Y(n_204)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_37),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_98),
.B(n_37),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_41),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_99),
.A2(n_18),
.B1(n_86),
.B2(n_82),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_101),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_185),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_97),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_192),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_195),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_99),
.A2(n_18),
.B1(n_89),
.B2(n_84),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_167),
.B(n_157),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_199),
.A2(n_109),
.B(n_134),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_148),
.A2(n_132),
.B1(n_77),
.B2(n_56),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_218),
.B1(n_220),
.B2(n_104),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_215),
.A2(n_226),
.B1(n_195),
.B2(n_192),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_123),
.B1(n_108),
.B2(n_111),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_68),
.B1(n_57),
.B2(n_92),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_170),
.A2(n_131),
.B1(n_124),
.B2(n_133),
.Y(n_226)
);

NAND2x1_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_94),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_205),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_95),
.B1(n_124),
.B2(n_131),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_151),
.B1(n_126),
.B2(n_187),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_237),
.A2(n_218),
.B1(n_234),
.B2(n_220),
.Y(n_279)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_165),
.B(n_147),
.C(n_94),
.Y(n_241)
);

AO21x2_ASAP7_75t_SL g288 ( 
.A1(n_241),
.A2(n_243),
.B(n_254),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_199),
.A2(n_109),
.B(n_185),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_269),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_166),
.B1(n_161),
.B2(n_169),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_244),
.B(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_246),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_247),
.A2(n_137),
.B(n_201),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_248),
.B(n_261),
.Y(n_278)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_249),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_179),
.Y(n_250)
);

BUFx24_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_153),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_251),
.B(n_260),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_149),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_272),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_253),
.A2(n_266),
.B1(n_261),
.B2(n_258),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_29),
.B(n_17),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_159),
.C(n_168),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_222),
.C(n_227),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_258),
.B(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_200),
.B(n_171),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_202),
.B(n_175),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_263),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_211),
.B(n_197),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_267),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_198),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_265),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_211),
.B(n_17),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_198),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_268),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_208),
.A2(n_29),
.B(n_38),
.C(n_31),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_271),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_40),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_216),
.B(n_40),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_259),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_213),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_276),
.B(n_293),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_279),
.A2(n_253),
.B1(n_266),
.B2(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_245),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_181),
.B1(n_189),
.B2(n_228),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_297),
.B1(n_232),
.B2(n_231),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_285),
.A2(n_243),
.B1(n_265),
.B2(n_268),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_204),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_224),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_224),
.C(n_221),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_298),
.C(n_269),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_238),
.A2(n_228),
.B1(n_29),
.B2(n_233),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_221),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_302),
.A2(n_249),
.B(n_255),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_250),
.B(n_233),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_232),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_303),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_275),
.A2(n_298),
.B(n_302),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_309),
.A2(n_310),
.B1(n_316),
.B2(n_329),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_279),
.A2(n_241),
.B1(n_239),
.B2(n_250),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_275),
.A2(n_252),
.B(n_254),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_333),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_241),
.C(n_254),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_326),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_278),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_286),
.B(n_256),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_319),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_306),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_315),
.B(n_328),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_241),
.B1(n_243),
.B2(n_263),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_291),
.A2(n_241),
.B(n_270),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_318),
.A2(n_321),
.B(n_305),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_289),
.B(n_246),
.Y(n_319)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_243),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_323),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_280),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_287),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_324),
.Y(n_342)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_273),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_327),
.A2(n_331),
.B1(n_288),
.B2(n_323),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_290),
.B(n_299),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_296),
.Y(n_343)
);

AO22x1_ASAP7_75t_L g331 ( 
.A1(n_281),
.A2(n_240),
.B1(n_231),
.B2(n_38),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_288),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_306),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_46),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_335),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_277),
.B(n_46),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_336),
.Y(n_359)
);

AOI21xp33_ASAP7_75t_SL g338 ( 
.A1(n_331),
.A2(n_283),
.B(n_304),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_337),
.C(n_355),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_343),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_341),
.A2(n_321),
.B1(n_318),
.B2(n_310),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_319),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_362),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_346),
.A2(n_351),
.B1(n_357),
.B2(n_309),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_274),
.Y(n_373)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_349),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_327),
.A2(n_288),
.B1(n_285),
.B2(n_276),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_281),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_356),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_281),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_334),
.A2(n_288),
.B1(n_300),
.B2(n_307),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_295),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_361),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_334),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_363),
.A2(n_370),
.B1(n_377),
.B2(n_359),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_332),
.C(n_313),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_366),
.C(n_382),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_374),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_312),
.C(n_326),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_308),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_383),
.Y(n_389)
);

AOI21xp33_ASAP7_75t_R g369 ( 
.A1(n_344),
.A2(n_311),
.B(n_317),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_369),
.B(n_379),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_360),
.A2(n_322),
.B1(n_320),
.B2(n_317),
.Y(n_370)
);

AOI221xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_336),
.B1(n_335),
.B2(n_301),
.C(n_324),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_373),
.Y(n_385)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_351),
.A2(n_295),
.B1(n_292),
.B2(n_134),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_380),
.B(n_1),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_38),
.C(n_31),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_38),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_346),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_384),
.A2(n_347),
.B(n_358),
.Y(n_387)
);

AOI21x1_ASAP7_75t_SL g386 ( 
.A1(n_373),
.A2(n_347),
.B(n_341),
.Y(n_386)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_401),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_356),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_393),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_361),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_368),
.Y(n_408)
);

FAx1_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_361),
.CI(n_350),
.CON(n_394),
.SN(n_394)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_394),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_342),
.C(n_353),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_398),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_370),
.A2(n_349),
.B1(n_2),
.B2(n_4),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_31),
.C(n_4),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_382),
.C(n_383),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_375),
.Y(n_403)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_406),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_396),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_389),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_377),
.C(n_365),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_412),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_399),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_381),
.C(n_378),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_415),
.C(n_400),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_372),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_414),
.A2(n_398),
.B(n_5),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_381),
.C(n_5),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_416),
.B(n_417),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_409),
.C(n_392),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_421),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_391),
.C(n_395),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_410),
.A2(n_385),
.B(n_394),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_422),
.B(n_423),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_403),
.A2(n_394),
.B(n_389),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_426),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_404),
.A2(n_4),
.B(n_6),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_414),
.B(n_6),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_6),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_402),
.Y(n_430)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_430),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_425),
.A2(n_402),
.B1(n_7),
.B2(n_8),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_435),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_436),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_6),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_417),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_439),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_418),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_429),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_445),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_432),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_442),
.Y(n_446)
);

AOI21xp33_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_441),
.B(n_431),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_443),
.C(n_421),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_449),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_447),
.B(n_427),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_451),
.B(n_9),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_9),
.Y(n_453)
);


endmodule