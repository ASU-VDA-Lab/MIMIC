module fake_jpeg_7862_n_319 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx12_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_26),
.B1(n_21),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_63),
.B1(n_23),
.B2(n_20),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_54),
.B1(n_23),
.B2(n_20),
.Y(n_88)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_27),
.B1(n_28),
.B2(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_33),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_29),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_68),
.B(n_8),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_60),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_34),
.B1(n_30),
.B2(n_25),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_67),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_19),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_43),
.B1(n_18),
.B2(n_33),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_87),
.B1(n_90),
.B2(n_46),
.Y(n_105)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_34),
.B1(n_30),
.B2(n_18),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_86),
.B1(n_53),
.B2(n_45),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_10),
.Y(n_83)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_95),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_33),
.B1(n_23),
.B2(n_20),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_0),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_99),
.B1(n_101),
.B2(n_87),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_108),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_68),
.B1(n_45),
.B2(n_53),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_45),
.B1(n_61),
.B2(n_62),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_96),
.B1(n_102),
.B2(n_115),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_90),
.B(n_82),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_94),
.B(n_73),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_77),
.Y(n_108)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_121),
.Y(n_130)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_116),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_57),
.A3(n_58),
.B1(n_59),
.B2(n_49),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_89),
.A3(n_85),
.B1(n_74),
.B2(n_69),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_46),
.B(n_50),
.C(n_10),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_123),
.A2(n_124),
.B1(n_148),
.B2(n_103),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_71),
.B1(n_94),
.B2(n_95),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_125),
.A2(n_16),
.B1(n_7),
.B2(n_4),
.Y(n_173)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_127),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_104),
.B1(n_116),
.B2(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_131),
.Y(n_170)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_85),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_118),
.B(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_134),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_85),
.C(n_73),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_151),
.C(n_105),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_141),
.B(n_147),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_140),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_59),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_79),
.B(n_80),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_59),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_80),
.B1(n_9),
.B2(n_11),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_80),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_79),
.C(n_49),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_97),
.A2(n_79),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_111),
.B1(n_113),
.B2(n_122),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_160),
.C(n_171),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_156),
.B(n_132),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_135),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_157),
.A2(n_167),
.B(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_173),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_118),
.C(n_111),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_166),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_175),
.B1(n_181),
.B2(n_155),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_6),
.B1(n_14),
.B2(n_4),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_147),
.B1(n_133),
.B2(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_0),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_79),
.C(n_2),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_79),
.B(n_2),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_130),
.B(n_7),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_7),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_130),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_145),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

XOR2x2_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_132),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_200),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_197),
.B1(n_199),
.B2(n_203),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_183),
.C(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_206),
.Y(n_236)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_208),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_182),
.A2(n_134),
.B1(n_142),
.B2(n_126),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_142),
.B1(n_143),
.B2(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_184),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_209),
.A2(n_204),
.B1(n_187),
.B2(n_203),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_153),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_215),
.C(n_217),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_201),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_218),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_156),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_157),
.C(n_168),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_225),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_189),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_168),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_171),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_174),
.C(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_231),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_173),
.B1(n_166),
.B2(n_176),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_172),
.B(n_162),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_178),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_234),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_177),
.C(n_169),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_235),
.Y(n_256)
);

CKINVDCx11_ASAP7_75t_R g237 ( 
.A(n_232),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_239),
.B1(n_245),
.B2(n_248),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_202),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_197),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_195),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_239),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_214),
.C(n_219),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_223),
.C(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_267),
.C(n_269),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_248),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_228),
.B1(n_209),
.B2(n_191),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_262),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_217),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_219),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_240),
.A2(n_186),
.B1(n_215),
.B2(n_190),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_254),
.B1(n_256),
.B2(n_238),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_226),
.C(n_196),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_246),
.C(n_252),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_268),
.B1(n_271),
.B2(n_251),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_277),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_256),
.B1(n_245),
.B2(n_250),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_279),
.C(n_284),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_253),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_260),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_1),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_255),
.B1(n_249),
.B2(n_241),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_292),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_275),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_272),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_12),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_285),
.C(n_282),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_278),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_167),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_296),
.Y(n_300)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_167),
.A3(n_259),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_296),
.B(n_11),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_291),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_305),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_12),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_14),
.B1(n_15),
.B2(n_3),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_15),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_287),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_309),
.Y(n_312)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_303),
.B(n_288),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_313),
.A2(n_314),
.B(n_306),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_306),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_312),
.B(n_308),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_307),
.C(n_314),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_15),
.B(n_3),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_3),
.Y(n_319)
);


endmodule