module fake_jpeg_2324_n_290 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_4),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_4),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_59),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_4),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_64),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_5),
.B(n_6),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_6),
.C(n_7),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_23),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_84),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_33),
.A2(n_27),
.B1(n_31),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_42),
.B1(n_43),
.B2(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_9),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_9),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_39),
.B(n_10),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_85),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_43),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_88),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_37),
.B1(n_44),
.B2(n_31),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_90),
.B(n_103),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_97),
.A2(n_113),
.B1(n_115),
.B2(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_102),
.B1(n_115),
.B2(n_111),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_50),
.A2(n_25),
.B1(n_41),
.B2(n_36),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_42),
.B1(n_36),
.B2(n_40),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_112),
.B1(n_120),
.B2(n_128),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_60),
.A2(n_26),
.B1(n_45),
.B2(n_12),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_26),
.B1(n_45),
.B2(n_12),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_72),
.B1(n_69),
.B2(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_10),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_11),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_77),
.B1(n_63),
.B2(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_111),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_35),
.B1(n_53),
.B2(n_60),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_85),
.A2(n_73),
.B1(n_57),
.B2(n_50),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_101),
.B1(n_90),
.B2(n_95),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_53),
.A2(n_35),
.B1(n_60),
.B2(n_31),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_89),
.B1(n_93),
.B2(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_107),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_137),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_124),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_174)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_149),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_153),
.B(n_141),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_89),
.A2(n_114),
.B1(n_129),
.B2(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_153),
.B(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_89),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_89),
.A2(n_93),
.B1(n_110),
.B2(n_125),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_98),
.B(n_105),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_103),
.A2(n_97),
.B1(n_114),
.B2(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_94),
.B(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_136),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_161),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_102),
.A2(n_96),
.B1(n_126),
.B2(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_169),
.Y(n_186)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_167),
.Y(n_185)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_131),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_98),
.B(n_105),
.Y(n_169)
);

NOR2x1_ASAP7_75t_R g171 ( 
.A(n_92),
.B(n_95),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_137),
.B(n_170),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_111),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_143),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_181),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_139),
.B(n_166),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_144),
.B(n_171),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_175),
.B(n_176),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_149),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_193),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_191),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_155),
.B1(n_143),
.B2(n_145),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_174),
.B1(n_191),
.B2(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_205),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_156),
.B1(n_166),
.B2(n_168),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_208),
.B(n_209),
.C(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_163),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_214),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_179),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_185),
.C(n_178),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_151),
.B1(n_165),
.B2(n_192),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_174),
.B1(n_188),
.B2(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_194),
.B(n_177),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_210),
.B1(n_204),
.B2(n_198),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_235),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_183),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_229),
.C(n_214),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_202),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_217),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_238),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_194),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_202),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_244),
.B1(n_248),
.B2(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_246),
.B1(n_201),
.B2(n_228),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_233),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_203),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_232),
.B1(n_231),
.B2(n_234),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_255),
.B1(n_231),
.B2(n_246),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_256),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_231),
.B1(n_214),
.B2(n_199),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_231),
.B1(n_196),
.B2(n_228),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_257),
.A2(n_245),
.B(n_247),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_231),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_264),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_266),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_242),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_269),
.A2(n_240),
.B(n_238),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_258),
.C(n_256),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_267),
.A2(n_255),
.B1(n_251),
.B2(n_257),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_275),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_268),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_248),
.B(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_262),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_273),
.B(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_272),
.B1(n_278),
.B2(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_278),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_224),
.B(n_219),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_287),
.C(n_270),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_268),
.Y(n_290)
);


endmodule