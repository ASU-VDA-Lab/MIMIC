module real_jpeg_33165_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_0),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_1),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_1),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_1),
.B(n_276),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_1),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_1),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_2),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_2),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_2),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_2),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_2),
.B(n_63),
.Y(n_159)
);

AND2x4_ASAP7_75t_SL g202 ( 
.A(n_2),
.B(n_203),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_3),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_3),
.B(n_137),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_R g184 ( 
.A(n_3),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_3),
.B(n_284),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_3),
.B(n_500),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_514),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_4),
.B(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_5),
.B(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_5),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_5),
.Y(n_247)
);

NAND2x1_ASAP7_75t_SL g278 ( 
.A(n_5),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_5),
.B(n_181),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g389 ( 
.A(n_5),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_5),
.B(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_8),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_9),
.Y(n_515)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_10),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_10),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_10),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_80),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_10),
.B(n_96),
.Y(n_95)
);

AND2x4_ASAP7_75t_SL g121 ( 
.A(n_10),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_10),
.B(n_63),
.Y(n_470)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_11),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_12),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_13),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_13),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_13),
.B(n_108),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_13),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_13),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_13),
.B(n_344),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_13),
.B(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_14),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_63),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_15),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_15),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_15),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_15),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_15),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_15),
.B(n_428),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_17),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_17),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_17),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_17),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_17),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_17),
.B(n_474),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_17),
.B(n_509),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_484),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_452),
.B(n_482),
.Y(n_20)
);

OA21x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_260),
.B(n_443),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_212),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_162),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_25),
.B(n_163),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_25),
.B(n_163),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_103),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_26),
.B(n_455),
.C(n_456),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_69),
.C(n_89),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_27),
.A2(n_28),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_44),
.C(n_56),
.Y(n_28)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_29),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_39),
.C(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_33),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_36),
.A2(n_42),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_38),
.Y(n_196)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_40),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_41),
.Y(n_145)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_41),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_42),
.B(n_468),
.C(n_470),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_44),
.B(n_56),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.C(n_51),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_45),
.A2(n_46),
.B1(n_201),
.B2(n_202),
.Y(n_510)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_49),
.Y(n_258)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_50),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_51),
.A2(n_52),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_52),
.B(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_52),
.B(n_121),
.C(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_55),
.Y(n_203)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_55),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_57),
.A2(n_141),
.B1(n_142),
.B2(n_146),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_57),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_57),
.B(n_65),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_57),
.B(n_65),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_57),
.B(n_144),
.C(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_57),
.A2(n_146),
.B1(n_343),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_59),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_68),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_61),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_65),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_65),
.A2(n_68),
.B1(n_236),
.B2(n_237),
.Y(n_272)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_69),
.A2(n_90),
.B1(n_91),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_81),
.C(n_86),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_70),
.A2(n_71),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.C(n_79),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_72),
.B(n_75),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_79),
.B(n_178),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g335 ( 
.A(n_79),
.B(n_116),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_80),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_83),
.Y(n_206)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_84),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_85),
.Y(n_341)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_88),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_94),
.C(n_100),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_94),
.A2(n_95),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_94),
.B(n_155),
.C(n_159),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_94),
.A2(n_95),
.B1(n_499),
.B2(n_504),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_96),
.Y(n_285)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_102),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_138),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_104),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_119),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_105),
.B(n_120),
.C(n_127),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_107),
.Y(n_115)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_110),
.A2(n_111),
.B1(n_242),
.B2(n_271),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_110),
.A2(n_111),
.B1(n_201),
.B2(n_202),
.Y(n_477)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_111),
.B(n_242),
.C(n_248),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_111),
.B(n_115),
.C(n_156),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_111),
.B(n_201),
.C(n_473),
.Y(n_512)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_118),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_118),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_124),
.Y(n_480)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.C(n_135),
.Y(n_127)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_129),
.B1(n_135),
.B2(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_131),
.B(n_201),
.C(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_131),
.A2(n_132),
.B1(n_204),
.B2(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_138),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_152),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_139),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.C(n_150),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_146),
.B(n_343),
.Y(n_342)
);

XOR2x1_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_149),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_161),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_160),
.B(n_459),
.C(n_460),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_161),
.Y(n_460)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.C(n_174),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_170),
.B1(n_171),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_215),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_215),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_197),
.C(n_208),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_186),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_177),
.B(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_179),
.A2(n_180),
.B1(n_186),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_SL g306 ( 
.A(n_180),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_184),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_186),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_194),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_196),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.C(n_207),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_201),
.B(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_204),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_207),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_213),
.A2(n_445),
.B(n_451),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_217),
.B(n_218),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g446 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.C(n_228),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_225),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_229),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_253),
.C(n_256),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_230),
.B(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.C(n_241),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_266),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_234),
.A2(n_235),
.B1(n_241),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_240),
.Y(n_431)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_246),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_247),
.B(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_256),
.Y(n_312)
);

XOR2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_319),
.C(n_325),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_310),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_262),
.B(n_310),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.C(n_286),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_264),
.A2(n_265),
.B1(n_288),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_328),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_328),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_272),
.B(n_274),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.C(n_283),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_275),
.B(n_278),
.Y(n_376)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_283),
.B(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_301),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_306),
.C(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_294),
.C(n_300),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_349)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_296),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_349),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_306),
.B2(n_309),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_314),
.C(n_316),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_320),
.A2(n_448),
.B(n_449),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_321),
.B(n_322),
.Y(n_449)
);

OAI21x1_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_350),
.B(n_442),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_330),
.B(n_331),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g442 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.C(n_347),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_332),
.B(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_348),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.C(n_342),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_335),
.A2(n_336),
.B1(n_337),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_379),
.B(n_441),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_377),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_352),
.B(n_377),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.C(n_374),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_357),
.A2(n_358),
.B1(n_375),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_364),
.C(n_369),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_359),
.A2(n_360),
.B1(n_364),
.B2(n_365),
.Y(n_384)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_369),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

OAI21x1_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_399),
.B(n_440),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_396),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_381),
.B(n_396),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.C(n_388),
.Y(n_381)
);

XNOR2x2_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_385),
.A2(n_386),
.B1(n_388),
.B2(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_393),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_389),
.B(n_393),
.Y(n_403)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI21x1_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_434),
.B(n_439),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_420),
.B(n_433),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_413),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_402),
.B(n_413),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_406),
.C(n_408),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_418),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_418),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_427),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_426),
.B(n_432),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_425),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_425),
.Y(n_432)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_436),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_447),
.B(n_450),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.Y(n_453)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_457),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_471),
.C(n_488),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_471),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_462),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g491 ( 
.A(n_463),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_491),
.C(n_492),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_466),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_468),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_478),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_479),
.C(n_481),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_477),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g484 ( 
.A(n_485),
.B(n_513),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

NOR2x1_ASAP7_75t_SL g513 ( 
.A(n_487),
.B(n_489),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_506),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_505),
.Y(n_497)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_499),
.Y(n_504)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_511),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.Y(n_507)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);


endmodule