module real_aes_6431_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_0), .Y(n_683) );
AOI22xp5_ASAP7_75t_SL g426 ( .A1(n_1), .A2(n_191), .B1(n_427), .B2(n_428), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_2), .A2(n_185), .B1(n_333), .B2(n_409), .Y(n_509) );
INVx1_ASAP7_75t_L g476 ( .A(n_3), .Y(n_476) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_4), .A2(n_66), .B1(n_207), .B2(n_359), .C1(n_361), .C2(n_527), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_5), .A2(n_15), .B1(n_242), .B2(n_258), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_6), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_7), .B(n_595), .Y(n_658) );
INVx1_ASAP7_75t_L g473 ( .A(n_8), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_9), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_10), .A2(n_102), .B1(n_412), .B2(n_546), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_11), .A2(n_141), .B1(n_304), .B2(n_368), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_12), .A2(n_94), .B1(n_287), .B2(n_333), .Y(n_574) );
AOI222xp33_ASAP7_75t_L g617 ( .A1(n_13), .A2(n_96), .B1(n_174), .B2(n_319), .C1(n_528), .C2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_14), .A2(n_119), .B1(n_521), .B2(n_522), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_16), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_17), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g311 ( .A1(n_18), .A2(n_63), .B1(n_117), .B2(n_312), .C1(n_314), .C2(n_318), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_19), .B(n_522), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_20), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_21), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_22), .Y(n_498) );
AO22x2_ASAP7_75t_L g257 ( .A1(n_23), .A2(n_67), .B1(n_248), .B2(n_253), .Y(n_257) );
INVx1_ASAP7_75t_L g636 ( .A(n_23), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_24), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_25), .A2(n_160), .B1(n_546), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_26), .A2(n_111), .B1(n_289), .B2(n_428), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_27), .A2(n_167), .B1(n_359), .B2(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_28), .A2(n_128), .B1(n_260), .B2(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_29), .A2(n_221), .B1(n_484), .B2(n_548), .Y(n_547) );
AOI222xp33_ASAP7_75t_L g526 ( .A1(n_30), .A2(n_157), .B1(n_203), .B2(n_361), .C1(n_527), .C2(n_528), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_31), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_32), .A2(n_200), .B1(n_289), .B2(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_33), .B(n_521), .Y(n_615) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_34), .A2(n_71), .B1(n_248), .B2(n_249), .Y(n_255) );
INVx1_ASAP7_75t_L g637 ( .A(n_34), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_35), .A2(n_109), .B1(n_308), .B2(n_320), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_36), .A2(n_133), .B1(n_260), .B2(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_37), .A2(n_64), .B1(n_278), .B2(n_281), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_38), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_39), .A2(n_99), .B1(n_271), .B2(n_335), .Y(n_334) );
AOI222xp33_ASAP7_75t_L g601 ( .A1(n_40), .A2(n_153), .B1(n_209), .B2(n_359), .C1(n_388), .C2(n_527), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_41), .A2(n_52), .B1(n_289), .B2(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_42), .Y(n_582) );
AOI22xp5_ASAP7_75t_SL g423 ( .A1(n_43), .A2(n_131), .B1(n_402), .B2(n_424), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_44), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_45), .A2(n_168), .B1(n_404), .B2(n_654), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_46), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_47), .A2(n_218), .B1(n_407), .B2(n_409), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_48), .A2(n_179), .B1(n_514), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_49), .A2(n_124), .B1(n_368), .B2(n_438), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_50), .A2(n_149), .B1(n_430), .B2(n_548), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_51), .Y(n_488) );
INVx1_ASAP7_75t_L g671 ( .A(n_53), .Y(n_671) );
AOI22xp5_ASAP7_75t_SL g420 ( .A1(n_54), .A2(n_118), .B1(n_421), .B2(n_422), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_55), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_56), .A2(n_178), .B1(n_298), .B2(n_302), .Y(n_439) );
AO22x2_ASAP7_75t_L g370 ( .A1(n_57), .A2(n_371), .B1(n_413), .B2(n_414), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_57), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g356 ( .A1(n_58), .A2(n_134), .B1(n_357), .B2(n_360), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_59), .A2(n_188), .B1(n_404), .B2(n_405), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_60), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_61), .A2(n_193), .B1(n_330), .B2(n_331), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_62), .A2(n_182), .B1(n_297), .B2(n_301), .Y(n_296) );
AOI22xp5_ASAP7_75t_SL g479 ( .A1(n_65), .A2(n_123), .B1(n_260), .B2(n_422), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_68), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_69), .A2(n_115), .B1(n_314), .B2(n_360), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_70), .A2(n_216), .B1(n_424), .B2(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_72), .Y(n_602) );
INVx1_ASAP7_75t_L g229 ( .A(n_73), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_74), .A2(n_105), .B1(n_347), .B2(n_421), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_75), .A2(n_211), .B1(n_516), .B2(n_518), .Y(n_515) );
INVx1_ASAP7_75t_L g554 ( .A(n_76), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_77), .A2(n_103), .B1(n_279), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_78), .A2(n_113), .B1(n_287), .B2(n_292), .Y(n_286) );
AOI22xp5_ASAP7_75t_SL g482 ( .A1(n_79), .A2(n_192), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_80), .A2(n_151), .B1(n_361), .B2(n_368), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_81), .Y(n_337) );
INVx1_ASAP7_75t_L g226 ( .A(n_82), .Y(n_226) );
XOR2x2_ASAP7_75t_L g501 ( .A(n_83), .B(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_84), .A2(n_152), .B1(n_653), .B2(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g449 ( .A(n_85), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_86), .A2(n_127), .B1(n_542), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_87), .A2(n_199), .B1(n_412), .B2(n_612), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_88), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_89), .A2(n_176), .B1(n_359), .B2(n_438), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_90), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_91), .A2(n_140), .B1(n_244), .B2(n_407), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_92), .B(n_521), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_93), .A2(n_146), .B1(n_411), .B2(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_95), .B(n_366), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_97), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_98), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_100), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g540 ( .A(n_101), .Y(n_540) );
INVx1_ASAP7_75t_L g474 ( .A(n_104), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_106), .A2(n_189), .B1(n_272), .B2(n_551), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_107), .A2(n_196), .B1(n_368), .B2(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_108), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_110), .A2(n_148), .B1(n_308), .B2(n_319), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_112), .B(n_528), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_114), .A2(n_217), .B1(n_271), .B2(n_516), .Y(n_575) );
AOI22xp5_ASAP7_75t_SL g559 ( .A1(n_116), .A2(n_560), .B1(n_584), .B2(n_585), .Y(n_559) );
INVx1_ASAP7_75t_L g585 ( .A(n_116), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_120), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_121), .Y(n_619) );
INVx2_ASAP7_75t_L g230 ( .A(n_122), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_125), .A2(n_187), .B1(n_304), .B2(n_308), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_126), .Y(n_563) );
AND2x6_ASAP7_75t_L g225 ( .A(n_129), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_129), .Y(n_630) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_130), .A2(n_186), .B1(n_248), .B2(n_249), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_132), .A2(n_166), .B1(n_524), .B2(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_135), .A2(n_205), .B1(n_339), .B2(n_407), .Y(n_606) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_136), .A2(n_223), .B(n_231), .C(n_638), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_137), .A2(n_164), .B1(n_421), .B2(n_592), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_138), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_139), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_142), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_143), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_144), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_145), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_147), .A2(n_161), .B1(n_343), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_150), .A2(n_208), .B1(n_411), .B2(n_412), .Y(n_410) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_154), .A2(n_201), .B1(n_248), .B2(n_253), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_155), .A2(n_215), .B1(n_319), .B2(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_156), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_158), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_159), .A2(n_204), .B1(n_387), .B2(n_388), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_162), .Y(n_348) );
INVx1_ASAP7_75t_L g446 ( .A(n_163), .Y(n_446) );
INVx1_ASAP7_75t_L g471 ( .A(n_165), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_169), .Y(n_687) );
XOR2xp5_ASAP7_75t_L g639 ( .A(n_170), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_171), .A2(n_220), .B1(n_267), .B2(n_271), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_172), .B(n_428), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_173), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_175), .A2(n_202), .B1(n_272), .B2(n_404), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_177), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_180), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_181), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_183), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_184), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_186), .B(n_635), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_190), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_194), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_195), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_197), .A2(n_206), .B1(n_364), .B2(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_198), .A2(n_325), .B1(n_326), .B2(n_369), .Y(n_324) );
INVx1_ASAP7_75t_L g369 ( .A(n_198), .Y(n_369) );
INVx1_ASAP7_75t_L g633 ( .A(n_201), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_210), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_212), .A2(n_214), .B1(n_505), .B2(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g248 ( .A(n_213), .Y(n_248) );
INVx1_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
OA22x2_ASAP7_75t_L g237 ( .A1(n_219), .A2(n_238), .B1(n_239), .B2(n_322), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_219), .Y(n_238) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_226), .Y(n_629) );
OA21x2_ASAP7_75t_L g669 ( .A1(n_227), .A2(n_628), .B(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_556), .B1(n_557), .B2(n_624), .C(n_625), .Y(n_231) );
INVx1_ASAP7_75t_L g624 ( .A(n_232), .Y(n_624) );
XOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_500), .Y(n_232) );
XOR2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_416), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AO22x1_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_323), .B2(n_415), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_SL g322 ( .A(n_239), .Y(n_322) );
NAND4xp75_ASAP7_75t_L g239 ( .A(n_240), .B(n_276), .C(n_295), .D(n_311), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_266), .Y(n_240) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_243), .A2(n_408), .B1(n_462), .B2(n_463), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_243), .A2(n_577), .B1(n_578), .B2(n_580), .Y(n_576) );
INVx2_ASAP7_75t_L g592 ( .A(n_243), .Y(n_592) );
INVx3_ASAP7_75t_L g610 ( .A(n_243), .Y(n_610) );
INVx6_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx3_ASAP7_75t_L g343 ( .A(n_244), .Y(n_343) );
BUFx3_ASAP7_75t_L g402 ( .A(n_244), .Y(n_402) );
BUFx3_ASAP7_75t_L g514 ( .A(n_244), .Y(n_514) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_254), .Y(n_244) );
AND2x2_ASAP7_75t_L g280 ( .A(n_245), .B(n_264), .Y(n_280) );
AND2x6_ASAP7_75t_L g283 ( .A(n_245), .B(n_284), .Y(n_283) );
AND2x6_ASAP7_75t_L g313 ( .A(n_245), .B(n_310), .Y(n_313) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_251), .Y(n_245) );
AND2x2_ASAP7_75t_L g291 ( .A(n_246), .B(n_252), .Y(n_291) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g262 ( .A(n_247), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_247), .B(n_252), .Y(n_275) );
AND2x2_ASAP7_75t_L g307 ( .A(n_247), .B(n_257), .Y(n_307) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g253 ( .A(n_250), .Y(n_253) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g263 ( .A(n_252), .Y(n_263) );
INVx1_ASAP7_75t_L g317 ( .A(n_252), .Y(n_317) );
AND2x2_ASAP7_75t_L g270 ( .A(n_254), .B(n_262), .Y(n_270) );
AND2x6_ASAP7_75t_L g302 ( .A(n_254), .B(n_291), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_254), .B(n_291), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_254), .B(n_262), .Y(n_469) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g265 ( .A(n_255), .Y(n_265) );
INVx1_ASAP7_75t_L g274 ( .A(n_255), .Y(n_274) );
OR2x2_ASAP7_75t_L g285 ( .A(n_255), .B(n_256), .Y(n_285) );
AND2x2_ASAP7_75t_L g310 ( .A(n_255), .B(n_257), .Y(n_310) );
AND2x2_ASAP7_75t_L g264 ( .A(n_256), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx3_ASAP7_75t_L g508 ( .A(n_261), .Y(n_508) );
BUFx3_ASAP7_75t_L g546 ( .A(n_261), .Y(n_546) );
BUFx3_ASAP7_75t_L g651 ( .A(n_261), .Y(n_651) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_262), .B(n_264), .Y(n_351) );
INVx1_ASAP7_75t_L g309 ( .A(n_263), .Y(n_309) );
AND2x4_ASAP7_75t_L g290 ( .A(n_264), .B(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g293 ( .A(n_264), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g316 ( .A(n_265), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g395 ( .A(n_265), .Y(n_395) );
BUFx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_268), .Y(n_335) );
INVx2_ASAP7_75t_L g517 ( .A(n_268), .Y(n_517) );
INVx4_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g404 ( .A(n_269), .Y(n_404) );
INVx3_ASAP7_75t_L g422 ( .A(n_269), .Y(n_422) );
INVx5_ASAP7_75t_L g551 ( .A(n_269), .Y(n_551) );
INVx1_ASAP7_75t_L g653 ( .A(n_269), .Y(n_653) );
INVx8_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g405 ( .A(n_272), .Y(n_405) );
BUFx2_ASAP7_75t_L g518 ( .A(n_272), .Y(n_518) );
INVx6_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g553 ( .A(n_273), .Y(n_553) );
INVx1_ASAP7_75t_L g654 ( .A(n_273), .Y(n_654) );
OR2x6_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g306 ( .A(n_274), .Y(n_306) );
INVx1_ASAP7_75t_L g294 ( .A(n_275), .Y(n_294) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_286), .Y(n_276) );
BUFx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_SL g347 ( .A(n_280), .Y(n_347) );
INVx2_ASAP7_75t_L g408 ( .A(n_280), .Y(n_408) );
BUFx2_ASAP7_75t_SL g424 ( .A(n_280), .Y(n_424) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g421 ( .A(n_282), .Y(n_421) );
INVx4_ASAP7_75t_L g483 ( .A(n_282), .Y(n_483) );
INVx4_ASAP7_75t_L g505 ( .A(n_282), .Y(n_505) );
INVx11_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx11_ASAP7_75t_L g340 ( .A(n_283), .Y(n_340) );
AND2x4_ASAP7_75t_L g300 ( .A(n_284), .B(n_291), .Y(n_300) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g377 ( .A(n_285), .B(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx4_ASAP7_75t_L g330 ( .A(n_288), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_288), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_685) );
INVx4_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx3_ASAP7_75t_L g409 ( .A(n_290), .Y(n_409) );
BUFx3_ASAP7_75t_L g430 ( .A(n_290), .Y(n_430) );
INVx2_ASAP7_75t_L g458 ( .A(n_290), .Y(n_458) );
BUFx3_ASAP7_75t_L g612 ( .A(n_290), .Y(n_612) );
INVx1_ASAP7_75t_L g378 ( .A(n_291), .Y(n_378) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx3_ASAP7_75t_L g333 ( .A(n_293), .Y(n_333) );
BUFx3_ASAP7_75t_L g412 ( .A(n_293), .Y(n_412) );
BUFx3_ASAP7_75t_L g427 ( .A(n_293), .Y(n_427) );
INVx1_ASAP7_75t_L g467 ( .A(n_293), .Y(n_467) );
BUFx3_ASAP7_75t_L g484 ( .A(n_293), .Y(n_484) );
BUFx2_ASAP7_75t_SL g647 ( .A(n_293), .Y(n_647) );
BUFx2_ASAP7_75t_SL g689 ( .A(n_293), .Y(n_689) );
AND2x2_ASAP7_75t_L g428 ( .A(n_294), .B(n_395), .Y(n_428) );
AND2x2_ASAP7_75t_SL g295 ( .A(n_296), .B(n_303), .Y(n_295) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_298), .Y(n_366) );
INVx5_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g521 ( .A(n_299), .Y(n_521) );
INVx2_ASAP7_75t_L g595 ( .A(n_299), .Y(n_595) );
INVx4_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx4f_ASAP7_75t_L g364 ( .A(n_302), .Y(n_364) );
BUFx2_ASAP7_75t_L g522 ( .A(n_302), .Y(n_522) );
BUFx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g438 ( .A(n_305), .Y(n_438) );
INVx1_ASAP7_75t_L g525 ( .A(n_305), .Y(n_525) );
BUFx2_ASAP7_75t_L g597 ( .A(n_305), .Y(n_597) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x4_ASAP7_75t_L g315 ( .A(n_307), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g320 ( .A(n_307), .B(n_321), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_307), .B(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_308), .Y(n_368) );
BUFx3_ASAP7_75t_L g542 ( .A(n_308), .Y(n_542) );
BUFx2_ASAP7_75t_SL g660 ( .A(n_308), .Y(n_660) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g399 ( .A(n_309), .Y(n_399) );
INVx1_ASAP7_75t_L g398 ( .A(n_310), .Y(n_398) );
INVx3_ASAP7_75t_L g385 ( .A(n_312), .Y(n_385) );
BUFx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx4_ASAP7_75t_L g354 ( .A(n_313), .Y(n_354) );
INVx2_ASAP7_75t_L g434 ( .A(n_313), .Y(n_434) );
INVx2_ASAP7_75t_SL g454 ( .A(n_313), .Y(n_454) );
INVx2_ASAP7_75t_L g539 ( .A(n_313), .Y(n_539) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_313), .Y(n_618) );
BUFx4f_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
BUFx2_ASAP7_75t_L g387 ( .A(n_315), .Y(n_387) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_315), .Y(n_528) );
INVx1_ASAP7_75t_L g321 ( .A(n_317), .Y(n_321) );
BUFx4f_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g389 ( .A(n_319), .Y(n_389) );
BUFx12f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_320), .Y(n_697) );
INVx1_ASAP7_75t_L g415 ( .A(n_323), .Y(n_415) );
XNOR2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_370), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_327), .B(n_352), .Y(n_326) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_336), .C(n_344), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_341), .B2(n_342), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx5_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_SL g411 ( .A(n_340), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_340), .B(n_473), .Y(n_472) );
INVx4_ASAP7_75t_L g579 ( .A(n_340), .Y(n_579) );
INVx1_ASAP7_75t_L g645 ( .A(n_340), .Y(n_645) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_348), .B2(n_349), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_346), .A2(n_349), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g684 ( .A(n_350), .Y(n_684) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_351), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_362), .Y(n_352) );
OAI21xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_355), .B(n_356), .Y(n_353) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_354), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
INVx4_ASAP7_75t_L g527 ( .A(n_354), .Y(n_527) );
OAI21xp5_ASAP7_75t_SL g565 ( .A1(n_354), .A2(n_566), .B(n_567), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_354), .A2(n_695), .B1(n_696), .B2(n_698), .C(n_699), .Y(n_694) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_358), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_452) );
INVx4_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g497 ( .A(n_359), .Y(n_497) );
BUFx4f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .C(n_367), .Y(n_362) );
INVx1_ASAP7_75t_SL g413 ( .A(n_371), .Y(n_413) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_372), .B(n_400), .Y(n_371) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_383), .C(n_390), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_379), .B2(n_380), .Y(n_373) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_377), .A2(n_446), .B(n_447), .Y(n_445) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_377), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g562 ( .A1(n_377), .A2(n_450), .B1(n_563), .B2(n_564), .Y(n_562) );
BUFx3_ASAP7_75t_L g702 ( .A(n_377), .Y(n_702) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_380), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_487) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g657 ( .A(n_381), .Y(n_657) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g450 ( .A(n_382), .Y(n_450) );
OAI21xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_386), .Y(n_383) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_396), .B2(n_397), .Y(n_390) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_SL g489 ( .A(n_393), .Y(n_489) );
INVx4_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_394), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_448) );
BUFx2_ASAP7_75t_L g570 ( .A(n_397), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_397), .A2(n_489), .B1(n_692), .B2(n_693), .Y(n_691) );
OR2x6_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
AND4x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .C(n_406), .D(n_410), .Y(n_400) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g548 ( .A(n_408), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_441), .B2(n_499), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
XOR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_440), .Y(n_418) );
NAND4xp75_ASAP7_75t_SL g419 ( .A(n_420), .B(n_423), .C(n_425), .D(n_431), .Y(n_419) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_436), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_435), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx2_ASAP7_75t_L g499 ( .A(n_441), .Y(n_499) );
XOR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_475), .Y(n_441) );
XNOR2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_474), .Y(n_442) );
AND3x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_456), .C(n_464), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .C(n_452), .Y(n_444) );
OA211x2_ASAP7_75t_L g613 ( .A1(n_450), .A2(n_614), .B(n_615), .C(n_616), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
OAI21xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_459), .B(n_460), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_470), .C(n_472), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_465) );
XNOR2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
NAND3x1_ASAP7_75t_SL g477 ( .A(n_478), .B(n_481), .C(n_486), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_491), .C(n_495), .Y(n_486) );
OAI22xp5_ASAP7_75t_SL g568 ( .A1(n_489), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
OAI21xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_493), .B(n_494), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_529), .B1(n_530), .B2(n_555), .Y(n_500) );
INVx1_ASAP7_75t_L g555 ( .A(n_501), .Y(n_555) );
NAND4xp75_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .C(n_519), .D(n_526), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_SL g519 ( .A(n_520), .B(n_523), .Y(n_519) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
XOR2x2_ASAP7_75t_SL g531 ( .A(n_532), .B(n_554), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_533), .B(n_543), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
NAND3xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .C(n_537), .Y(n_534) );
OAI21xp5_ASAP7_75t_SL g538 ( .A1(n_539), .A2(n_540), .B(n_541), .Y(n_538) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_549), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
CKINVDCx14_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_586), .B1(n_622), .B2(n_623), .Y(n_557) );
INVx1_ASAP7_75t_L g622 ( .A(n_558), .Y(n_622) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g584 ( .A(n_560), .Y(n_584) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_572), .Y(n_560) );
NOR3xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .C(n_568), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .C(n_581), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g623 ( .A(n_586), .Y(n_623) );
AO22x1_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_603), .B1(n_620), .B2(n_621), .Y(n_586) );
INVx2_ASAP7_75t_SL g620 ( .A(n_587), .Y(n_620) );
XOR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_602), .Y(n_587) );
NAND4xp75_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .C(n_598), .D(n_601), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_SL g593 ( .A(n_594), .B(n_596), .Y(n_593) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_SL g621 ( .A(n_603), .Y(n_621) );
XOR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_619), .Y(n_603) );
NAND4xp75_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .C(n_613), .D(n_617), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g682 ( .A(n_610), .Y(n_682) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .Y(n_626) );
OR2x2_ASAP7_75t_SL g706 ( .A(n_627), .B(n_632), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_628), .Y(n_663) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_629), .B(n_666), .Y(n_670) );
CKINVDCx16_ASAP7_75t_R g666 ( .A(n_630), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OAI322xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_662), .A3(n_664), .B1(n_667), .B2(n_671), .C1(n_672), .C2(n_704), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND4xp75_ASAP7_75t_L g642 ( .A(n_643), .B(n_648), .C(n_655), .D(n_661), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
BUFx4f_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
OA211x2_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B(n_658), .C(n_659), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_657), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_669), .Y(n_668) );
XOR2xp5_ASAP7_75t_SL g674 ( .A(n_671), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_690), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .C(n_685), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_680) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .C(n_700), .Y(n_690) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_705), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
endmodule