module fake_jpeg_23804_n_131 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_12),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_34),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_32),
.B(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_41),
.B1(n_22),
.B2(n_20),
.Y(n_43)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_3),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_21),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_5),
.C(n_7),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_27),
.B(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_25),
.B1(n_40),
.B2(n_35),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_15),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_9),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_19),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_14),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_33),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_14),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_68),
.B1(n_74),
.B2(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_38),
.B1(n_35),
.B2(n_39),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_72),
.Y(n_84)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_57),
.B1(n_62),
.B2(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_45),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_27),
.B(n_14),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_77),
.B(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_8),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_14),
.B1(n_29),
.B2(n_18),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_78),
.B1(n_73),
.B2(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_85),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_50),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_78),
.B(n_65),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_44),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_81),
.B1(n_78),
.B2(n_74),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_100),
.C(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_69),
.C(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_45),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_69),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_69),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.C(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_65),
.C(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_47),
.B1(n_90),
.B2(n_70),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_104),
.C(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_89),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_116),
.C(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_102),
.C(n_84),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_108),
.C(n_117),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_83),
.B1(n_70),
.B2(n_47),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_89),
.C(n_55),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

AOI31xp67_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_120),
.A3(n_72),
.B(n_13),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_125),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_128),
.B(n_10),
.Y(n_131)
);


endmodule