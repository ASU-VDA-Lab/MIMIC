module real_aes_8715_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_0), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_1), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_2), .A2(n_10), .B1(n_422), .B2(n_424), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_3), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_4), .A2(n_190), .B1(n_280), .B2(n_285), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_5), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_6), .A2(n_399), .B1(n_438), .B2(n_439), .Y(n_398) );
INVx1_ASAP7_75t_L g438 ( .A(n_6), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g335 ( .A1(n_7), .A2(n_137), .B1(n_291), .B2(n_296), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_8), .A2(n_77), .B1(n_285), .B2(n_307), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_9), .A2(n_93), .B1(n_293), .B2(n_619), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_11), .A2(n_46), .B1(n_435), .B2(n_436), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_12), .A2(n_179), .B1(n_497), .B2(n_498), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_13), .Y(n_355) );
XOR2x2_ASAP7_75t_L g538 ( .A(n_14), .B(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_15), .A2(n_219), .B1(n_318), .B2(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_16), .A2(n_68), .B1(n_460), .B2(n_605), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_17), .Y(n_712) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_18), .A2(n_60), .B1(n_246), .B2(n_251), .Y(n_255) );
INVx1_ASAP7_75t_L g651 ( .A(n_18), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_19), .A2(n_121), .B1(n_241), .B2(n_256), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_20), .A2(n_23), .B1(n_337), .B2(n_422), .Y(n_489) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_21), .A2(n_76), .B1(n_96), .B2(n_411), .C1(n_476), .C2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_22), .A2(n_185), .B1(n_348), .B2(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g632 ( .A(n_24), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g299 ( .A1(n_25), .A2(n_67), .B1(n_201), .B2(n_300), .C1(n_303), .C2(n_306), .Y(n_299) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_26), .A2(n_45), .B1(n_318), .B2(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_27), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_28), .A2(n_124), .B1(n_423), .B2(n_465), .Y(n_572) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_29), .A2(n_63), .B1(n_246), .B2(n_247), .Y(n_253) );
INVx1_ASAP7_75t_L g652 ( .A(n_29), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_30), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_31), .A2(n_33), .B1(n_368), .B2(n_558), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_32), .A2(n_89), .B1(n_332), .B2(n_348), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_34), .A2(n_212), .B1(n_411), .B2(n_588), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_35), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_36), .A2(n_116), .B1(n_435), .B2(n_436), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_37), .B(n_321), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_38), .A2(n_186), .B1(n_453), .B2(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_39), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_40), .A2(n_90), .B1(n_432), .B2(n_433), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_41), .A2(n_161), .B1(n_436), .B2(n_452), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_42), .Y(n_726) );
XOR2x2_ASAP7_75t_L g595 ( .A(n_43), .B(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_44), .A2(n_166), .B1(n_351), .B2(n_352), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_47), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_48), .B(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_49), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_50), .A2(n_66), .B1(n_427), .B2(n_429), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_51), .B(n_457), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_52), .A2(n_127), .B1(n_523), .B2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g395 ( .A(n_53), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_54), .A2(n_146), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g316 ( .A1(n_55), .A2(n_119), .B1(n_317), .B2(n_318), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_56), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_57), .A2(n_88), .B1(n_262), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_58), .A2(n_206), .B1(n_486), .B2(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_59), .A2(n_213), .B1(n_273), .B2(n_278), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_61), .A2(n_655), .B1(n_687), .B2(n_688), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_61), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_62), .A2(n_114), .B1(n_325), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_64), .A2(n_209), .B1(n_262), .B2(n_267), .Y(n_261) );
AOI22xp33_ASAP7_75t_SL g328 ( .A1(n_65), .A2(n_169), .B1(n_256), .B2(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g230 ( .A(n_69), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_70), .A2(n_97), .B1(n_348), .B2(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_71), .B(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_72), .Y(n_481) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_73), .A2(n_147), .B1(n_293), .B2(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_74), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g226 ( .A(n_75), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_78), .A2(n_211), .B1(n_293), .B2(n_349), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_79), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_80), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_81), .A2(n_136), .B1(n_296), .B2(n_298), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_82), .A2(n_154), .B1(n_523), .B2(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_83), .A2(n_92), .B1(n_291), .B2(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g634 ( .A(n_84), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_85), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_86), .B(n_414), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_87), .A2(n_98), .B1(n_173), .B2(n_385), .C1(n_684), .C2(n_686), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_91), .Y(n_670) );
INVx1_ASAP7_75t_L g628 ( .A(n_94), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_95), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_99), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_100), .A2(n_200), .B1(n_491), .B2(n_493), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_101), .A2(n_104), .B1(n_449), .B2(n_619), .Y(n_618) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_102), .A2(n_223), .B(n_231), .C(n_653), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_103), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_105), .A2(n_133), .B1(n_452), .B2(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_106), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g630 ( .A(n_107), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g635 ( .A1(n_108), .A2(n_144), .B1(n_151), .B2(n_280), .C1(n_301), .C2(n_414), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g468 ( .A1(n_109), .A2(n_138), .B1(n_168), .B2(n_301), .C1(n_325), .C2(n_469), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_110), .A2(n_198), .B1(n_385), .B2(n_518), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_111), .A2(n_160), .B1(n_560), .B2(n_562), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_112), .A2(n_221), .B1(n_456), .B2(n_487), .C(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_113), .A2(n_216), .B1(n_436), .B2(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g698 ( .A(n_115), .Y(n_698) );
AOI22xp5_ASAP7_75t_SL g701 ( .A1(n_115), .A2(n_698), .B1(n_702), .B2(n_729), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_117), .A2(n_148), .B1(n_531), .B2(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_L g229 ( .A(n_118), .B(n_230), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_120), .A2(n_191), .B1(n_317), .B2(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_122), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_123), .A2(n_204), .B1(n_574), .B2(n_575), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_125), .A2(n_192), .B1(n_318), .B2(n_460), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_126), .A2(n_175), .B1(n_429), .B2(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_128), .Y(n_705) );
AND2x6_ASAP7_75t_L g225 ( .A(n_129), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_129), .Y(n_645) );
AO22x2_ASAP7_75t_L g245 ( .A1(n_130), .A2(n_183), .B1(n_246), .B2(n_247), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_131), .A2(n_210), .B1(n_453), .B2(n_565), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_132), .A2(n_163), .B1(n_414), .B2(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g338 ( .A(n_134), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_135), .B(n_273), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_139), .A2(n_205), .B1(n_527), .B2(n_528), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_140), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_141), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_142), .A2(n_215), .B1(n_464), .B2(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g622 ( .A(n_143), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_145), .Y(n_590) );
INVx1_ASAP7_75t_L g636 ( .A(n_149), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_150), .A2(n_177), .B1(n_267), .B2(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_152), .B(n_323), .Y(n_322) );
AO22x2_ASAP7_75t_L g250 ( .A1(n_153), .A2(n_193), .B1(n_246), .B2(n_251), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_155), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_156), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_157), .B(n_457), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_158), .Y(n_416) );
XOR2x2_ASAP7_75t_L g445 ( .A(n_159), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_162), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_164), .A2(n_199), .B1(n_306), .B2(n_460), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_165), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_167), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_170), .B(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g324 ( .A1(n_171), .A2(n_217), .B1(n_286), .B2(n_325), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_172), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_174), .A2(n_214), .B1(n_241), .B2(n_612), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_176), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_178), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_180), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_181), .Y(n_708) );
XOR2x2_ASAP7_75t_L g504 ( .A(n_182), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_183), .B(n_650), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_184), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_187), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_188), .A2(n_195), .B1(n_429), .B2(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_189), .Y(n_680) );
INVx1_ASAP7_75t_L g648 ( .A(n_193), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_194), .A2(n_218), .B1(n_456), .B2(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g508 ( .A(n_196), .Y(n_508) );
OA22x2_ASAP7_75t_L g470 ( .A1(n_197), .A2(n_471), .B1(n_472), .B2(n_500), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_197), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_202), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_203), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_207), .Y(n_402) );
INVx1_ASAP7_75t_L g246 ( .A(n_208), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_220), .B(n_273), .Y(n_603) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_226), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_227), .A2(n_643), .B(n_697), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_534), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_231) );
INVx1_ASAP7_75t_L g638 ( .A(n_232), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_441), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B1(n_340), .B2(n_440), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AO22x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_310), .B2(n_339), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
XOR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_309), .Y(n_237) );
NAND4xp75_ASAP7_75t_L g238 ( .A(n_239), .B(n_271), .C(n_289), .D(n_299), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_261), .Y(n_239) );
BUFx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx3_ASAP7_75t_L g337 ( .A(n_242), .Y(n_337) );
INVx6_ASAP7_75t_L g358 ( .A(n_242), .Y(n_358) );
BUFx3_ASAP7_75t_L g586 ( .A(n_242), .Y(n_586) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
AND2x2_ASAP7_75t_L g297 ( .A(n_243), .B(n_264), .Y(n_297) );
AND2x6_ASAP7_75t_L g298 ( .A(n_243), .B(n_276), .Y(n_298) );
AND2x6_ASAP7_75t_L g301 ( .A(n_243), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_249), .Y(n_243) );
AND2x2_ASAP7_75t_L g266 ( .A(n_244), .B(n_250), .Y(n_266) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g259 ( .A(n_245), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_245), .B(n_250), .Y(n_270) );
AND2x2_ASAP7_75t_L g284 ( .A(n_245), .B(n_255), .Y(n_284) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g251 ( .A(n_248), .Y(n_251) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g260 ( .A(n_250), .Y(n_260) );
INVx1_ASAP7_75t_L g283 ( .A(n_250), .Y(n_283) );
AND2x2_ASAP7_75t_L g258 ( .A(n_252), .B(n_259), .Y(n_258) );
AND2x6_ASAP7_75t_L g278 ( .A(n_252), .B(n_266), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_252), .B(n_266), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_252), .B(n_259), .Y(n_665) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g265 ( .A(n_253), .Y(n_265) );
OR2x2_ASAP7_75t_L g277 ( .A(n_253), .B(n_254), .Y(n_277) );
INVx1_ASAP7_75t_L g288 ( .A(n_253), .Y(n_288) );
AND2x2_ASAP7_75t_L g302 ( .A(n_253), .B(n_255), .Y(n_302) );
AND2x2_ASAP7_75t_L g264 ( .A(n_254), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx2_ASAP7_75t_L g435 ( .A(n_256), .Y(n_435) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_256), .Y(n_452) );
INVx5_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g351 ( .A(n_257), .Y(n_351) );
INVx1_ASAP7_75t_L g492 ( .A(n_257), .Y(n_492) );
BUFx3_ASAP7_75t_L g566 ( .A(n_257), .Y(n_566) );
INVx3_ASAP7_75t_L g574 ( .A(n_257), .Y(n_574) );
INVx4_ASAP7_75t_L g720 ( .A(n_257), .Y(n_720) );
INVx8_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g292 ( .A(n_259), .B(n_264), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_259), .B(n_264), .Y(n_362) );
INVx1_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
INVx4_ASAP7_75t_L g365 ( .A(n_262), .Y(n_365) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g333 ( .A(n_263), .Y(n_333) );
BUFx3_ASAP7_75t_L g433 ( .A(n_263), .Y(n_433) );
BUFx3_ASAP7_75t_L g568 ( .A(n_263), .Y(n_568) );
BUFx3_ASAP7_75t_L g584 ( .A(n_263), .Y(n_584) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x4_ASAP7_75t_L g294 ( .A(n_264), .B(n_269), .Y(n_294) );
INVx1_ASAP7_75t_L g268 ( .A(n_265), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_265), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g275 ( .A(n_266), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g390 ( .A(n_266), .Y(n_390) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_268), .B(n_284), .Y(n_374) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x6_ASAP7_75t_L g353 ( .A(n_270), .B(n_288), .Y(n_353) );
AND2x2_ASAP7_75t_SL g271 ( .A(n_272), .B(n_279), .Y(n_271) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_273), .Y(n_456) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_273), .Y(n_550) );
INVx5_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g321 ( .A(n_274), .Y(n_321) );
INVx2_ASAP7_75t_L g486 ( .A(n_274), .Y(n_486) );
INVx2_ASAP7_75t_L g516 ( .A(n_274), .Y(n_516) );
INVx4_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g389 ( .A(n_277), .B(n_390), .Y(n_389) );
BUFx4f_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
INVx1_ASAP7_75t_SL g458 ( .A(n_278), .Y(n_458) );
BUFx2_ASAP7_75t_L g487 ( .A(n_278), .Y(n_487) );
BUFx2_ASAP7_75t_L g552 ( .A(n_278), .Y(n_552) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_280), .Y(n_411) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx4f_ASAP7_75t_SL g325 ( .A(n_281), .Y(n_325) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_281), .Y(n_385) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_281), .Y(n_512) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g305 ( .A(n_283), .Y(n_305) );
AND2x4_ASAP7_75t_L g286 ( .A(n_284), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g304 ( .A(n_284), .B(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g461 ( .A(n_286), .Y(n_461) );
BUFx2_ASAP7_75t_L g484 ( .A(n_286), .Y(n_484) );
BUFx2_ASAP7_75t_L g518 ( .A(n_286), .Y(n_518) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_295), .Y(n_289) );
INVx1_ASAP7_75t_L g529 ( .A(n_291), .Y(n_529) );
BUFx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g423 ( .A(n_292), .Y(n_423) );
BUFx3_ASAP7_75t_L g464 ( .A(n_292), .Y(n_464) );
BUFx3_ASAP7_75t_L g558 ( .A(n_292), .Y(n_558) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_SL g368 ( .A(n_294), .Y(n_368) );
BUFx3_ASAP7_75t_L g425 ( .A(n_294), .Y(n_425) );
BUFx3_ASAP7_75t_L g465 ( .A(n_294), .Y(n_465) );
BUFx2_ASAP7_75t_SL g532 ( .A(n_294), .Y(n_532) );
BUFx3_ASAP7_75t_L g562 ( .A(n_294), .Y(n_562) );
BUFx3_ASAP7_75t_L g432 ( .A(n_296), .Y(n_432) );
BUFx3_ASAP7_75t_L g497 ( .A(n_296), .Y(n_497) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_296), .Y(n_527) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_SL g348 ( .A(n_297), .Y(n_348) );
BUFx2_ASAP7_75t_SL g449 ( .A(n_297), .Y(n_449) );
INVx2_ASAP7_75t_L g561 ( .A(n_297), .Y(n_561) );
INVx11_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
INVx11_ASAP7_75t_L g428 ( .A(n_298), .Y(n_428) );
BUFx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g314 ( .A(n_301), .Y(n_314) );
INVx4_ASAP7_75t_L g380 ( .A(n_301), .Y(n_380) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_301), .Y(n_408) );
INVx2_ASAP7_75t_SL g542 ( .A(n_301), .Y(n_542) );
AND2x4_ASAP7_75t_L g307 ( .A(n_302), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g377 ( .A(n_302), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g469 ( .A(n_303), .Y(n_469) );
INVx2_ASAP7_75t_L g589 ( .A(n_303), .Y(n_589) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_304), .Y(n_317) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_304), .Y(n_414) );
BUFx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_SL g318 ( .A(n_307), .Y(n_318) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_307), .Y(n_547) );
BUFx2_ASAP7_75t_SL g605 ( .A(n_307), .Y(n_605) );
INVx1_ASAP7_75t_L g378 ( .A(n_308), .Y(n_378) );
INVx2_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
XOR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_338), .Y(n_310) );
NAND2x1_ASAP7_75t_L g311 ( .A(n_312), .B(n_326), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_319), .Y(n_312) );
OAI21xp5_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_315), .B(n_316), .Y(n_313) );
INVx2_ASAP7_75t_L g382 ( .A(n_317), .Y(n_382) );
BUFx3_ASAP7_75t_L g686 ( .A(n_317), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .C(n_324), .Y(n_319) );
INVx1_ASAP7_75t_L g478 ( .A(n_325), .Y(n_478) );
NOR2x1_ASAP7_75t_L g326 ( .A(n_327), .B(n_334), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx4_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g349 ( .A(n_330), .Y(n_349) );
INVx2_ASAP7_75t_SL g612 ( .A(n_330), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_330), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g440 ( .A(n_340), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_396), .B2(n_397), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
XOR2xp5_ASAP7_75t_SL g343 ( .A(n_344), .B(n_395), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_369), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_354), .C(n_363), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_350), .Y(n_346) );
INVx1_ASAP7_75t_L g727 ( .A(n_348), .Y(n_727) );
INVx1_ASAP7_75t_L g633 ( .A(n_349), .Y(n_633) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx6_ASAP7_75t_SL g437 ( .A(n_353), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_359), .B2(n_360), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_356), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g429 ( .A(n_358), .Y(n_429) );
INVx2_ASAP7_75t_L g531 ( .A(n_358), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_358), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_360), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g675 ( .A(n_361), .Y(n_675) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_366), .B2(n_367), .Y(n_363) );
INVx4_ASAP7_75t_L g450 ( .A(n_365), .Y(n_450) );
INVx3_ASAP7_75t_L g619 ( .A(n_365), .Y(n_619) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NOR3xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_379), .C(n_386), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_375), .B2(n_376), .Y(n_370) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_372), .A2(n_418), .B1(n_712), .B2(n_713), .Y(n_711) );
INVx3_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx4_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_374), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_415) );
BUFx3_ASAP7_75t_L g681 ( .A(n_374), .Y(n_681) );
BUFx2_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
OR2x6_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_382), .B2(n_383), .C(n_384), .Y(n_379) );
INVx4_ASAP7_75t_L g476 ( .A(n_380), .Y(n_476) );
BUFx2_ASAP7_75t_L g685 ( .A(n_380), .Y(n_685) );
OAI21xp5_ASAP7_75t_SL g707 ( .A1(n_380), .A2(n_708), .B(n_709), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_391), .B2(n_392), .Y(n_386) );
BUFx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_389), .Y(n_403) );
OAI22xp5_ASAP7_75t_SL g704 ( .A1(n_389), .A2(n_579), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g405 ( .A(n_393), .Y(n_405) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx3_ASAP7_75t_L g579 ( .A(n_394), .Y(n_579) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_419), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_406), .C(n_415), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B1(n_410), .B2(n_412), .C(n_413), .Y(n_406) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_407), .A2(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g480 ( .A(n_414), .Y(n_480) );
BUFx4f_ASAP7_75t_L g710 ( .A(n_414), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_418), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_430), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_426), .Y(n_420) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g677 ( .A(n_424), .Y(n_677) );
BUFx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g723 ( .A(n_427), .Y(n_723) );
INVx4_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g467 ( .A(n_428), .Y(n_467) );
INVx2_ASAP7_75t_SL g523 ( .A(n_428), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g499 ( .A(n_433), .Y(n_499) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g453 ( .A(n_437), .Y(n_453) );
BUFx2_ASAP7_75t_L g493 ( .A(n_437), .Y(n_493) );
BUFx2_ASAP7_75t_L g575 ( .A(n_437), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_443), .B1(n_502), .B2(n_533), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_470), .B2(n_501), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND4xp75_ASAP7_75t_L g446 ( .A(n_447), .B(n_454), .C(n_462), .D(n_468), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
AND2x2_ASAP7_75t_SL g454 ( .A(n_455), .B(n_459), .Y(n_454) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .Y(n_462) );
INVxp67_ASAP7_75t_L g629 ( .A(n_465), .Y(n_629) );
INVx1_ASAP7_75t_L g501 ( .A(n_470), .Y(n_501) );
INVx2_ASAP7_75t_L g500 ( .A(n_472), .Y(n_500) );
NAND3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_488), .C(n_494), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
OAI222xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B1(n_478), .B2(n_479), .C1(n_480), .C2(n_481), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g507 ( .A1(n_475), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
BUFx2_ASAP7_75t_L g624 ( .A(n_486), .Y(n_624) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_L g667 ( .A(n_493), .Y(n_667) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g533 ( .A(n_502), .Y(n_533) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND3x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_519), .C(n_525), .Y(n_505) );
NOR2x1_ASAP7_75t_SL g506 ( .A(n_507), .B(n_513), .Y(n_506) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .C(n_517), .Y(n_513) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g639 ( .A(n_534), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_593), .B2(n_594), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AO22x2_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_569), .B1(n_591), .B2(n_592), .Y(n_537) );
INVx2_ASAP7_75t_L g591 ( .A(n_538), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_554), .Y(n_539) );
NOR2xp33_ASAP7_75t_SL g540 ( .A(n_541), .B(n_548), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_543), .B(n_544), .Y(n_541) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .C(n_553), .Y(n_548) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_563), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
BUFx4f_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_561), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx3_ASAP7_75t_SL g592 ( .A(n_569), .Y(n_592) );
XOR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_590), .Y(n_569) );
NAND4xp75_ASAP7_75t_L g570 ( .A(n_571), .B(n_576), .C(n_582), .D(n_587), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OA211x2_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_580), .C(n_581), .Y(n_576) );
OA211x2_ASAP7_75t_L g621 ( .A1(n_578), .A2(n_622), .B(n_623), .C(n_625), .Y(n_621) );
BUFx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
BUFx2_ASAP7_75t_L g661 ( .A(n_584), .Y(n_661) );
INVx1_ASAP7_75t_L g672 ( .A(n_586), .Y(n_672) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI22xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_613), .B1(n_614), .B2(n_637), .Y(n_594) );
INVx1_ASAP7_75t_L g637 ( .A(n_595), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_606), .C(n_609), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .C(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
XOR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_636), .Y(n_615) );
NAND4xp75_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .C(n_626), .D(n_635), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .Y(n_626) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_646), .Y(n_641) );
OR2x2_ASAP7_75t_SL g732 ( .A(n_642), .B(n_647), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_643), .Y(n_690) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_644), .B(n_694), .Y(n_697) );
CKINVDCx16_ASAP7_75t_R g694 ( .A(n_645), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
OAI322xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_689), .A3(n_691), .B1(n_695), .B2(n_698), .C1(n_699), .C2(n_730), .Y(n_653) );
INVx1_ASAP7_75t_L g688 ( .A(n_655), .Y(n_688) );
AND4x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_668), .C(n_678), .D(n_683), .Y(n_655) );
NOR2xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_662), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_666), .B2(n_667), .Y(n_662) );
BUFx2_ASAP7_75t_R g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_SL g668 ( .A(n_669), .B(n_673), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_675), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g729 ( .A(n_702), .Y(n_729) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_714), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .C(n_711), .Y(n_703) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_721), .C(n_725), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
endmodule