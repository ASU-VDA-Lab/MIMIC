module fake_jpeg_127_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_67),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_49),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_1),
.C(n_2),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_42),
.B(n_36),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_23),
.Y(n_89)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_54),
.Y(n_110)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_4),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_73),
.B(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_79),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_80),
.Y(n_102)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_82),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_41),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_89),
.B(n_92),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_40),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_72),
.B(n_109),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_44),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_109),
.B1(n_120),
.B2(n_122),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_113),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_28),
.B1(n_27),
.B2(n_37),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_19),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_111),
.B(n_125),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_28),
.B1(n_38),
.B2(n_37),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_115),
.B1(n_64),
.B2(n_60),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_23),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_36),
.B1(n_34),
.B2(n_6),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_10),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_34),
.B1(n_5),
.B2(n_7),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_5),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_62),
.A2(n_9),
.B1(n_11),
.B2(n_79),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_92),
.B1(n_126),
.B2(n_121),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_68),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_133),
.C(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_137),
.B1(n_141),
.B2(n_147),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_135),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_117),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_90),
.B1(n_104),
.B2(n_124),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_157),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_94),
.B1(n_96),
.B2(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_156),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_95),
.B1(n_96),
.B2(n_112),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_160),
.B1(n_130),
.B2(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_153),
.Y(n_170)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_123),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_90),
.A2(n_84),
.B1(n_97),
.B2(n_100),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_162),
.B(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_118),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_149),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_116),
.B1(n_97),
.B2(n_100),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_112),
.B1(n_115),
.B2(n_102),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_102),
.B1(n_51),
.B2(n_49),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_145),
.B(n_147),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_181),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_178),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_142),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_140),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_171),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_179),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_141),
.B1(n_159),
.B2(n_144),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_190),
.B1(n_173),
.B2(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_159),
.B1(n_138),
.B2(n_136),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_148),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

AOI22x1_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_152),
.B1(n_159),
.B2(n_178),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_200),
.B(n_201),
.Y(n_205)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_198),
.B(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_159),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_176),
.B(n_169),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_196),
.B(n_194),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_177),
.C(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_206),
.C(n_215),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_190),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_174),
.B1(n_173),
.B2(n_180),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_182),
.B1(n_170),
.B2(n_180),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_213),
.A2(n_198),
.B(n_186),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_186),
.C(n_197),
.Y(n_215)
);

XNOR2x2_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_225),
.B1(n_210),
.B2(n_191),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_209),
.B(n_211),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_221),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_196),
.C(n_183),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_226),
.C(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_192),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_213),
.C(n_203),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_218),
.B(n_211),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_217),
.B1(n_226),
.B2(n_219),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_233),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_205),
.C(n_209),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_211),
.B(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_230),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_244),
.B(n_240),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_247),
.B(n_243),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_230),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_214),
.CI(n_201),
.CON(n_249),
.SN(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_214),
.C(n_195),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_200),
.B1(n_189),
.B2(n_185),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_250),
.Y(n_253)
);


endmodule