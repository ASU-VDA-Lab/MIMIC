module fake_jpeg_26735_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_25),
.B1(n_17),
.B2(n_22),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_27),
.B1(n_29),
.B2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_15),
.B(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_38),
.B1(n_17),
.B2(n_40),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_73),
.B1(n_74),
.B2(n_23),
.Y(n_109)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2x1_ASAP7_75t_R g62 ( 
.A(n_44),
.B(n_16),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_34),
.B1(n_54),
.B2(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_38),
.B1(n_17),
.B2(n_34),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_34),
.B1(n_32),
.B2(n_24),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_24),
.B1(n_18),
.B2(n_26),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_54),
.B1(n_16),
.B2(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_95),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_98),
.B1(n_65),
.B2(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_39),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_39),
.C(n_36),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_101),
.C(n_23),
.Y(n_140)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_107),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_53),
.B1(n_57),
.B2(n_82),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_79),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_106),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_80),
.B1(n_75),
.B2(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_19),
.B1(n_28),
.B2(n_16),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_36),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_112),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_77),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_114),
.A2(n_91),
.B(n_1),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_69),
.B1(n_68),
.B2(n_58),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_134),
.B1(n_100),
.B2(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_122),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_68),
.B(n_69),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_119),
.B(n_128),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_70),
.B1(n_76),
.B2(n_65),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_99),
.B1(n_102),
.B2(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_14),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_14),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_28),
.B(n_19),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_137),
.B(n_0),
.Y(n_169)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_133),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_36),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_99),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_36),
.B1(n_21),
.B2(n_23),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_93),
.B1(n_90),
.B2(n_99),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_114),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_19),
.B(n_31),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_31),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_112),
.B(n_90),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_96),
.C(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_140),
.C(n_119),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_149),
.B1(n_173),
.B2(n_133),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_94),
.B1(n_95),
.B2(n_86),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_153),
.B1(n_165),
.B2(n_166),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_156),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_155),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_152),
.B(n_169),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_159),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_0),
.B(n_1),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_100),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_23),
.A3(n_21),
.B1(n_91),
.B2(n_14),
.C1(n_12),
.C2(n_5),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_21),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_138),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_91),
.B1(n_1),
.B2(n_2),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_91),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_189),
.C(n_169),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_140),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_184),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_171),
.A2(n_131),
.B1(n_129),
.B2(n_119),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_183),
.B1(n_190),
.B2(n_193),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_173),
.B1(n_170),
.B2(n_162),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_120),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_187),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_123),
.C(n_137),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_123),
.B1(n_122),
.B2(n_116),
.Y(n_190)
);

AOI22x1_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_138),
.B1(n_125),
.B2(n_134),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_124),
.B1(n_130),
.B2(n_139),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_202),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_149),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_2),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_4),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_206),
.C(n_207),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_168),
.C(n_159),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_168),
.C(n_148),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_167),
.C(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_212),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_152),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_164),
.C(n_158),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_147),
.B(n_4),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_191),
.B(n_186),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_3),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_224),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_174),
.B(n_4),
.CI(n_6),
.CON(n_222),
.SN(n_222)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_225),
.A2(n_177),
.B1(n_208),
.B2(n_214),
.Y(n_234)
);

FAx1_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_191),
.CI(n_210),
.CON(n_229),
.SN(n_229)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_229),
.A2(n_243),
.B1(n_230),
.B2(n_228),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_175),
.B1(n_194),
.B2(n_182),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_188),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_239),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_194),
.B1(n_186),
.B2(n_225),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_188),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_195),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_201),
.B(n_177),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_240),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_217),
.C(n_216),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_252),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_217),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_235),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_201),
.B1(n_215),
.B2(n_205),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_254),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_246),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_226),
.C(n_211),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_200),
.B1(n_185),
.B2(n_222),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_257),
.Y(n_271)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_229),
.B1(n_239),
.B2(n_222),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_231),
.C(n_229),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_247),
.C(n_250),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_199),
.B1(n_220),
.B2(n_221),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_235),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_275),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_224),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_278),
.B1(n_273),
.B2(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_254),
.C(n_260),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_6),
.C(n_7),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_258),
.C(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_285),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_6),
.C(n_7),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_292),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_271),
.B1(n_266),
.B2(n_8),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_10),
.B1(n_11),
.B2(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_6),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_280),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_7),
.B(n_8),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_9),
.B(n_10),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_293),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_296),
.C(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_301),
.B(n_298),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_302),
.C(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_291),
.C(n_297),
.Y(n_307)
);

NAND4xp25_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_290),
.C(n_10),
.D(n_11),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_11),
.B(n_211),
.Y(n_309)
);


endmodule