module fake_ibex_626_n_2615 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_407, n_102, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_460, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2615);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_407;
input n_102;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_460;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2615;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2475;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_641;
wire n_557;
wire n_2311;
wire n_1937;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_787;
wire n_523;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_709;
wire n_499;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2509;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_737;
wire n_606;
wire n_2445;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2470;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2424;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2252;
wire n_1982;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_2590;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_2484;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2524;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_1331;
wire n_634;
wire n_1349;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_1340;
wire n_2562;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1839;
wire n_1617;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2611;
wire n_1538;
wire n_487;
wire n_2528;
wire n_2548;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_484;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_1362;
wire n_707;
wire n_1586;
wire n_1097;
wire n_2518;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_645;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2487;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1385;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_704;
wire n_2357;
wire n_2104;
wire n_924;
wire n_2331;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_2430;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

BUFx10_ASAP7_75t_L g467 ( 
.A(n_365),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_214),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_335),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_164),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_144),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_55),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_6),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_328),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_58),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_426),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_36),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_83),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_164),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_181),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_226),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_290),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_388),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_80),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_132),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_376),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_196),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_75),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_120),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_246),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_229),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_451),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_26),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_308),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_424),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_341),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_318),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_35),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_217),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_337),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_316),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_105),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_34),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_198),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_423),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_44),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_61),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_286),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_303),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_84),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_41),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_393),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_296),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_360),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_19),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_272),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_455),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_332),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_223),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_357),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_383),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_97),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_79),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_117),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_154),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_325),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_275),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_226),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_329),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_199),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_183),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_179),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_162),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_359),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_373),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_179),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_218),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_389),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_261),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_47),
.Y(n_544)
);

BUFx5_ASAP7_75t_L g545 ( 
.A(n_66),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_285),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_155),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_95),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_183),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_103),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_139),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_213),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_322),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_149),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_380),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_284),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_22),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_76),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_188),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_338),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_465),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_43),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_21),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_174),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_137),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_244),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_219),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_199),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_76),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_448),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_366),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_31),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_347),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_402),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_429),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_409),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_92),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_234),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_282),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_412),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_297),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_215),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_432),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_342),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_125),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_82),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_410),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_34),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_407),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_81),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_364),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_30),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_385),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_441),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_281),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_10),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_343),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_127),
.Y(n_600)
);

CKINVDCx14_ASAP7_75t_R g601 ( 
.A(n_422),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_382),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_168),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_461),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_390),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_54),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_21),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_370),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_438),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_149),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_300),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_36),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_5),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_94),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_334),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_163),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_252),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_458),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_295),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_27),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_98),
.Y(n_621)
);

CKINVDCx14_ASAP7_75t_R g622 ( 
.A(n_259),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_330),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_243),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_119),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_278),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_299),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_114),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_387),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_134),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_175),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_350),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_16),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_411),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_2),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_456),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_79),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_430),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_192),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_344),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_356),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_6),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_225),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_257),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_449),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_240),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_395),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_354),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_440),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_120),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_425),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_118),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_408),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_123),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_102),
.Y(n_655)
);

CKINVDCx14_ASAP7_75t_R g656 ( 
.A(n_362),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_113),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_443),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_206),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_250),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_87),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_55),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_283),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_309),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_435),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_258),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_67),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_406),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_457),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_302),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_3),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_154),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_225),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_401),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_44),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_415),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_170),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_294),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_100),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_363),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_320),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_403),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_452),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_127),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_136),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_185),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_258),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_156),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_73),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_119),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_84),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_229),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_236),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_391),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_419),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_287),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_278),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_8),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_47),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_118),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_117),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_78),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_353),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_289),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_340),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_396),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_405),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_349),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_352),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_459),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_135),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_445),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_301),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_420),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_3),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_112),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_195),
.Y(n_717)
);

BUFx10_ASAP7_75t_L g718 ( 
.A(n_367),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_235),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_305),
.Y(n_720)
);

BUFx10_ASAP7_75t_L g721 ( 
.A(n_273),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_450),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_454),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_94),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_205),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_291),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_428),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_142),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_319),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_169),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_186),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_221),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_163),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_146),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_227),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_123),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_355),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_151),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_386),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_377),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_134),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_126),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_314),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_273),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_87),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_90),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_22),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_346),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_250),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_37),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_361),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_321),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_222),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_170),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_1),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_327),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_394),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_392),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_217),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_311),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_60),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_172),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_444),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_184),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_64),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_381),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_351),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_77),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_90),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_27),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_184),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_336),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_167),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_133),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_23),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_358),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_169),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_15),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_166),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_464),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_339),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_158),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_31),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_213),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_201),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_103),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_472),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_571),
.B(n_0),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_674),
.Y(n_789)
);

XNOR2xp5_ASAP7_75t_L g790 ( 
.A(n_482),
.B(n_0),
.Y(n_790)
);

INVxp33_ASAP7_75t_SL g791 ( 
.A(n_683),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_545),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_609),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_662),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_662),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_692),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_487),
.Y(n_797)
);

BUFx2_ASAP7_75t_SL g798 ( 
.A(n_487),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_504),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_499),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_499),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_504),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_539),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_505),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_622),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_527),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_601),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_482),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_660),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_534),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_539),
.Y(n_811)
);

CKINVDCx16_ASAP7_75t_R g812 ( 
.A(n_534),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_687),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_527),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_551),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_545),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_608),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_551),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_592),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_608),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_619),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_765),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_592),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_632),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_594),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_473),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_632),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_594),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_553),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_489),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_649),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_489),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_529),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_627),
.B(n_1),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_553),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_529),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_536),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_536),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_537),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_537),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_649),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_544),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_568),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_568),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_651),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_471),
.B(n_2),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_569),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_544),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_559),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_569),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_559),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_545),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_570),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_651),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_480),
.B(n_4),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_570),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_579),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_579),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_696),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_696),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_623),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_590),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_590),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_625),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_643),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_625),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_534),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_631),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_643),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_703),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_703),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_661),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_627),
.B(n_4),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_473),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_656),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_631),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_661),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_704),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_679),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_704),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_742),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_721),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_644),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_644),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_742),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_647),
.B(n_5),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_768),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_545),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_714),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_545),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_545),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_545),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_714),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_623),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_720),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_533),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_479),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_481),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_491),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_659),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_721),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_506),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_659),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_506),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_647),
.B(n_7),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_720),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_721),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_492),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_509),
.B(n_8),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_689),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_508),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_533),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_640),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_757),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_512),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_794),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_795),
.B(n_528),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_791),
.A2(n_513),
.B1(n_519),
.B2(n_508),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_792),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_792),
.A2(n_549),
.B(n_538),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_816),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_816),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_852),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_813),
.B(n_796),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_R g925 ( 
.A(n_791),
.B(n_513),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_852),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_888),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_822),
.B(n_467),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_890),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_808),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_806),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_789),
.B(n_682),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_799),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_809),
.B(n_467),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_787),
.B(n_682),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_896),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_892),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_802),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_896),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_804),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_897),
.B(n_535),
.Y(n_941)
);

OA21x2_ASAP7_75t_L g942 ( 
.A1(n_891),
.A2(n_549),
.B(n_538),
.Y(n_942)
);

OA21x2_ASAP7_75t_L g943 ( 
.A1(n_886),
.A2(n_638),
.B(n_602),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_904),
.B(n_467),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_912),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_912),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_858),
.B(n_540),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_819),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_823),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_826),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_814),
.B(n_730),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_825),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_828),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_861),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_894),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_877),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_807),
.B(n_757),
.Y(n_957)
);

CKINVDCx8_ASAP7_75t_R g958 ( 
.A(n_798),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_898),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_894),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_805),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_913),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_899),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_SL g964 ( 
.A1(n_808),
.A2(n_719),
.B1(n_733),
.B2(n_689),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_810),
.B(n_476),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_913),
.B(n_731),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_830),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_832),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_874),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_902),
.Y(n_970)
);

BUFx8_ASAP7_75t_L g971 ( 
.A(n_846),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_833),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_915),
.B(n_543),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_836),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_837),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_838),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_812),
.B(n_476),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_839),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_840),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_842),
.Y(n_980)
);

NAND2x1_ASAP7_75t_L g981 ( 
.A(n_788),
.B(n_469),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_848),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_849),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_851),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_853),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_867),
.B(n_882),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_856),
.Y(n_987)
);

BUFx8_ASAP7_75t_L g988 ( 
.A(n_857),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_911),
.A2(n_734),
.B1(n_738),
.B2(n_731),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_865),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_908),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_807),
.B(n_734),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_869),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_SL g994 ( 
.A(n_875),
.B(n_474),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_872),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_879),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_834),
.B(n_602),
.Y(n_997)
);

CKINVDCx6p67_ASAP7_75t_R g998 ( 
.A(n_815),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_881),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_875),
.B(n_901),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_885),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_887),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_805),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_873),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_905),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_909),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_907),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_855),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_793),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_790),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_878),
.A2(n_680),
.B(n_638),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_880),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_880),
.B(n_680),
.Y(n_1013)
);

OA21x2_ASAP7_75t_L g1014 ( 
.A1(n_797),
.A2(n_510),
.B(n_497),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_800),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_801),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_803),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_811),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_817),
.A2(n_521),
.B(n_516),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_820),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_821),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_824),
.A2(n_526),
.B(n_524),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_827),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_831),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_841),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_845),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_854),
.B(n_554),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_859),
.B(n_572),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_860),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_870),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_914),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_871),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_889),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_893),
.B(n_495),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_895),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_906),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_910),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_910),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_815),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_818),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_903),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_829),
.B(n_749),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_835),
.A2(n_582),
.B(n_577),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_903),
.B(n_548),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_835),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_900),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_843),
.B(n_783),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_900),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_843),
.Y(n_1049)
);

XOR2xp5_ASAP7_75t_L g1050 ( 
.A(n_844),
.B(n_847),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_844),
.B(n_586),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_847),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_884),
.B(n_565),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_884),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_850),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_850),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_883),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_862),
.A2(n_591),
.B(n_589),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_883),
.B(n_574),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_862),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_876),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_876),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_863),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_863),
.B(n_783),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_868),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_864),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_864),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_866),
.Y(n_1068)
);

BUFx8_ASAP7_75t_L g1069 ( 
.A(n_866),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_868),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_792),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_806),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_792),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_904),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_794),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_792),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_794),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_794),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_806),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_794),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_794),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_794),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_806),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_791),
.B(n_511),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_794),
.B(n_584),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_794),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_794),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_794),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_792),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_904),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_792),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_792),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_792),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_794),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_792),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_813),
.B(n_476),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_794),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_792),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_794),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_904),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_813),
.B(n_503),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_904),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_792),
.Y(n_1103)
);

XNOR2xp5_ASAP7_75t_L g1104 ( 
.A(n_808),
.B(n_719),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_794),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_794),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_813),
.B(n_503),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_791),
.A2(n_470),
.B1(n_475),
.B2(n_468),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_792),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_904),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_806),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_792),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_792),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_794),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_806),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_794),
.Y(n_1116)
);

AND2x6_ASAP7_75t_L g1117 ( 
.A(n_965),
.B(n_640),
.Y(n_1117)
);

OR2x2_ASAP7_75t_SL g1118 ( 
.A(n_1049),
.B(n_733),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_986),
.B(n_588),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_916),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1074),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_991),
.B(n_478),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1004),
.B(n_593),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_991),
.B(n_514),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1007),
.B(n_771),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_988),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_955),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_973),
.B(n_514),
.Y(n_1128)
);

AO22x2_ASAP7_75t_L g1129 ( 
.A1(n_1051),
.A2(n_607),
.B1(n_614),
.B2(n_603),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1075),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1005),
.B(n_503),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1077),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1078),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1007),
.B(n_718),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_973),
.B(n_515),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1090),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1115),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1080),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_955),
.Y(n_1139)
);

OR2x2_ASAP7_75t_SL g1140 ( 
.A(n_1049),
.B(n_736),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_988),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_955),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_930),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_924),
.B(n_518),
.Y(n_1144)
);

INVx4_ASAP7_75t_SL g1145 ( 
.A(n_1004),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1004),
.B(n_780),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_988),
.Y(n_1147)
);

AND2x6_ASAP7_75t_L g1148 ( 
.A(n_977),
.B(n_678),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1081),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1082),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1086),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_950),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1100),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1087),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_973),
.B(n_515),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_917),
.B(n_620),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_959),
.B(n_963),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1088),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1094),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1102),
.B(n_485),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_919),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1115),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1110),
.B(n_486),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1004),
.B(n_596),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1069),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1097),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1115),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_969),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_979),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_927),
.B(n_597),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_917),
.B(n_621),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1042),
.B(n_541),
.Y(n_1172)
);

OR2x6_ASAP7_75t_L g1173 ( 
.A(n_1020),
.B(n_628),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_956),
.B(n_718),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_950),
.B(n_488),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1099),
.Y(n_1176)
);

INVx5_ASAP7_75t_L g1177 ( 
.A(n_919),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_981),
.B(n_718),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_927),
.B(n_781),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_941),
.A2(n_642),
.B1(n_646),
.B2(n_633),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_970),
.Y(n_1181)
);

OA22x2_ASAP7_75t_L g1182 ( 
.A1(n_918),
.A2(n_654),
.B1(n_667),
.B2(n_650),
.Y(n_1182)
);

AND2x6_ASAP7_75t_L g1183 ( 
.A(n_1003),
.B(n_678),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1058),
.A2(n_741),
.B1(n_754),
.B2(n_736),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1105),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_979),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_970),
.B(n_490),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1106),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_962),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_917),
.B(n_1085),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1085),
.B(n_672),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_941),
.A2(n_685),
.B1(n_691),
.B2(n_675),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_958),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_971),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_962),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1084),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1085),
.B(n_517),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_962),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_971),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_929),
.B(n_636),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_941),
.B(n_699),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_954),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_958),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_954),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_960),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_999),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1011),
.Y(n_1207)
);

AND2x2_ASAP7_75t_SL g1208 ( 
.A(n_1058),
.B(n_501),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_937),
.B(n_641),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1114),
.Y(n_1210)
);

BUFx4f_ASAP7_75t_L g1211 ( 
.A(n_1014),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_931),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_937),
.B(n_663),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_931),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_947),
.B(n_1003),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1116),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_944),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_921),
.B(n_668),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1079),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1079),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_934),
.A2(n_782),
.B1(n_778),
.B2(n_500),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_936),
.Y(n_1222)
);

INVx6_ASAP7_75t_L g1223 ( 
.A(n_999),
.Y(n_1223)
);

AND2x6_ASAP7_75t_L g1224 ( 
.A(n_931),
.B(n_670),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1083),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1083),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1111),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1111),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1072),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1072),
.Y(n_1230)
);

AND2x6_ASAP7_75t_L g1231 ( 
.A(n_1009),
.B(n_695),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_936),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_1034),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_942),
.A2(n_711),
.B1(n_715),
.B2(n_702),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_999),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_980),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1069),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_951),
.B(n_743),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_928),
.B(n_494),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_980),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_995),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_995),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_995),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1096),
.B(n_522),
.Y(n_1244)
);

CKINVDCx8_ASAP7_75t_R g1245 ( 
.A(n_1040),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_936),
.Y(n_1246)
);

NOR2x1p5_ASAP7_75t_L g1247 ( 
.A(n_998),
.B(n_525),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_961),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_921),
.B(n_706),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_942),
.A2(n_724),
.B1(n_725),
.B2(n_716),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1101),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_936),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1011),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_947),
.B(n_732),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1107),
.B(n_531),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1069),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_967),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_998),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_971),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_989),
.B(n_532),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_947),
.B(n_708),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1008),
.B(n_735),
.Y(n_1262)
);

AND2x6_ASAP7_75t_L g1263 ( 
.A(n_935),
.B(n_723),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_942),
.B(n_727),
.Y(n_1264)
);

OR2x6_ASAP7_75t_L g1265 ( 
.A(n_1020),
.B(n_745),
.Y(n_1265)
);

INVx8_ASAP7_75t_L g1266 ( 
.A(n_1020),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1108),
.B(n_547),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_975),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1047),
.B(n_613),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_925),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_968),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_978),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_925),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_982),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_984),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_932),
.B(n_737),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_985),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_968),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_943),
.B(n_739),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_930),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_996),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_992),
.B(n_550),
.Y(n_1282)
);

BUFx4f_ASAP7_75t_L g1283 ( 
.A(n_1014),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_939),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_919),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1104),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_920),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_932),
.B(n_751),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1006),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_939),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_945),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_966),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_945),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_972),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_972),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_974),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_974),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_976),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_SL g1299 ( 
.A(n_1000),
.B(n_477),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_983),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_964),
.Y(n_1301)
);

AND3x2_ASAP7_75t_L g1302 ( 
.A(n_1054),
.B(n_744),
.C(n_741),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_983),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1044),
.B(n_552),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_946),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_987),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1022),
.B(n_747),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_987),
.Y(n_1308)
);

NOR3xp33_ASAP7_75t_L g1309 ( 
.A(n_1051),
.B(n_677),
.C(n_639),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1063),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_990),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_943),
.B(n_756),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_990),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_993),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_943),
.Y(n_1315)
);

BUFx8_ASAP7_75t_SL g1316 ( 
.A(n_1055),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_993),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_922),
.B(n_560),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_933),
.B(n_483),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1001),
.Y(n_1320)
);

AND2x6_ASAP7_75t_L g1321 ( 
.A(n_1018),
.B(n_560),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1001),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1002),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1006),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1002),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_938),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_940),
.Y(n_1327)
);

INVx4_ASAP7_75t_SL g1328 ( 
.A(n_1006),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1006),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1022),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_948),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_997),
.B(n_507),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1058),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1050),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_949),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_919),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_952),
.Y(n_1337)
);

INVx5_ASAP7_75t_L g1338 ( 
.A(n_926),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_953),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_997),
.B(n_484),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1043),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1043),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1019),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_922),
.B(n_560),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1044),
.B(n_555),
.Y(n_1345)
);

BUFx4f_ASAP7_75t_L g1346 ( 
.A(n_1019),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1019),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1031),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1013),
.B(n_573),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1031),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1023),
.B(n_750),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_923),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1064),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1013),
.B(n_611),
.Y(n_1354)
);

CKINVDCx8_ASAP7_75t_R g1355 ( 
.A(n_1049),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1113),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1071),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1071),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_957),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1044),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1023),
.B(n_753),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1017),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1027),
.B(n_664),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1278),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1190),
.B(n_1025),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1190),
.B(n_1025),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1196),
.B(n_1027),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1196),
.B(n_1028),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1141),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1297),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1168),
.B(n_1029),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1152),
.B(n_1017),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1121),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1181),
.A2(n_994),
.B1(n_1028),
.B2(n_1030),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1236),
.Y(n_1375)
);

OAI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1180),
.A2(n_957),
.B1(n_1032),
.B2(n_1030),
.C(n_1016),
.Y(n_1376)
);

OAI221xp5_ASAP7_75t_L g1377 ( 
.A1(n_1180),
.A2(n_1032),
.B1(n_1024),
.B2(n_1026),
.C(n_1021),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1184),
.A2(n_1055),
.B1(n_1057),
.B2(n_1054),
.Y(n_1378)
);

OAI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1192),
.A2(n_1035),
.B1(n_1036),
.B2(n_1033),
.C(n_1015),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1157),
.Y(n_1380)
);

AO22x2_ASAP7_75t_L g1381 ( 
.A1(n_1184),
.A2(n_1055),
.B1(n_1060),
.B2(n_1057),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1181),
.Y(n_1382)
);

NOR2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1165),
.B(n_1017),
.Y(n_1383)
);

AND2x2_ASAP7_75t_SL g1384 ( 
.A(n_1194),
.B(n_1049),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1136),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1292),
.B(n_994),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1157),
.Y(n_1387)
);

OAI221xp5_ASAP7_75t_L g1388 ( 
.A1(n_1192),
.A2(n_1012),
.B1(n_1062),
.B2(n_1065),
.C(n_1060),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1120),
.Y(n_1389)
);

AO22x2_ASAP7_75t_L g1390 ( 
.A1(n_1343),
.A2(n_1065),
.B1(n_1062),
.B2(n_1038),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1130),
.Y(n_1391)
);

OAI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1360),
.A2(n_1012),
.B1(n_1037),
.B2(n_1041),
.C(n_1039),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1132),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1133),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1153),
.Y(n_1395)
);

AO22x2_ASAP7_75t_L g1396 ( 
.A1(n_1341),
.A2(n_1045),
.B1(n_1048),
.B2(n_1046),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1126),
.B(n_1053),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1175),
.B(n_1187),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1215),
.A2(n_1053),
.B1(n_1059),
.B2(n_1010),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1138),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1149),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1122),
.B(n_1059),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1236),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1360),
.A2(n_1144),
.B1(n_1309),
.B2(n_1251),
.C(n_1128),
.Y(n_1404)
);

AO22x2_ASAP7_75t_L g1405 ( 
.A1(n_1342),
.A2(n_1056),
.B1(n_1061),
.B2(n_1052),
.Y(n_1405)
);

OR2x6_ASAP7_75t_SL g1406 ( 
.A(n_1237),
.B(n_1066),
.Y(n_1406)
);

AO22x2_ASAP7_75t_L g1407 ( 
.A1(n_1307),
.A2(n_1147),
.B1(n_1309),
.B2(n_1347),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1215),
.A2(n_1059),
.B1(n_561),
.B2(n_564),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_SL g1409 ( 
.A(n_1199),
.B(n_744),
.Y(n_1409)
);

OR2x2_ASAP7_75t_SL g1410 ( 
.A(n_1143),
.B(n_1067),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1256),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1248),
.B(n_1068),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1150),
.Y(n_1413)
);

AO22x2_ASAP7_75t_L g1414 ( 
.A1(n_1307),
.A2(n_1347),
.B1(n_1253),
.B2(n_1070),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1151),
.Y(n_1415)
);

INVx8_ASAP7_75t_L g1416 ( 
.A(n_1266),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1154),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_SL g1418 ( 
.A(n_1193),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1203),
.B(n_690),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1158),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1310),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1362),
.B(n_761),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1128),
.B(n_558),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1159),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1239),
.A2(n_567),
.B1(n_580),
.B2(n_566),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1166),
.Y(n_1426)
);

OAI221xp5_ASAP7_75t_L g1427 ( 
.A1(n_1135),
.A2(n_755),
.B1(n_693),
.B2(n_598),
.C(n_610),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1135),
.B(n_587),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1176),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1185),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1143),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1188),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1244),
.A2(n_1255),
.B1(n_1353),
.B2(n_1260),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1280),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1243),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1155),
.B(n_606),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1217),
.A2(n_616),
.B1(n_617),
.B2(n_612),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1155),
.B(n_624),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1210),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1333),
.A2(n_779),
.B1(n_786),
.B2(n_754),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1243),
.Y(n_1441)
);

NAND2x1p5_ASAP7_75t_L g1442 ( 
.A(n_1259),
.B(n_762),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1216),
.Y(n_1443)
);

NAND2x1p5_ASAP7_75t_L g1444 ( 
.A(n_1348),
.B(n_773),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1124),
.Y(n_1445)
);

AO22x2_ASAP7_75t_L g1446 ( 
.A1(n_1273),
.A2(n_779),
.B1(n_786),
.B2(n_784),
.Y(n_1446)
);

NAND2x1p5_ASAP7_75t_L g1447 ( 
.A(n_1350),
.B(n_777),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1124),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1326),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_L g1450 ( 
.A(n_1258),
.B(n_9),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1119),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1327),
.Y(n_1452)
);

NAND2x1p5_ASAP7_75t_L g1453 ( 
.A(n_1247),
.B(n_501),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1156),
.B(n_501),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1160),
.B(n_1163),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1335),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1337),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1339),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1221),
.A2(n_626),
.B1(n_637),
.B2(n_635),
.C(n_630),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1268),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1272),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1304),
.B(n_652),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1274),
.Y(n_1463)
);

AO22x2_ASAP7_75t_L g1464 ( 
.A1(n_1273),
.A2(n_740),
.B1(n_748),
.B2(n_681),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1275),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1277),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1267),
.A2(n_657),
.B1(n_671),
.B2(n_655),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1156),
.B(n_600),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1316),
.Y(n_1469)
);

AO22x2_ASAP7_75t_L g1470 ( 
.A1(n_1330),
.A2(n_776),
.B1(n_11),
.B2(n_9),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1281),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1282),
.A2(n_684),
.B1(n_686),
.B2(n_673),
.Y(n_1472)
);

AO22x2_ASAP7_75t_L g1473 ( 
.A1(n_1118),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1197),
.B(n_688),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1359),
.A2(n_698),
.B1(n_700),
.B2(n_697),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_1119),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1331),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1331),
.Y(n_1478)
);

AO22x2_ASAP7_75t_L g1479 ( 
.A1(n_1140),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1345),
.B(n_701),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1119),
.Y(n_1481)
);

AO22x2_ASAP7_75t_L g1482 ( 
.A1(n_1302),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1171),
.Y(n_1483)
);

AO22x2_ASAP7_75t_L g1484 ( 
.A1(n_1302),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1191),
.B(n_600),
.Y(n_1485)
);

AO22x2_ASAP7_75t_L g1486 ( 
.A1(n_1129),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1261),
.A2(n_728),
.B1(n_746),
.B2(n_717),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1298),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1303),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1306),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1191),
.B(n_600),
.Y(n_1491)
);

CKINVDCx16_ASAP7_75t_R g1492 ( 
.A(n_1299),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1173),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1240),
.Y(n_1494)
);

AO22x2_ASAP7_75t_L g1495 ( 
.A1(n_1129),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1265),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1299),
.B(n_493),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1241),
.Y(n_1498)
);

AO22x2_ASAP7_75t_L g1499 ( 
.A1(n_1129),
.A2(n_28),
.B1(n_25),
.B2(n_26),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1125),
.B(n_759),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1242),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1284),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1172),
.A2(n_769),
.B1(n_774),
.B2(n_770),
.C(n_764),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1284),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1290),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1254),
.B(n_666),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1266),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1351),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1261),
.A2(n_775),
.B1(n_1076),
.B2(n_1073),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_SL g1510 ( 
.A(n_1245),
.B(n_498),
.C(n_496),
.Y(n_1510)
);

AO22x2_ASAP7_75t_L g1511 ( 
.A1(n_1254),
.A2(n_29),
.B1(n_25),
.B2(n_28),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1238),
.B(n_1076),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1131),
.A2(n_1091),
.B1(n_1092),
.B2(n_1089),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1351),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1208),
.A2(n_1089),
.B1(n_1092),
.B2(n_1091),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1290),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1361),
.Y(n_1517)
);

AO22x2_ASAP7_75t_L g1518 ( 
.A1(n_1279),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_SL g1519 ( 
.A(n_1355),
.B(n_520),
.C(n_502),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1291),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1361),
.B(n_1201),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1211),
.A2(n_1093),
.B1(n_1098),
.B2(n_1095),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1308),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1313),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1269),
.B(n_1112),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_SL g1526 ( 
.A(n_1334),
.B(n_1301),
.C(n_1286),
.Y(n_1526)
);

NOR2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1316),
.B(n_523),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1315),
.Y(n_1528)
);

AO22x2_ASAP7_75t_L g1529 ( 
.A1(n_1279),
.A2(n_37),
.B1(n_33),
.B2(n_35),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1314),
.Y(n_1530)
);

INVx2_ASAP7_75t_SL g1531 ( 
.A(n_1266),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1201),
.B(n_38),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1291),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1224),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1317),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1322),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1263),
.B(n_530),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1325),
.Y(n_1538)
);

AO22x2_ASAP7_75t_L g1539 ( 
.A1(n_1312),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1229),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1230),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1212),
.Y(n_1542)
);

AO22x2_ASAP7_75t_L g1543 ( 
.A1(n_1312),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1293),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1289),
.B(n_785),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1293),
.Y(n_1546)
);

AO22x2_ASAP7_75t_L g1547 ( 
.A1(n_1145),
.A2(n_1264),
.B1(n_1283),
.B2(n_1211),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1263),
.B(n_542),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1352),
.Y(n_1549)
);

AO22x2_ASAP7_75t_L g1550 ( 
.A1(n_1145),
.A2(n_46),
.B1(n_42),
.B2(n_45),
.Y(n_1550)
);

BUFx8_ASAP7_75t_L g1551 ( 
.A(n_1117),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1182),
.A2(n_1174),
.B1(n_1276),
.B2(n_1288),
.C(n_1134),
.Y(n_1552)
);

AO22x2_ASAP7_75t_L g1553 ( 
.A1(n_1145),
.A2(n_46),
.B1(n_42),
.B2(n_45),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1263),
.B(n_1276),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1357),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1263),
.B(n_546),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1289),
.B(n_785),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1270),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1182),
.A2(n_785),
.B1(n_562),
.B2(n_563),
.C(n_557),
.Y(n_1559)
);

OAI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1174),
.A2(n_575),
.B1(n_578),
.B2(n_576),
.C(n_556),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1358),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1233),
.B(n_581),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1305),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1134),
.A2(n_585),
.B1(n_605),
.B2(n_599),
.C(n_595),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1283),
.B(n_615),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1212),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1214),
.Y(n_1567)
);

AO22x2_ASAP7_75t_L g1568 ( 
.A1(n_1264),
.A2(n_1346),
.B1(n_1328),
.B2(n_1329),
.Y(n_1568)
);

AO22x2_ASAP7_75t_L g1569 ( 
.A1(n_1346),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1324),
.B(n_1103),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1214),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1219),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1220),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1225),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1226),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1227),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1270),
.B(n_618),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1228),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1305),
.Y(n_1579)
);

AO22x2_ASAP7_75t_L g1580 ( 
.A1(n_1328),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1580)
);

AO22x2_ASAP7_75t_L g1581 ( 
.A1(n_1328),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1257),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1262),
.B(n_52),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1148),
.B(n_1231),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1271),
.Y(n_1585)
);

AND2x6_ASAP7_75t_L g1586 ( 
.A(n_1137),
.B(n_560),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1294),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1295),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1296),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1300),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1311),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1320),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1148),
.B(n_629),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1323),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1324),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1262),
.B(n_53),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1319),
.Y(n_1597)
);

AO22x2_ASAP7_75t_L g1598 ( 
.A1(n_1329),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1170),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1363),
.A2(n_648),
.B1(n_653),
.B2(n_645),
.C(n_634),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1224),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1207),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1183),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1137),
.Y(n_1604)
);

AO22x2_ASAP7_75t_L g1605 ( 
.A1(n_1301),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1492),
.B(n_1162),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1395),
.B(n_1162),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1398),
.B(n_1382),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1380),
.B(n_1387),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1385),
.B(n_1167),
.Y(n_1610)
);

NAND2xp33_ASAP7_75t_SL g1611 ( 
.A(n_1534),
.B(n_1315),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1534),
.B(n_1315),
.Y(n_1612)
);

AND3x1_ASAP7_75t_L g1613 ( 
.A(n_1409),
.B(n_1399),
.C(n_1433),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_SL g1614 ( 
.A(n_1601),
.B(n_1287),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1372),
.B(n_1319),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1373),
.B(n_1189),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1451),
.B(n_1189),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1445),
.B(n_1234),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1448),
.B(n_1234),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1525),
.B(n_1363),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1442),
.B(n_1250),
.Y(n_1621)
);

NAND2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1528),
.B(n_1287),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1597),
.B(n_1231),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1521),
.B(n_1349),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1493),
.B(n_1250),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1521),
.B(n_1231),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1496),
.B(n_1161),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1476),
.B(n_1177),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1481),
.B(n_1444),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1528),
.B(n_1287),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1455),
.B(n_1389),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1447),
.B(n_1507),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1397),
.B(n_1177),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1397),
.B(n_1177),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1371),
.B(n_1177),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1419),
.B(n_1285),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1391),
.B(n_1195),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1421),
.B(n_1285),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1384),
.B(n_1285),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1416),
.B(n_1285),
.Y(n_1640)
);

NAND2xp33_ASAP7_75t_SL g1641 ( 
.A(n_1596),
.B(n_1340),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1393),
.B(n_1231),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1416),
.B(n_1338),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1551),
.B(n_1338),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1551),
.B(n_1531),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1394),
.B(n_1400),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1402),
.B(n_1349),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1367),
.B(n_1354),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1368),
.B(n_1354),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1374),
.B(n_1178),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1401),
.B(n_1332),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1596),
.B(n_1178),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1413),
.B(n_1332),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1386),
.B(n_1340),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1440),
.B(n_1412),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1554),
.B(n_1123),
.Y(n_1656)
);

NAND2xp33_ASAP7_75t_SL g1657 ( 
.A(n_1418),
.B(n_1123),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1562),
.B(n_1169),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1472),
.B(n_1169),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1415),
.B(n_1417),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1420),
.B(n_1224),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1437),
.B(n_1169),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1528),
.B(n_1146),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1424),
.B(n_1224),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1475),
.B(n_1186),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1426),
.B(n_1429),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1602),
.B(n_1164),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1593),
.B(n_1206),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1584),
.B(n_1164),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1430),
.B(n_1198),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_SL g1671 ( 
.A(n_1603),
.B(n_1206),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1509),
.B(n_1425),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1487),
.B(n_1537),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1548),
.B(n_658),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1556),
.B(n_665),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1485),
.B(n_669),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1491),
.B(n_1369),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1408),
.B(n_676),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1506),
.B(n_694),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1432),
.B(n_1183),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1462),
.B(n_705),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1480),
.B(n_707),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1532),
.B(n_1170),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1364),
.B(n_709),
.Y(n_1684)
);

NAND2xp33_ASAP7_75t_SL g1685 ( 
.A(n_1370),
.B(n_1179),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_SL g1686 ( 
.A(n_1370),
.B(n_1179),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1375),
.B(n_710),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1403),
.B(n_712),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1435),
.B(n_713),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1441),
.B(n_722),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1500),
.B(n_726),
.Y(n_1691)
);

NAND2xp33_ASAP7_75t_SL g1692 ( 
.A(n_1488),
.B(n_1200),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1365),
.B(n_729),
.Y(n_1693)
);

NAND2xp33_ASAP7_75t_SL g1694 ( 
.A(n_1488),
.B(n_1489),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1365),
.B(n_752),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1366),
.B(n_758),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_SL g1697 ( 
.A(n_1489),
.B(n_1200),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1366),
.B(n_763),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1422),
.B(n_766),
.Y(n_1699)
);

NAND2xp33_ASAP7_75t_SL g1700 ( 
.A(n_1490),
.B(n_1209),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1422),
.B(n_767),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1450),
.B(n_772),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1512),
.B(n_1549),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1439),
.B(n_1209),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1549),
.B(n_1356),
.Y(n_1705)
);

NAND2xp33_ASAP7_75t_SL g1706 ( 
.A(n_1490),
.B(n_1213),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1443),
.B(n_1213),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1555),
.B(n_1561),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1446),
.B(n_1218),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1449),
.B(n_1218),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1452),
.B(n_1249),
.Y(n_1711)
);

NAND2xp33_ASAP7_75t_SL g1712 ( 
.A(n_1515),
.B(n_1249),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1474),
.B(n_1483),
.Y(n_1713)
);

AND2x2_ASAP7_75t_SL g1714 ( 
.A(n_1547),
.B(n_583),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1456),
.B(n_1202),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1467),
.B(n_1235),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1457),
.B(n_1204),
.Y(n_1717)
);

NAND2xp33_ASAP7_75t_R g1718 ( 
.A(n_1411),
.B(n_1235),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_SL g1719 ( 
.A(n_1522),
.B(n_1205),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1458),
.B(n_1127),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1423),
.B(n_1428),
.Y(n_1721)
);

NAND2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1477),
.B(n_1139),
.Y(n_1722)
);

NAND2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1478),
.B(n_1142),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1436),
.B(n_1438),
.Y(n_1724)
);

AND3x1_ASAP7_75t_L g1725 ( 
.A(n_1431),
.B(n_59),
.C(n_60),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1460),
.B(n_1223),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1446),
.B(n_59),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_SL g1728 ( 
.A(n_1523),
.B(n_1222),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1434),
.B(n_1109),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1454),
.B(n_1468),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1524),
.B(n_1232),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1461),
.B(n_1463),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_SL g1733 ( 
.A(n_1530),
.B(n_1246),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1392),
.B(n_1223),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1465),
.B(n_1252),
.Y(n_1735)
);

NAND2xp33_ASAP7_75t_SL g1736 ( 
.A(n_1535),
.B(n_1318),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1508),
.B(n_1514),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1536),
.B(n_1318),
.Y(n_1738)
);

NAND2xp33_ASAP7_75t_SL g1739 ( 
.A(n_1538),
.B(n_1344),
.Y(n_1739)
);

AND3x1_ASAP7_75t_L g1740 ( 
.A(n_1583),
.B(n_62),
.C(n_63),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1517),
.B(n_1582),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1466),
.B(n_1223),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1471),
.B(n_1321),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_SL g1744 ( 
.A(n_1418),
.B(n_583),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_SL g1745 ( 
.A(n_1527),
.B(n_604),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1577),
.B(n_1497),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1453),
.B(n_760),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1410),
.B(n_62),
.Y(n_1748)
);

AND2x2_ASAP7_75t_SL g1749 ( 
.A(n_1547),
.B(n_63),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_SL g1750 ( 
.A(n_1383),
.B(n_64),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1552),
.B(n_1336),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1585),
.B(n_1336),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1587),
.B(n_65),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_SL g1754 ( 
.A(n_1558),
.B(n_65),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1588),
.B(n_66),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1572),
.B(n_67),
.Y(n_1756)
);

NAND2xp33_ASAP7_75t_SL g1757 ( 
.A(n_1595),
.B(n_68),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1589),
.B(n_68),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1590),
.B(n_69),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1469),
.B(n_69),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1591),
.B(n_70),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1592),
.B(n_70),
.Y(n_1762)
);

NAND2xp33_ASAP7_75t_SL g1763 ( 
.A(n_1594),
.B(n_71),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1513),
.B(n_71),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1545),
.B(n_72),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1557),
.B(n_72),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1501),
.B(n_74),
.Y(n_1767)
);

NAND2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1604),
.B(n_75),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1604),
.B(n_78),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1502),
.B(n_81),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1504),
.B(n_82),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1505),
.B(n_83),
.Y(n_1772)
);

NAND2xp33_ASAP7_75t_SL g1773 ( 
.A(n_1516),
.B(n_85),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1520),
.B(n_85),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1533),
.B(n_86),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1544),
.B(n_86),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1546),
.B(n_88),
.Y(n_1777)
);

NAND2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1563),
.B(n_88),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1579),
.B(n_89),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1599),
.B(n_89),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1573),
.B(n_91),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1494),
.B(n_91),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1498),
.B(n_92),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1570),
.B(n_93),
.Y(n_1784)
);

NAND2xp33_ASAP7_75t_SL g1785 ( 
.A(n_1542),
.B(n_1566),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1574),
.B(n_93),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1575),
.B(n_95),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1576),
.B(n_96),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1578),
.B(n_96),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1567),
.B(n_97),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1378),
.B(n_98),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1378),
.B(n_99),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1571),
.B(n_99),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_SL g1794 ( 
.A(n_1565),
.B(n_101),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1404),
.B(n_101),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1407),
.B(n_102),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1540),
.B(n_1541),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1510),
.B(n_1519),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1407),
.B(n_104),
.Y(n_1799)
);

NAND2xp33_ASAP7_75t_SL g1800 ( 
.A(n_1568),
.B(n_105),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1379),
.B(n_106),
.Y(n_1801)
);

NAND2xp33_ASAP7_75t_SL g1802 ( 
.A(n_1568),
.B(n_106),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1406),
.B(n_107),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1414),
.B(n_108),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1396),
.B(n_108),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1381),
.B(n_109),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1381),
.B(n_109),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1464),
.B(n_110),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1427),
.B(n_111),
.Y(n_1809)
);

NAND2xp33_ASAP7_75t_SL g1810 ( 
.A(n_1486),
.B(n_111),
.Y(n_1810)
);

NAND2xp33_ASAP7_75t_SL g1811 ( 
.A(n_1486),
.B(n_112),
.Y(n_1811)
);

NAND2xp33_ASAP7_75t_SL g1812 ( 
.A(n_1495),
.B(n_113),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1511),
.B(n_114),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1376),
.B(n_115),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1388),
.B(n_115),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1377),
.B(n_116),
.Y(n_1816)
);

AND2x2_ASAP7_75t_SL g1817 ( 
.A(n_1470),
.B(n_116),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1503),
.B(n_121),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1390),
.B(n_121),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1390),
.B(n_122),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1586),
.B(n_1396),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1586),
.B(n_1405),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1586),
.B(n_122),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1586),
.B(n_124),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1405),
.B(n_124),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1470),
.B(n_125),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1600),
.B(n_126),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1459),
.B(n_1564),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1560),
.B(n_128),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1495),
.B(n_128),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1499),
.B(n_129),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1559),
.B(n_129),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1473),
.B(n_130),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1499),
.B(n_130),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1473),
.B(n_131),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1479),
.B(n_131),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1479),
.B(n_132),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1550),
.B(n_133),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1511),
.B(n_135),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1518),
.B(n_136),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1605),
.B(n_137),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1550),
.B(n_138),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1553),
.B(n_138),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1553),
.B(n_140),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1518),
.B(n_140),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1529),
.B(n_141),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1529),
.B(n_141),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1539),
.B(n_142),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1539),
.B(n_143),
.Y(n_1849)
);

NAND2xp33_ASAP7_75t_SL g1850 ( 
.A(n_1580),
.B(n_1581),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1543),
.B(n_144),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1543),
.B(n_145),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1526),
.B(n_146),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_SL g1854 ( 
.A(n_1580),
.B(n_147),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1581),
.B(n_147),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1482),
.B(n_148),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1598),
.B(n_148),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1598),
.B(n_150),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1569),
.B(n_150),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1569),
.B(n_151),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1605),
.B(n_152),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1482),
.B(n_152),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1484),
.B(n_153),
.Y(n_1863)
);

NAND2xp33_ASAP7_75t_SL g1864 ( 
.A(n_1484),
.B(n_153),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1609),
.B(n_1647),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1715),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1620),
.A2(n_155),
.B(n_156),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1637),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1719),
.A2(n_292),
.B(n_288),
.Y(n_1869)
);

OAI22x1_ASAP7_75t_L g1870 ( 
.A1(n_1859),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1608),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1655),
.B(n_157),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1714),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1714),
.Y(n_1874)
);

OA21x2_ASAP7_75t_L g1875 ( 
.A1(n_1806),
.A2(n_298),
.B(n_293),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1613),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1641),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1756),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1631),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1629),
.B(n_165),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1618),
.A2(n_165),
.B(n_166),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1624),
.B(n_167),
.Y(n_1882)
);

OR2x6_ASAP7_75t_L g1883 ( 
.A(n_1859),
.B(n_168),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1756),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1619),
.A2(n_171),
.B(n_172),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1694),
.A2(n_306),
.B(n_304),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1801),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1694),
.A2(n_310),
.B(n_307),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1718),
.Y(n_1889)
);

O2A1O1Ixp5_ASAP7_75t_L g1890 ( 
.A1(n_1665),
.A2(n_313),
.B(n_315),
.C(n_312),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1859),
.A2(n_177),
.B1(n_173),
.B2(n_176),
.Y(n_1891)
);

OAI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1651),
.A2(n_176),
.B(n_177),
.Y(n_1892)
);

NOR2xp67_ASAP7_75t_L g1893 ( 
.A(n_1748),
.B(n_178),
.Y(n_1893)
);

OAI21x1_ASAP7_75t_L g1894 ( 
.A1(n_1705),
.A2(n_323),
.B(n_317),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1653),
.B(n_178),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1841),
.A2(n_180),
.B(n_181),
.Y(n_1896)
);

AO31x2_ASAP7_75t_L g1897 ( 
.A1(n_1796),
.A2(n_180),
.A3(n_182),
.B(n_185),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1672),
.A2(n_182),
.B(n_187),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1646),
.B(n_187),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1828),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1721),
.A2(n_326),
.B(n_324),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1756),
.Y(n_1902)
);

AO21x2_ASAP7_75t_L g1903 ( 
.A1(n_1807),
.A2(n_333),
.B(n_331),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1660),
.B(n_189),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1850),
.Y(n_1905)
);

AO31x2_ASAP7_75t_L g1906 ( 
.A1(n_1805),
.A2(n_190),
.A3(n_191),
.B(n_192),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1644),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1717),
.Y(n_1908)
);

CKINVDCx14_ASAP7_75t_R g1909 ( 
.A(n_1745),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1749),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1781),
.Y(n_1911)
);

INVxp67_ASAP7_75t_SL g1912 ( 
.A(n_1781),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1666),
.Y(n_1913)
);

AO22x2_ASAP7_75t_L g1914 ( 
.A1(n_1826),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1645),
.B(n_193),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1732),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_SL g1917 ( 
.A1(n_1840),
.A2(n_194),
.B(n_195),
.Y(n_1917)
);

INVx2_ASAP7_75t_SL g1918 ( 
.A(n_1632),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1813),
.B(n_196),
.Y(n_1919)
);

OR2x6_ASAP7_75t_L g1920 ( 
.A(n_1781),
.B(n_197),
.Y(n_1920)
);

AOI21x1_ASAP7_75t_SL g1921 ( 
.A1(n_1795),
.A2(n_197),
.B(n_198),
.Y(n_1921)
);

OAI21x1_ASAP7_75t_L g1922 ( 
.A1(n_1668),
.A2(n_348),
.B(n_345),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1749),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1709),
.B(n_200),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1637),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1652),
.B(n_1724),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1637),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1615),
.B(n_200),
.Y(n_1928)
);

INVx1_ASAP7_75t_SL g1929 ( 
.A(n_1636),
.Y(n_1929)
);

AO31x2_ASAP7_75t_L g1930 ( 
.A1(n_1751),
.A2(n_201),
.A3(n_202),
.B(n_203),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1648),
.A2(n_203),
.B(n_204),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1649),
.A2(n_1815),
.B(n_1816),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1711),
.B(n_204),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1711),
.B(n_1621),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1727),
.B(n_205),
.Y(n_1935)
);

NAND2x1p5_ASAP7_75t_L g1936 ( 
.A(n_1677),
.B(n_206),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1711),
.B(n_207),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1713),
.B(n_207),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_SL g1939 ( 
.A1(n_1847),
.A2(n_208),
.B(n_209),
.Y(n_1939)
);

AO31x2_ASAP7_75t_L g1940 ( 
.A1(n_1833),
.A2(n_208),
.A3(n_209),
.B(n_210),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1830),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1625),
.B(n_210),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1691),
.B(n_211),
.Y(n_1943)
);

INVx5_ASAP7_75t_L g1944 ( 
.A(n_1791),
.Y(n_1944)
);

INVx3_ASAP7_75t_SL g1945 ( 
.A(n_1817),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1704),
.B(n_211),
.Y(n_1946)
);

O2A1O1Ixp5_ASAP7_75t_L g1947 ( 
.A1(n_1821),
.A2(n_378),
.B(n_463),
.C(n_462),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1822),
.A2(n_369),
.B(n_368),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1850),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1831),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1707),
.B(n_212),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1810),
.A2(n_212),
.B(n_214),
.C(n_215),
.Y(n_1952)
);

INVxp67_ASAP7_75t_SL g1953 ( 
.A(n_1730),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1744),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1720),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1650),
.B(n_216),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_SL g1957 ( 
.A1(n_1839),
.A2(n_216),
.B(n_218),
.Y(n_1957)
);

OA21x2_ASAP7_75t_L g1958 ( 
.A1(n_1799),
.A2(n_384),
.B(n_460),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1818),
.B(n_219),
.Y(n_1959)
);

O2A1O1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1808),
.A2(n_220),
.B(n_221),
.C(n_222),
.Y(n_1960)
);

AOI221x1_ASAP7_75t_L g1961 ( 
.A1(n_1810),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.C(n_227),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1708),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1817),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1814),
.A2(n_228),
.B(n_230),
.Y(n_1964)
);

A2O1A1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1811),
.A2(n_231),
.B(n_232),
.C(n_233),
.Y(n_1965)
);

NAND3xp33_ASAP7_75t_L g1966 ( 
.A(n_1854),
.B(n_233),
.C(n_234),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1654),
.A2(n_235),
.B(n_237),
.Y(n_1967)
);

A2O1A1Ixp33_ASAP7_75t_L g1968 ( 
.A1(n_1811),
.A2(n_237),
.B(n_238),
.C(n_239),
.Y(n_1968)
);

NOR2xp67_ASAP7_75t_L g1969 ( 
.A(n_1803),
.B(n_238),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1710),
.B(n_239),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1812),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1728),
.A2(n_397),
.B(n_453),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1703),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1797),
.B(n_241),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1639),
.Y(n_1975)
);

AO32x2_ASAP7_75t_L g1976 ( 
.A1(n_1812),
.A2(n_242),
.A3(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1734),
.B(n_245),
.Y(n_1977)
);

AND2x6_ASAP7_75t_SL g1978 ( 
.A(n_1856),
.B(n_246),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1670),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1804),
.A2(n_398),
.B(n_447),
.Y(n_1980)
);

OAI21x1_ASAP7_75t_SL g1981 ( 
.A1(n_1623),
.A2(n_247),
.B(n_248),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1678),
.B(n_247),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1670),
.B(n_1809),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1725),
.B(n_248),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1764),
.A2(n_249),
.B(n_251),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1670),
.B(n_249),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1731),
.A2(n_400),
.B(n_446),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1735),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1834),
.Y(n_1989)
);

OAI21x1_ASAP7_75t_SL g1990 ( 
.A1(n_1642),
.A2(n_251),
.B(n_252),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_SL g1991 ( 
.A1(n_1862),
.A2(n_253),
.B(n_254),
.Y(n_1991)
);

AO21x2_ASAP7_75t_L g1992 ( 
.A1(n_1819),
.A2(n_399),
.B(n_439),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1626),
.B(n_253),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1798),
.B(n_254),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1735),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1760),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1737),
.B(n_255),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1827),
.B(n_256),
.Y(n_1998)
);

NAND3xp33_ASAP7_75t_SL g1999 ( 
.A(n_1861),
.B(n_257),
.C(n_260),
.Y(n_1999)
);

INVx2_ASAP7_75t_SL g2000 ( 
.A(n_1640),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1829),
.B(n_260),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1857),
.Y(n_2002)
);

O2A1O1Ixp33_ASAP7_75t_SL g2003 ( 
.A1(n_1838),
.A2(n_379),
.B(n_434),
.C(n_433),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1699),
.B(n_261),
.Y(n_2004)
);

OAI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1858),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1616),
.B(n_262),
.Y(n_2006)
);

AO21x1_ASAP7_75t_L g2007 ( 
.A1(n_1800),
.A2(n_263),
.B(n_264),
.Y(n_2007)
);

AO21x1_ASAP7_75t_L g2008 ( 
.A1(n_1800),
.A2(n_265),
.B(n_266),
.Y(n_2008)
);

NOR4xp25_ASAP7_75t_L g2009 ( 
.A(n_1835),
.B(n_265),
.C(n_266),
.D(n_267),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1643),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1610),
.B(n_267),
.Y(n_2011)
);

NOR2xp67_ASAP7_75t_L g2012 ( 
.A(n_1853),
.B(n_268),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1750),
.Y(n_2013)
);

NOR2xp67_ASAP7_75t_SL g2014 ( 
.A(n_1842),
.B(n_1843),
.Y(n_2014)
);

A2O1A1Ixp33_ASAP7_75t_L g2015 ( 
.A1(n_1864),
.A2(n_1683),
.B(n_1763),
.C(n_1754),
.Y(n_2015)
);

CKINVDCx20_ASAP7_75t_R g2016 ( 
.A(n_1864),
.Y(n_2016)
);

A2O1A1Ixp33_ASAP7_75t_L g2017 ( 
.A1(n_1683),
.A2(n_268),
.B(n_269),
.C(n_270),
.Y(n_2017)
);

AOI21x1_ASAP7_75t_L g2018 ( 
.A1(n_1820),
.A2(n_1846),
.B(n_1845),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1726),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1673),
.A2(n_269),
.B(n_270),
.Y(n_2020)
);

AO31x2_ASAP7_75t_L g2021 ( 
.A1(n_1832),
.A2(n_271),
.A3(n_272),
.B(n_274),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1740),
.B(n_271),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1733),
.A2(n_413),
.B(n_427),
.Y(n_2023)
);

AO31x2_ASAP7_75t_L g2024 ( 
.A1(n_1680),
.A2(n_274),
.A3(n_275),
.B(n_276),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1607),
.B(n_276),
.Y(n_2025)
);

INVx2_ASAP7_75t_SL g2026 ( 
.A(n_1638),
.Y(n_2026)
);

INVxp67_ASAP7_75t_L g2027 ( 
.A(n_1792),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1681),
.B(n_277),
.Y(n_2028)
);

AO21x2_ASAP7_75t_L g2029 ( 
.A1(n_1848),
.A2(n_1851),
.B(n_1849),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1661),
.A2(n_277),
.B(n_279),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1701),
.B(n_279),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1741),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1742),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1860),
.A2(n_280),
.B1(n_371),
.B2(n_372),
.Y(n_2034)
);

INVx5_ASAP7_75t_L g2035 ( 
.A(n_1802),
.Y(n_2035)
);

OAI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1664),
.A2(n_280),
.B(n_374),
.Y(n_2036)
);

OAI21x1_ASAP7_75t_L g2037 ( 
.A1(n_1658),
.A2(n_375),
.B(n_416),
.Y(n_2037)
);

OAI21x1_ASAP7_75t_L g2038 ( 
.A1(n_1743),
.A2(n_417),
.B(n_418),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1633),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1606),
.B(n_421),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1634),
.Y(n_2041)
);

A2O1A1Ixp33_ASAP7_75t_L g2042 ( 
.A1(n_1836),
.A2(n_466),
.B(n_1837),
.C(n_1768),
.Y(n_2042)
);

INVx4_ASAP7_75t_L g2043 ( 
.A(n_1802),
.Y(n_2043)
);

AO32x2_ASAP7_75t_L g2044 ( 
.A1(n_1852),
.A2(n_1855),
.A3(n_1844),
.B1(n_1825),
.B2(n_1863),
.Y(n_2044)
);

AND2x4_ASAP7_75t_L g2045 ( 
.A(n_1676),
.B(n_1679),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_1657),
.Y(n_2046)
);

AO32x2_ASAP7_75t_L g2047 ( 
.A1(n_1757),
.A2(n_1778),
.A3(n_1777),
.B1(n_1776),
.B2(n_1773),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1682),
.B(n_1693),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1695),
.B(n_1696),
.Y(n_2049)
);

NOR2x1_ASAP7_75t_SL g2050 ( 
.A(n_1659),
.B(n_1662),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1698),
.B(n_1628),
.Y(n_2051)
);

AO31x2_ASAP7_75t_L g2052 ( 
.A1(n_1622),
.A2(n_1630),
.A3(n_1712),
.B(n_1667),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1769),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1617),
.B(n_1716),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1794),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1786),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1685),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1685),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1746),
.B(n_1787),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_SL g2060 ( 
.A1(n_1611),
.A2(n_1612),
.B(n_1614),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1879),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1913),
.B(n_1686),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1871),
.B(n_1883),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1883),
.B(n_1788),
.Y(n_2064)
);

INVx1_ASAP7_75t_SL g2065 ( 
.A(n_1902),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_2016),
.A2(n_1706),
.B1(n_1700),
.B2(n_1697),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1912),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1889),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1919),
.B(n_1789),
.Y(n_2069)
);

INVxp67_ASAP7_75t_SL g2070 ( 
.A(n_1873),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1913),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_1920),
.Y(n_2072)
);

INVx1_ASAP7_75t_SL g2073 ( 
.A(n_1920),
.Y(n_2073)
);

NAND3xp33_ASAP7_75t_L g2074 ( 
.A(n_1961),
.B(n_1782),
.C(n_1783),
.Y(n_2074)
);

AOI221x1_ASAP7_75t_L g2075 ( 
.A1(n_1870),
.A2(n_1963),
.B1(n_1914),
.B2(n_1965),
.C(n_1952),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1916),
.Y(n_2076)
);

OA21x2_ASAP7_75t_L g2077 ( 
.A1(n_2057),
.A2(n_1780),
.B(n_1759),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_2060),
.A2(n_1752),
.B(n_1729),
.Y(n_2078)
);

OR2x6_ASAP7_75t_L g2079 ( 
.A(n_1878),
.B(n_1884),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1880),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1865),
.Y(n_2081)
);

NAND3xp33_ASAP7_75t_L g2082 ( 
.A(n_1876),
.B(n_1784),
.C(n_1766),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_1866),
.B(n_1635),
.Y(n_2083)
);

NAND2x1p5_ASAP7_75t_L g2084 ( 
.A(n_1878),
.B(n_1747),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_SL g2085 ( 
.A(n_2043),
.B(n_1611),
.Y(n_2085)
);

BUFx8_ASAP7_75t_L g2086 ( 
.A(n_1915),
.Y(n_2086)
);

INVxp33_ASAP7_75t_L g2087 ( 
.A(n_1915),
.Y(n_2087)
);

NAND2xp33_ASAP7_75t_L g2088 ( 
.A(n_1873),
.B(n_1612),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_2027),
.B(n_1684),
.Y(n_2089)
);

NAND2x1p5_ASAP7_75t_L g2090 ( 
.A(n_1884),
.B(n_1765),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1866),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1940),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1945),
.B(n_1702),
.Y(n_2093)
);

O2A1O1Ixp5_ASAP7_75t_L g2094 ( 
.A1(n_2043),
.A2(n_1614),
.B(n_1669),
.C(n_1663),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1907),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1908),
.B(n_1955),
.Y(n_2096)
);

NAND2x1p5_ASAP7_75t_L g2097 ( 
.A(n_1911),
.B(n_1954),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1935),
.B(n_1790),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1908),
.Y(n_2099)
);

A2O1A1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_2015),
.A2(n_1896),
.B(n_2042),
.C(n_1867),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1955),
.Y(n_2101)
);

OAI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_1887),
.A2(n_1706),
.B1(n_1692),
.B2(n_1762),
.C(n_1761),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1873),
.Y(n_2103)
);

AOI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1893),
.A2(n_1656),
.B1(n_1793),
.B2(n_1755),
.Y(n_2104)
);

OAI21x1_ASAP7_75t_L g2105 ( 
.A1(n_2038),
.A2(n_1767),
.B(n_1753),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1940),
.Y(n_2106)
);

AOI221xp5_ASAP7_75t_L g2107 ( 
.A1(n_1891),
.A2(n_1758),
.B1(n_1770),
.B2(n_1774),
.C(n_1779),
.Y(n_2107)
);

OAI222xp33_ASAP7_75t_L g2108 ( 
.A1(n_2014),
.A2(n_1824),
.B1(n_1823),
.B2(n_1775),
.C1(n_1772),
.C2(n_1771),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2019),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1940),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1906),
.Y(n_2111)
);

AOI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_1910),
.A2(n_1785),
.B1(n_1675),
.B2(n_1674),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1934),
.B(n_1723),
.Y(n_2113)
);

BUFx2_ASAP7_75t_R g2114 ( 
.A(n_1996),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1906),
.Y(n_2115)
);

OAI21x1_ASAP7_75t_L g2116 ( 
.A1(n_1922),
.A2(n_1627),
.B(n_1671),
.Y(n_2116)
);

AO31x2_ASAP7_75t_L g2117 ( 
.A1(n_2058),
.A2(n_1663),
.A3(n_1723),
.B(n_1722),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1984),
.B(n_1690),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1973),
.B(n_1736),
.Y(n_2119)
);

OAI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1932),
.A2(n_1736),
.B(n_1738),
.Y(n_2120)
);

NAND2x1_ASAP7_75t_L g2121 ( 
.A(n_1911),
.B(n_1738),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_1910),
.A2(n_1739),
.B1(n_1688),
.B2(n_1689),
.Y(n_2122)
);

BUFx3_ASAP7_75t_L g2123 ( 
.A(n_1907),
.Y(n_2123)
);

NAND2x1p5_ASAP7_75t_L g2124 ( 
.A(n_1874),
.B(n_1687),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1868),
.Y(n_2125)
);

INVx6_ASAP7_75t_L g2126 ( 
.A(n_1907),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1914),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_SL g2128 ( 
.A1(n_2007),
.A2(n_1739),
.B(n_2008),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_SL g2129 ( 
.A1(n_1957),
.A2(n_1991),
.B(n_1939),
.Y(n_2129)
);

NOR2xp67_ASAP7_75t_L g2130 ( 
.A(n_2035),
.B(n_2013),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_1882),
.B(n_2004),
.Y(n_2131)
);

NAND2x1p5_ASAP7_75t_L g2132 ( 
.A(n_1874),
.B(n_2035),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_1874),
.Y(n_2133)
);

OAI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_1964),
.A2(n_1898),
.B(n_1942),
.Y(n_2134)
);

INVx8_ASAP7_75t_L g2135 ( 
.A(n_2006),
.Y(n_2135)
);

OAI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1881),
.A2(n_1885),
.B(n_1956),
.Y(n_2136)
);

BUFx12f_ASAP7_75t_L g2137 ( 
.A(n_1978),
.Y(n_2137)
);

NAND2x1p5_ASAP7_75t_L g2138 ( 
.A(n_2035),
.B(n_2046),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1925),
.Y(n_2139)
);

OAI21x1_ASAP7_75t_L g2140 ( 
.A1(n_1894),
.A2(n_1921),
.B(n_2037),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_1918),
.Y(n_2141)
);

AOI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_1910),
.A2(n_1923),
.B1(n_2002),
.B2(n_1989),
.Y(n_2142)
);

BUFx8_ASAP7_75t_L g2143 ( 
.A(n_1976),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_1905),
.A2(n_1949),
.B1(n_1909),
.B2(n_1923),
.Y(n_2144)
);

AO21x2_ASAP7_75t_L g2145 ( 
.A1(n_2018),
.A2(n_1917),
.B(n_1981),
.Y(n_2145)
);

O2A1O1Ixp33_ASAP7_75t_SL g2146 ( 
.A1(n_1968),
.A2(n_2017),
.B(n_1892),
.C(n_1966),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_2022),
.Y(n_2147)
);

BUFx2_ASAP7_75t_SL g2148 ( 
.A(n_1969),
.Y(n_2148)
);

CKINVDCx11_ASAP7_75t_R g2149 ( 
.A(n_2045),
.Y(n_2149)
);

AND2x4_ASAP7_75t_L g2150 ( 
.A(n_1927),
.B(n_1979),
.Y(n_2150)
);

INVxp67_ASAP7_75t_L g2151 ( 
.A(n_1938),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_2049),
.B(n_2048),
.Y(n_2152)
);

OA21x2_ASAP7_75t_L g2153 ( 
.A1(n_1869),
.A2(n_1980),
.B(n_2036),
.Y(n_2153)
);

AO21x2_ASAP7_75t_L g2154 ( 
.A1(n_2020),
.A2(n_1990),
.B(n_2050),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_2052),
.Y(n_2155)
);

AOI21xp5_ASAP7_75t_L g2156 ( 
.A1(n_1983),
.A2(n_1972),
.B(n_1987),
.Y(n_2156)
);

OA21x2_ASAP7_75t_L g2157 ( 
.A1(n_1890),
.A2(n_1947),
.B(n_2030),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1995),
.B(n_1962),
.Y(n_2158)
);

AOI21x1_ASAP7_75t_SL g2159 ( 
.A1(n_2040),
.A2(n_1977),
.B(n_1924),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2021),
.Y(n_2160)
);

AO21x2_ASAP7_75t_L g2161 ( 
.A1(n_2029),
.A2(n_1941),
.B(n_1950),
.Y(n_2161)
);

AO32x2_ASAP7_75t_L g2162 ( 
.A1(n_2005),
.A2(n_2034),
.A3(n_2026),
.B1(n_2000),
.B2(n_2010),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2032),
.Y(n_2163)
);

AOI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_1923),
.A2(n_1999),
.B1(n_1944),
.B2(n_2012),
.Y(n_2164)
);

OA21x2_ASAP7_75t_L g2165 ( 
.A1(n_1886),
.A2(n_1888),
.B(n_2023),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_2040),
.Y(n_2166)
);

BUFx2_ASAP7_75t_SL g2167 ( 
.A(n_2006),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1897),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1927),
.Y(n_2169)
);

INVx3_ASAP7_75t_L g2170 ( 
.A(n_1988),
.Y(n_2170)
);

AO21x2_ASAP7_75t_L g2171 ( 
.A1(n_1985),
.A2(n_1967),
.B(n_2054),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2031),
.B(n_1943),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_1979),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1944),
.B(n_1988),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_1975),
.Y(n_2175)
);

INVxp67_ASAP7_75t_SL g2176 ( 
.A(n_1938),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2071),
.B(n_1976),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_2103),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2158),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2127),
.B(n_1897),
.Y(n_2180)
);

INVxp67_ASAP7_75t_R g2181 ( 
.A(n_2063),
.Y(n_2181)
);

BUFx2_ASAP7_75t_L g2182 ( 
.A(n_2070),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2076),
.B(n_1976),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_2072),
.B(n_2045),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2092),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2106),
.Y(n_2186)
);

INVxp67_ASAP7_75t_L g2187 ( 
.A(n_2081),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2176),
.B(n_1944),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2061),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2067),
.B(n_1930),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2091),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2099),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2101),
.Y(n_2193)
);

NAND2x1p5_ASAP7_75t_L g2194 ( 
.A(n_2166),
.B(n_2033),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2067),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2096),
.B(n_1872),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2110),
.Y(n_2197)
);

NAND2x1_ASAP7_75t_L g2198 ( 
.A(n_2166),
.B(n_1948),
.Y(n_2198)
);

INVx4_ASAP7_75t_L g2199 ( 
.A(n_2135),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_2096),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2109),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_2072),
.B(n_1926),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2073),
.B(n_2028),
.Y(n_2203)
);

BUFx2_ASAP7_75t_L g2204 ( 
.A(n_2070),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2080),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_2103),
.Y(n_2206)
);

HB1xp67_ASAP7_75t_L g2207 ( 
.A(n_2175),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2083),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2111),
.B(n_1930),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2163),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2125),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2139),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2062),
.Y(n_2213)
);

AO21x2_ASAP7_75t_L g2214 ( 
.A1(n_2128),
.A2(n_2009),
.B(n_1931),
.Y(n_2214)
);

AOI22xp33_ASAP7_75t_SL g2215 ( 
.A1(n_2135),
.A2(n_2055),
.B1(n_1936),
.B2(n_1958),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2115),
.B(n_1930),
.Y(n_2216)
);

AO21x2_ASAP7_75t_L g2217 ( 
.A1(n_2160),
.A2(n_1971),
.B(n_1877),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_2176),
.B(n_2052),
.Y(n_2218)
);

INVx1_ASAP7_75t_SL g2219 ( 
.A(n_2149),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2175),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2168),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_2073),
.Y(n_2222)
);

BUFx2_ASAP7_75t_L g2223 ( 
.A(n_2133),
.Y(n_2223)
);

INVxp67_ASAP7_75t_L g2224 ( 
.A(n_2086),
.Y(n_2224)
);

OR2x6_ASAP7_75t_L g2225 ( 
.A(n_2135),
.B(n_1875),
.Y(n_2225)
);

AOI22xp33_ASAP7_75t_L g2226 ( 
.A1(n_2167),
.A2(n_1994),
.B1(n_2056),
.B2(n_2033),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_2130),
.B(n_1958),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2147),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2152),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2151),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2119),
.Y(n_2231)
);

AND2x4_ASAP7_75t_L g2232 ( 
.A(n_2133),
.B(n_2052),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2119),
.Y(n_2233)
);

HB1xp67_ASAP7_75t_L g2234 ( 
.A(n_2065),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2151),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2095),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2117),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2123),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_2132),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_2114),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2141),
.Y(n_2241)
);

AND2x4_ASAP7_75t_L g2242 ( 
.A(n_2103),
.B(n_2155),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_2132),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2174),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2174),
.Y(n_2245)
);

INVx4_ASAP7_75t_L g2246 ( 
.A(n_2138),
.Y(n_2246)
);

AO21x1_ASAP7_75t_L g2247 ( 
.A1(n_2136),
.A2(n_2134),
.B(n_2120),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_2065),
.Y(n_2248)
);

INVx1_ASAP7_75t_SL g2249 ( 
.A(n_2114),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2069),
.B(n_2131),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2155),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_2126),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2098),
.B(n_2172),
.Y(n_2253)
);

OA21x2_ASAP7_75t_L g2254 ( 
.A1(n_2156),
.A2(n_2053),
.B(n_2059),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2161),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2161),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_2086),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_2144),
.B(n_2113),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2137),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2117),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2253),
.B(n_2169),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_R g2262 ( 
.A(n_2257),
.B(n_2068),
.Y(n_2262)
);

XOR2xp5_ASAP7_75t_L g2263 ( 
.A(n_2257),
.B(n_2087),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2181),
.B(n_2118),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2200),
.B(n_2064),
.Y(n_2265)
);

BUFx24_ASAP7_75t_SL g2266 ( 
.A(n_2226),
.Y(n_2266)
);

NAND2xp33_ASAP7_75t_R g2267 ( 
.A(n_2182),
.B(n_2093),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2195),
.B(n_2142),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2207),
.B(n_2144),
.Y(n_2269)
);

OR2x6_ASAP7_75t_L g2270 ( 
.A(n_2199),
.B(n_2148),
.Y(n_2270)
);

OR2x2_ASAP7_75t_L g2271 ( 
.A(n_2220),
.B(n_2113),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2187),
.B(n_2143),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2181),
.B(n_2150),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_2182),
.B(n_2142),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2204),
.B(n_2117),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2204),
.B(n_2150),
.Y(n_2276)
);

XOR2x2_ASAP7_75t_SL g2277 ( 
.A(n_2188),
.B(n_2066),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_R g2278 ( 
.A(n_2199),
.B(n_2085),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_R g2279 ( 
.A(n_2199),
.B(n_2085),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_2188),
.B(n_2079),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2205),
.B(n_2143),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2208),
.B(n_2066),
.Y(n_2282)
);

NAND2xp33_ASAP7_75t_R g2283 ( 
.A(n_2188),
.B(n_2089),
.Y(n_2283)
);

INVx4_ASAP7_75t_L g2284 ( 
.A(n_2246),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2229),
.B(n_2100),
.Y(n_2285)
);

NAND2xp33_ASAP7_75t_R g2286 ( 
.A(n_2239),
.B(n_2153),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2202),
.B(n_2170),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2189),
.B(n_2170),
.Y(n_2288)
);

OR2x6_ASAP7_75t_L g2289 ( 
.A(n_2246),
.B(n_2138),
.Y(n_2289)
);

NAND2xp33_ASAP7_75t_R g2290 ( 
.A(n_2239),
.B(n_2153),
.Y(n_2290)
);

BUFx3_ASAP7_75t_L g2291 ( 
.A(n_2241),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2234),
.B(n_2044),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2191),
.B(n_2075),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2192),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_R g2295 ( 
.A(n_2259),
.B(n_2088),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_2232),
.B(n_2079),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2248),
.B(n_2044),
.Y(n_2297)
);

OR2x6_ASAP7_75t_L g2298 ( 
.A(n_2246),
.B(n_2097),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_R g2299 ( 
.A(n_2239),
.B(n_2157),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_2250),
.B(n_2097),
.Y(n_2300)
);

INVxp67_ASAP7_75t_L g2301 ( 
.A(n_2222),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_R g2302 ( 
.A(n_2224),
.B(n_2126),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2193),
.B(n_2171),
.Y(n_2303)
);

BUFx3_ASAP7_75t_L g2304 ( 
.A(n_2252),
.Y(n_2304)
);

NAND2xp33_ASAP7_75t_R g2305 ( 
.A(n_2243),
.B(n_2223),
.Y(n_2305)
);

XNOR2xp5_ASAP7_75t_L g2306 ( 
.A(n_2240),
.B(n_2164),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_R g2307 ( 
.A(n_2243),
.B(n_2223),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2184),
.B(n_2044),
.Y(n_2308)
);

CKINVDCx11_ASAP7_75t_R g2309 ( 
.A(n_2219),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2244),
.B(n_2171),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2245),
.B(n_2173),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2215),
.B(n_2164),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_2232),
.B(n_2079),
.Y(n_2313)
);

OR2x6_ASAP7_75t_L g2314 ( 
.A(n_2228),
.B(n_2124),
.Y(n_2314)
);

NAND2xp33_ASAP7_75t_SL g2315 ( 
.A(n_2258),
.B(n_2243),
.Y(n_2315)
);

INVxp67_ASAP7_75t_L g2316 ( 
.A(n_2203),
.Y(n_2316)
);

XNOR2xp5_ASAP7_75t_L g2317 ( 
.A(n_2249),
.B(n_2124),
.Y(n_2317)
);

NAND2xp33_ASAP7_75t_R g2318 ( 
.A(n_2225),
.B(n_2157),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2211),
.B(n_1933),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_R g2320 ( 
.A(n_2178),
.B(n_2126),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2232),
.B(n_2145),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2230),
.B(n_2145),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2218),
.B(n_2242),
.Y(n_2323)
);

NAND2xp33_ASAP7_75t_R g2324 ( 
.A(n_2225),
.B(n_2165),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_2218),
.B(n_2078),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_R g2326 ( 
.A(n_2178),
.B(n_2051),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2294),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2303),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_SL g2329 ( 
.A1(n_2278),
.A2(n_2218),
.B1(n_2258),
.B2(n_2194),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2285),
.B(n_2235),
.Y(n_2330)
);

OR2x2_ASAP7_75t_L g2331 ( 
.A(n_2271),
.B(n_2180),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2310),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2293),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2322),
.Y(n_2334)
);

AOI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2283),
.A2(n_2196),
.B1(n_2214),
.B2(n_2247),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2323),
.B(n_2209),
.Y(n_2336)
);

NAND4xp25_ASAP7_75t_L g2337 ( 
.A(n_2312),
.B(n_1960),
.C(n_1900),
.D(n_2180),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2323),
.B(n_2209),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2292),
.B(n_2216),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2325),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2288),
.Y(n_2341)
);

BUFx3_ASAP7_75t_L g2342 ( 
.A(n_2289),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_SL g2343 ( 
.A1(n_2306),
.A2(n_2194),
.B(n_2190),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2297),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2321),
.B(n_2237),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2279),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2301),
.B(n_2177),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2275),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2263),
.B(n_2236),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2316),
.B(n_2238),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_2326),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2275),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2325),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2289),
.A2(n_2190),
.B1(n_2194),
.B2(n_2122),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2308),
.B(n_2216),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2321),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2269),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2265),
.B(n_2177),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2296),
.B(n_2231),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2282),
.A2(n_2247),
.B1(n_2217),
.B2(n_2214),
.Y(n_2360)
);

OAI22xp5_ASAP7_75t_L g2361 ( 
.A1(n_2284),
.A2(n_2122),
.B1(n_2225),
.B2(n_2179),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2281),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2272),
.B(n_2231),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_2362),
.B(n_2309),
.Y(n_2364)
);

AOI22xp33_ASAP7_75t_L g2365 ( 
.A1(n_2351),
.A2(n_2264),
.B1(n_2315),
.B2(n_2214),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2327),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2357),
.B(n_2233),
.Y(n_2367)
);

INVx3_ASAP7_75t_L g2368 ( 
.A(n_2346),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2357),
.B(n_2261),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2327),
.Y(n_2370)
);

NAND4xp25_ASAP7_75t_L g2371 ( 
.A(n_2335),
.B(n_2267),
.C(n_2262),
.D(n_2311),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2332),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2339),
.B(n_2296),
.Y(n_2373)
);

INVx1_ASAP7_75t_SL g2374 ( 
.A(n_2351),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2332),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2333),
.B(n_2183),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2339),
.B(n_2313),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2355),
.B(n_2313),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2328),
.Y(n_2379)
);

INVx2_ASAP7_75t_SL g2380 ( 
.A(n_2342),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2355),
.B(n_2260),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2334),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2331),
.B(n_2233),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2328),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2346),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2334),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2333),
.B(n_2183),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2336),
.B(n_2260),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2331),
.Y(n_2389)
);

NAND3xp33_ASAP7_75t_L g2390 ( 
.A(n_2335),
.B(n_2291),
.C(n_2270),
.Y(n_2390)
);

AOI221xp5_ASAP7_75t_L g2391 ( 
.A1(n_2360),
.A2(n_2295),
.B1(n_2287),
.B2(n_2319),
.C(n_2146),
.Y(n_2391)
);

AND2x2_ASAP7_75t_SL g2392 ( 
.A(n_2345),
.B(n_2280),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2336),
.B(n_2237),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2344),
.B(n_2213),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_2368),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2389),
.B(n_2341),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2381),
.B(n_2348),
.Y(n_2397)
);

OR2x2_ASAP7_75t_L g2398 ( 
.A(n_2389),
.B(n_2344),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2368),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2383),
.B(n_2347),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2381),
.B(n_2348),
.Y(n_2401)
);

OR2x2_ASAP7_75t_L g2402 ( 
.A(n_2383),
.B(n_2341),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2388),
.B(n_2352),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2372),
.Y(n_2404)
);

AND3x2_ASAP7_75t_L g2405 ( 
.A(n_2364),
.B(n_2349),
.C(n_2350),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2372),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2382),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2388),
.B(n_2352),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2378),
.B(n_2356),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2375),
.Y(n_2410)
);

A2O1A1Ixp33_ASAP7_75t_L g2411 ( 
.A1(n_2390),
.A2(n_2342),
.B(n_2343),
.C(n_2329),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2382),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2386),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2375),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2378),
.B(n_2373),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2379),
.B(n_2330),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2379),
.B(n_2358),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2386),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2366),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2384),
.B(n_2362),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2373),
.B(n_2356),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2377),
.B(n_2338),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2390),
.B(n_2340),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2366),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2384),
.B(n_2363),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2425),
.B(n_2374),
.Y(n_2426)
);

AOI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2411),
.A2(n_2371),
.B1(n_2391),
.B2(n_2368),
.Y(n_2427)
);

NAND2xp33_ASAP7_75t_SL g2428 ( 
.A(n_2395),
.B(n_2385),
.Y(n_2428)
);

OAI22xp33_ASAP7_75t_L g2429 ( 
.A1(n_2395),
.A2(n_2371),
.B1(n_2385),
.B2(n_2343),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_2399),
.Y(n_2430)
);

OAI221xp5_ASAP7_75t_L g2431 ( 
.A1(n_2399),
.A2(n_2365),
.B1(n_2385),
.B2(n_2380),
.C(n_2361),
.Y(n_2431)
);

AO221x2_ASAP7_75t_L g2432 ( 
.A1(n_2405),
.A2(n_2354),
.B1(n_2392),
.B2(n_2277),
.C(n_2425),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2420),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2416),
.B(n_2376),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2397),
.B(n_2387),
.Y(n_2435)
);

HB1xp67_ASAP7_75t_L g2436 ( 
.A(n_2404),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2397),
.B(n_2369),
.Y(n_2437)
);

NOR2xp33_ASAP7_75t_L g2438 ( 
.A(n_2396),
.B(n_2380),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2401),
.B(n_2370),
.Y(n_2439)
);

AND2x4_ASAP7_75t_L g2440 ( 
.A(n_2423),
.B(n_2415),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_2423),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_2423),
.Y(n_2442)
);

OAI221xp5_ASAP7_75t_L g2443 ( 
.A1(n_2417),
.A2(n_2337),
.B1(n_2363),
.B2(n_2307),
.C(n_2305),
.Y(n_2443)
);

NOR2x1_ASAP7_75t_L g2444 ( 
.A(n_2429),
.B(n_2270),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2430),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2440),
.B(n_2401),
.Y(n_2446)
);

INVx1_ASAP7_75t_SL g2447 ( 
.A(n_2426),
.Y(n_2447)
);

INVx1_ASAP7_75t_SL g2448 ( 
.A(n_2428),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2427),
.B(n_2402),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2440),
.B(n_2403),
.Y(n_2450)
);

AOI22xp33_ASAP7_75t_SL g2451 ( 
.A1(n_2432),
.A2(n_2423),
.B1(n_2392),
.B2(n_2302),
.Y(n_2451)
);

HB1xp67_ASAP7_75t_L g2452 ( 
.A(n_2436),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2433),
.B(n_2403),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2442),
.Y(n_2454)
);

INVx4_ASAP7_75t_L g2455 ( 
.A(n_2441),
.Y(n_2455)
);

NAND3xp33_ASAP7_75t_L g2456 ( 
.A(n_2432),
.B(n_2337),
.C(n_2082),
.Y(n_2456)
);

NAND2xp33_ASAP7_75t_SL g2457 ( 
.A(n_2441),
.B(n_2320),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2442),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2439),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2438),
.B(n_2408),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2434),
.B(n_2408),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2435),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2437),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2458),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2452),
.Y(n_2465)
);

O2A1O1Ixp33_ASAP7_75t_L g2466 ( 
.A1(n_2456),
.A2(n_2444),
.B(n_2445),
.C(n_2454),
.Y(n_2466)
);

XNOR2xp5_ASAP7_75t_L g2467 ( 
.A(n_2456),
.B(n_2443),
.Y(n_2467)
);

AOI21xp33_ASAP7_75t_L g2468 ( 
.A1(n_2455),
.A2(n_2431),
.B(n_1982),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2445),
.B(n_2398),
.Y(n_2469)
);

OAI32xp33_ASAP7_75t_L g2470 ( 
.A1(n_2455),
.A2(n_2398),
.A3(n_2402),
.B1(n_2400),
.B2(n_2415),
.Y(n_2470)
);

AOI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_2451),
.A2(n_2392),
.B1(n_2410),
.B2(n_2404),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2459),
.Y(n_2472)
);

NOR2x1p5_ASAP7_75t_L g2473 ( 
.A(n_2455),
.B(n_2400),
.Y(n_2473)
);

O2A1O1Ixp33_ASAP7_75t_L g2474 ( 
.A1(n_2444),
.A2(n_2129),
.B(n_2108),
.C(n_2102),
.Y(n_2474)
);

OAI21xp33_ASAP7_75t_L g2475 ( 
.A1(n_2449),
.A2(n_2448),
.B(n_2458),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2463),
.B(n_2422),
.Y(n_2476)
);

OAI222xp33_ASAP7_75t_L g2477 ( 
.A1(n_2447),
.A2(n_2317),
.B1(n_2298),
.B2(n_2422),
.C1(n_2314),
.C2(n_2377),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2473),
.B(n_2446),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2475),
.B(n_2463),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2469),
.B(n_2465),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2472),
.B(n_2462),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2467),
.B(n_2462),
.Y(n_2482)
);

NAND2x1_ASAP7_75t_L g2483 ( 
.A(n_2464),
.B(n_2446),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2476),
.Y(n_2484)
);

AOI22xp33_ASAP7_75t_L g2485 ( 
.A1(n_2468),
.A2(n_2457),
.B1(n_2459),
.B2(n_2450),
.Y(n_2485)
);

INVx1_ASAP7_75t_SL g2486 ( 
.A(n_2468),
.Y(n_2486)
);

NOR2xp67_ASAP7_75t_L g2487 ( 
.A(n_2471),
.B(n_2466),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2477),
.A2(n_2450),
.B1(n_2460),
.B2(n_2453),
.Y(n_2488)
);

NAND2x1_ASAP7_75t_SL g2489 ( 
.A(n_2470),
.B(n_2460),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2474),
.B(n_2461),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2465),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2480),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2478),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2491),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_2482),
.B(n_2490),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2483),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2479),
.B(n_2406),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2481),
.Y(n_2498)
);

INVxp33_ASAP7_75t_L g2499 ( 
.A(n_2489),
.Y(n_2499)
);

INVxp67_ASAP7_75t_L g2500 ( 
.A(n_2486),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2481),
.Y(n_2501)
);

CKINVDCx16_ASAP7_75t_R g2502 ( 
.A(n_2484),
.Y(n_2502)
);

INVx2_ASAP7_75t_SL g2503 ( 
.A(n_2485),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2488),
.Y(n_2504)
);

CKINVDCx6p67_ASAP7_75t_R g2505 ( 
.A(n_2487),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2480),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2480),
.Y(n_2507)
);

NAND4xp25_ASAP7_75t_L g2508 ( 
.A(n_2495),
.B(n_2112),
.C(n_2304),
.D(n_2104),
.Y(n_2508)
);

NOR4xp25_ASAP7_75t_L g2509 ( 
.A(n_2500),
.B(n_1895),
.C(n_2011),
.D(n_2003),
.Y(n_2509)
);

NOR4xp25_ASAP7_75t_L g2510 ( 
.A(n_2500),
.B(n_1899),
.C(n_1904),
.D(n_1928),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2504),
.B(n_2406),
.Y(n_2511)
);

NAND3xp33_ASAP7_75t_SL g2512 ( 
.A(n_2499),
.B(n_1959),
.C(n_1998),
.Y(n_2512)
);

OAI21xp33_ASAP7_75t_L g2513 ( 
.A1(n_2499),
.A2(n_2314),
.B(n_2409),
.Y(n_2513)
);

NOR4xp25_ASAP7_75t_L g2514 ( 
.A(n_2495),
.B(n_2025),
.C(n_2001),
.D(n_1974),
.Y(n_2514)
);

NOR2xp67_ASAP7_75t_L g2515 ( 
.A(n_2496),
.B(n_2410),
.Y(n_2515)
);

NAND3xp33_ASAP7_75t_SL g2516 ( 
.A(n_2492),
.B(n_2107),
.C(n_1937),
.Y(n_2516)
);

AOI211xp5_ASAP7_75t_L g2517 ( 
.A1(n_2503),
.A2(n_2102),
.B(n_2108),
.C(n_2074),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2493),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2505),
.B(n_2409),
.Y(n_2519)
);

OAI211xp5_ASAP7_75t_L g2520 ( 
.A1(n_2506),
.A2(n_2507),
.B(n_2498),
.C(n_2501),
.Y(n_2520)
);

NOR2xp67_ASAP7_75t_L g2521 ( 
.A(n_2496),
.B(n_2414),
.Y(n_2521)
);

NAND4xp75_ASAP7_75t_L g2522 ( 
.A(n_2494),
.B(n_2497),
.C(n_2502),
.D(n_1986),
.Y(n_2522)
);

OAI211xp5_ASAP7_75t_SL g2523 ( 
.A1(n_2497),
.A2(n_2107),
.B(n_1997),
.C(n_2136),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2504),
.B(n_2414),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2518),
.Y(n_2525)
);

AOI221xp5_ASAP7_75t_SL g2526 ( 
.A1(n_2511),
.A2(n_2421),
.B1(n_2266),
.B2(n_2424),
.C(n_2407),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2519),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_2524),
.Y(n_2528)
);

OAI21x1_ASAP7_75t_SL g2529 ( 
.A1(n_2522),
.A2(n_2520),
.B(n_2510),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2515),
.Y(n_2530)
);

AOI221xp5_ASAP7_75t_L g2531 ( 
.A1(n_2516),
.A2(n_2424),
.B1(n_2407),
.B2(n_2412),
.C(n_2413),
.Y(n_2531)
);

AOI221xp5_ASAP7_75t_L g2532 ( 
.A1(n_2514),
.A2(n_2407),
.B1(n_2412),
.B2(n_2413),
.C(n_2418),
.Y(n_2532)
);

AOI211xp5_ASAP7_75t_L g2533 ( 
.A1(n_2512),
.A2(n_1929),
.B(n_2134),
.C(n_2273),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2513),
.B(n_2421),
.Y(n_2534)
);

AOI221xp5_ASAP7_75t_L g2535 ( 
.A1(n_2509),
.A2(n_2418),
.B1(n_2412),
.B2(n_2413),
.C(n_2419),
.Y(n_2535)
);

OAI211xp5_ASAP7_75t_L g2536 ( 
.A1(n_2517),
.A2(n_2198),
.B(n_1993),
.C(n_1946),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2521),
.B(n_2418),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2508),
.Y(n_2538)
);

INVxp67_ASAP7_75t_SL g2539 ( 
.A(n_2525),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2527),
.Y(n_2540)
);

NAND4xp75_ASAP7_75t_L g2541 ( 
.A(n_2530),
.B(n_2523),
.C(n_1970),
.D(n_1951),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2538),
.A2(n_2318),
.B1(n_2324),
.B2(n_2298),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2538),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2538),
.B(n_2419),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2537),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2528),
.Y(n_2546)
);

XNOR2xp5_ASAP7_75t_L g2547 ( 
.A(n_2533),
.B(n_2300),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2526),
.B(n_2419),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2534),
.B(n_2536),
.Y(n_2549)
);

NAND3xp33_ASAP7_75t_L g2550 ( 
.A(n_2543),
.B(n_2531),
.C(n_2532),
.Y(n_2550)
);

NOR2xp67_ASAP7_75t_L g2551 ( 
.A(n_2546),
.B(n_2529),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2540),
.B(n_2535),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_R g2553 ( 
.A(n_2544),
.B(n_2252),
.Y(n_2553)
);

NAND2xp33_ASAP7_75t_SL g2554 ( 
.A(n_2545),
.B(n_2198),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_R g2555 ( 
.A(n_2549),
.B(n_2299),
.Y(n_2555)
);

NAND2xp33_ASAP7_75t_SL g2556 ( 
.A(n_2547),
.B(n_2039),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2539),
.B(n_2039),
.Y(n_2557)
);

NAND3xp33_ASAP7_75t_L g2558 ( 
.A(n_2542),
.B(n_1901),
.C(n_2039),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2541),
.B(n_2206),
.Y(n_2559)
);

NAND3xp33_ASAP7_75t_L g2560 ( 
.A(n_2542),
.B(n_2548),
.C(n_2041),
.Y(n_2560)
);

NAND2xp33_ASAP7_75t_SL g2561 ( 
.A(n_2543),
.B(n_2041),
.Y(n_2561)
);

OAI21x1_ASAP7_75t_L g2562 ( 
.A1(n_2543),
.A2(n_2159),
.B(n_2090),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2551),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_2550),
.Y(n_2564)
);

OAI22xp5_ASAP7_75t_SL g2565 ( 
.A1(n_2559),
.A2(n_2560),
.B1(n_2558),
.B2(n_2552),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2557),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2562),
.Y(n_2567)
);

AOI221xp5_ASAP7_75t_L g2568 ( 
.A1(n_2561),
.A2(n_2041),
.B1(n_1953),
.B2(n_2370),
.C(n_2120),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2553),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2554),
.Y(n_2570)
);

AOI221xp5_ASAP7_75t_L g2571 ( 
.A1(n_2556),
.A2(n_2555),
.B1(n_2094),
.B2(n_2255),
.C(n_2256),
.Y(n_2571)
);

OA22x2_ASAP7_75t_L g2572 ( 
.A1(n_2552),
.A2(n_2225),
.B1(n_2340),
.B2(n_2353),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2551),
.A2(n_2280),
.B1(n_2268),
.B2(n_2290),
.Y(n_2573)
);

OAI211xp5_ASAP7_75t_L g2574 ( 
.A1(n_2551),
.A2(n_2367),
.B(n_2353),
.C(n_2121),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_2562),
.Y(n_2575)
);

AOI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2551),
.A2(n_2268),
.B1(n_2286),
.B2(n_2217),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2564),
.B(n_2393),
.Y(n_2577)
);

OA21x2_ASAP7_75t_L g2578 ( 
.A1(n_2563),
.A2(n_2140),
.B(n_2105),
.Y(n_2578)
);

OA22x2_ASAP7_75t_L g2579 ( 
.A1(n_2569),
.A2(n_2206),
.B1(n_2345),
.B2(n_2276),
.Y(n_2579)
);

OAI31xp33_ASAP7_75t_L g2580 ( 
.A1(n_2566),
.A2(n_2090),
.A3(n_2227),
.B(n_2084),
.Y(n_2580)
);

INVx1_ASAP7_75t_SL g2581 ( 
.A(n_2570),
.Y(n_2581)
);

OAI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2573),
.A2(n_2367),
.B1(n_2394),
.B2(n_2227),
.Y(n_2582)
);

NOR3xp33_ASAP7_75t_SL g2583 ( 
.A(n_2565),
.B(n_2156),
.C(n_2210),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2575),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2575),
.Y(n_2585)
);

XNOR2xp5_ASAP7_75t_L g2586 ( 
.A(n_2567),
.B(n_2276),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2576),
.Y(n_2587)
);

OAI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2581),
.A2(n_2572),
.B(n_2571),
.Y(n_2588)
);

OAI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2586),
.A2(n_2574),
.B1(n_2568),
.B2(n_2394),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2584),
.Y(n_2590)
);

AOI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2577),
.A2(n_2585),
.B1(n_2587),
.B2(n_2579),
.Y(n_2591)
);

AOI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_2583),
.A2(n_2582),
.B1(n_2578),
.B2(n_2580),
.Y(n_2592)
);

XNOR2xp5_ASAP7_75t_L g2593 ( 
.A(n_2578),
.B(n_2084),
.Y(n_2593)
);

AOI31xp33_ASAP7_75t_L g2594 ( 
.A1(n_2581),
.A2(n_2227),
.A3(n_2274),
.B(n_2359),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2581),
.B(n_2345),
.Y(n_2595)
);

OAI211xp5_ASAP7_75t_L g2596 ( 
.A1(n_2581),
.A2(n_2393),
.B(n_2338),
.C(n_2359),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2584),
.Y(n_2597)
);

AOI22xp33_ASAP7_75t_L g2598 ( 
.A1(n_2597),
.A2(n_2345),
.B1(n_2217),
.B2(n_2274),
.Y(n_2598)
);

AOI31xp33_ASAP7_75t_L g2599 ( 
.A1(n_2590),
.A2(n_2212),
.A3(n_2024),
.B(n_2179),
.Y(n_2599)
);

AOI31xp33_ASAP7_75t_L g2600 ( 
.A1(n_2591),
.A2(n_2024),
.A3(n_2251),
.B(n_2047),
.Y(n_2600)
);

AOI31xp33_ASAP7_75t_L g2601 ( 
.A1(n_2588),
.A2(n_2592),
.A3(n_2595),
.B(n_2589),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_2593),
.A2(n_2256),
.B1(n_2255),
.B2(n_2254),
.Y(n_2602)
);

AOI31xp33_ASAP7_75t_L g2603 ( 
.A1(n_2596),
.A2(n_2024),
.A3(n_2251),
.B(n_2047),
.Y(n_2603)
);

AOI31xp33_ASAP7_75t_L g2604 ( 
.A1(n_2594),
.A2(n_2047),
.A3(n_2242),
.B(n_2201),
.Y(n_2604)
);

XNOR2x2_ASAP7_75t_L g2605 ( 
.A(n_2601),
.B(n_2116),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_SL g2606 ( 
.A1(n_2598),
.A2(n_2077),
.B1(n_2254),
.B2(n_2165),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2604),
.Y(n_2607)
);

AOI22xp33_ASAP7_75t_L g2608 ( 
.A1(n_2602),
.A2(n_2254),
.B1(n_2242),
.B2(n_2154),
.Y(n_2608)
);

OAI21x1_ASAP7_75t_L g2609 ( 
.A1(n_2603),
.A2(n_2599),
.B(n_2600),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2607),
.A2(n_1992),
.B(n_1903),
.Y(n_2610)
);

AOI222xp33_ASAP7_75t_L g2611 ( 
.A1(n_2606),
.A2(n_2185),
.B1(n_2186),
.B2(n_2221),
.C1(n_2197),
.C2(n_2201),
.Y(n_2611)
);

AOI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2609),
.A2(n_2605),
.B(n_2608),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2612),
.Y(n_2613)
);

OAI221xp5_ASAP7_75t_R g2614 ( 
.A1(n_2613),
.A2(n_2611),
.B1(n_2610),
.B2(n_2159),
.C(n_2162),
.Y(n_2614)
);

AOI211xp5_ASAP7_75t_L g2615 ( 
.A1(n_2614),
.A2(n_2221),
.B(n_2197),
.C(n_2186),
.Y(n_2615)
);


endmodule