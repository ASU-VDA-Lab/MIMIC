module fake_jpeg_31218_n_446 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_446);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_58),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_82),
.Y(n_98)
);

CKINVDCx11_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_59),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_70),
.Y(n_137)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_65),
.Y(n_134)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_79),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_30),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_84),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_16),
.B(n_14),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_86),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_35),
.B(n_0),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_29),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_90),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_29),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_28),
.B1(n_44),
.B2(n_31),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_95),
.A2(n_103),
.B1(n_104),
.B2(n_131),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_45),
.B(n_43),
.C(n_38),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_99),
.B(n_82),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_28),
.B1(n_44),
.B2(n_31),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_27),
.B1(n_46),
.B2(n_26),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_114),
.A2(n_136),
.B1(n_47),
.B2(n_62),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_36),
.B1(n_43),
.B2(n_38),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_121),
.B1(n_126),
.B2(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_45),
.B1(n_34),
.B2(n_32),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_120),
.A2(n_132),
.B1(n_64),
.B2(n_84),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_36),
.B1(n_34),
.B2(n_46),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_27),
.B1(n_26),
.B2(n_20),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_7),
.B(n_8),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_74),
.A2(n_33),
.B1(n_29),
.B2(n_4),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_81),
.A2(n_33),
.B1(n_29),
.B2(n_4),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_33),
.B1(n_29),
.B2(n_5),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_72),
.A2(n_33),
.B1(n_3),
.B2(n_5),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_80),
.A2(n_33),
.B1(n_3),
.B2(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_78),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_51),
.B1(n_73),
.B2(n_61),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_71),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_145),
.Y(n_221)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_149),
.B(n_153),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_55),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_150),
.B(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_97),
.A2(n_52),
.B(n_50),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_154),
.A2(n_156),
.B(n_10),
.C(n_11),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_98),
.A2(n_84),
.B(n_77),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_59),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_163),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_99),
.A2(n_91),
.B1(n_66),
.B2(n_69),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_122),
.B1(n_118),
.B2(n_112),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

BUFx16f_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_119),
.B(n_53),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_162),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_51),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_140),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_166),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_120),
.B1(n_124),
.B2(n_127),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_65),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

HAxp5_ASAP7_75t_SL g230 ( 
.A(n_170),
.B(n_187),
.CON(n_230),
.SN(n_230)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_54),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_173),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_97),
.B(n_7),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_48),
.Y(n_173)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_7),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_182),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_127),
.B1(n_125),
.B2(n_101),
.Y(n_199)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_77),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_135),
.B(n_48),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_179),
.B(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_180),
.Y(n_232)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_128),
.Y(n_182)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_188),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_107),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_8),
.Y(n_189)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_12),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_92),
.C(n_109),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_192),
.B(n_213),
.C(n_231),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_202),
.B1(n_206),
.B2(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_199),
.A2(n_200),
.B1(n_204),
.B2(n_185),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_125),
.B1(n_107),
.B2(n_142),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_110),
.B1(n_142),
.B2(n_116),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_110),
.B1(n_116),
.B2(n_92),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_96),
.B1(n_109),
.B2(n_112),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_132),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_122),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_12),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_220),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_147),
.A2(n_10),
.B1(n_11),
.B2(n_166),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_179),
.B1(n_169),
.B2(n_151),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_145),
.B(n_11),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_177),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_156),
.B(n_154),
.Y(n_231)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_235),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_144),
.B1(n_170),
.B2(n_178),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_249),
.B1(n_250),
.B2(n_259),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_239),
.A2(n_198),
.B1(n_224),
.B2(n_203),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_161),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_240),
.B(n_243),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_207),
.B(n_178),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_148),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_148),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_244),
.B(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_148),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_246),
.A2(n_266),
.B1(n_268),
.B2(n_195),
.Y(n_305)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_161),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_248),
.B(n_251),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_207),
.A2(n_146),
.B1(n_157),
.B2(n_188),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_209),
.A2(n_155),
.B1(n_186),
.B2(n_180),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_161),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_254),
.B(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_209),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_181),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_264),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_155),
.B1(n_186),
.B2(n_165),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_205),
.A2(n_187),
.B1(n_143),
.B2(n_190),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_261),
.A2(n_233),
.B1(n_194),
.B2(n_193),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_196),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_263),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_152),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_202),
.A2(n_174),
.B1(n_184),
.B2(n_158),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_205),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_270),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_219),
.A2(n_192),
.B1(n_230),
.B2(n_211),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_211),
.B(n_226),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_233),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_222),
.B(n_215),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_273),
.A2(n_281),
.B(n_287),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_215),
.B(n_201),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_232),
.C(n_198),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_270),
.C(n_238),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_284),
.B(n_303),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_197),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_286),
.B(n_294),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_241),
.B(n_258),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_237),
.A2(n_193),
.B(n_194),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_217),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_214),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_305),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_249),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_236),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_301),
.B1(n_246),
.B2(n_259),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_206),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_298),
.B(n_224),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_262),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_238),
.C(n_252),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_308),
.Y(n_355)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_332),
.B1(n_334),
.B2(n_295),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_261),
.C(n_239),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_250),
.C(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_247),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_325),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_236),
.B1(n_242),
.B2(n_255),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_317),
.A2(n_274),
.B1(n_300),
.B2(n_290),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_271),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_333),
.C(n_281),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_260),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_321),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_299),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_322),
.B(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_327),
.A2(n_302),
.B1(n_235),
.B2(n_304),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_264),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_329),
.A2(n_334),
.B(n_314),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_290),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_330),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_253),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_195),
.C(n_203),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_254),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_280),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_316),
.A2(n_291),
.B1(n_288),
.B2(n_289),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_344),
.B1(n_350),
.B2(n_358),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_340),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_287),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_273),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_346),
.Y(n_381)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_317),
.A2(n_324),
.B1(n_319),
.B2(n_329),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_306),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_348),
.C(n_352),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_274),
.C(n_304),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_315),
.Y(n_364)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_292),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_295),
.C(n_296),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_333),
.C(n_330),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_324),
.A2(n_329),
.B1(n_311),
.B2(n_320),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_321),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_329),
.A2(n_302),
.B(n_296),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_361),
.B(n_326),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_356),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_371),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_359),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_364),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_345),
.Y(n_366)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_374),
.Y(n_398)
);

BUFx12_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_356),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_309),
.Y(n_375)
);

OAI21x1_ASAP7_75t_L g392 ( 
.A1(n_375),
.A2(n_380),
.B(n_308),
.Y(n_392)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_376),
.A2(n_378),
.B(n_379),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_355),
.Y(n_379)
);

BUFx12_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_347),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_342),
.C(n_348),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_390),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_395),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_373),
.A2(n_351),
.B1(n_352),
.B2(n_336),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_364),
.A2(n_358),
.B1(n_344),
.B2(n_354),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_387),
.A2(n_389),
.B1(n_378),
.B2(n_365),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_367),
.A2(n_342),
.B1(n_325),
.B2(n_339),
.Y(n_389)
);

INVx11_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_341),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_340),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_381),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_323),
.C(n_300),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_383),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_366),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_374),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_406),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_412),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_376),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_393),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_407),
.B(n_409),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_371),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_371),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_410),
.B(n_411),
.Y(n_419)
);

AOI22x1_ASAP7_75t_L g414 ( 
.A1(n_400),
.A2(n_384),
.B1(n_365),
.B2(n_380),
.Y(n_414)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_414),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_400),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_418),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_390),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_420),
.B(n_327),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_406),
.B(n_385),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_421),
.B(n_402),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_387),
.B1(n_397),
.B2(n_372),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_404),
.C(n_412),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_425),
.B(n_427),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_419),
.A2(n_403),
.B(n_386),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_430),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_416),
.A2(n_380),
.B(n_323),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_429),
.B(n_432),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_389),
.C(n_396),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_422),
.B(n_381),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_431),
.B(n_420),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_435),
.Y(n_441)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_424),
.A2(n_415),
.A3(n_414),
.B1(n_417),
.B2(n_395),
.C1(n_368),
.C2(n_235),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_426),
.B(n_217),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_438),
.B(n_432),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_439),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_437),
.Y(n_440)
);

AOI21x1_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_442),
.B(n_436),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_433),
.A2(n_430),
.B(n_436),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_441),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_444),
.Y(n_446)
);


endmodule