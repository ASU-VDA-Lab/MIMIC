module real_jpeg_32278_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_0),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_0),
.B(n_82),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_0),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_0),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_0),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_0),
.B(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_2),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_2),
.B(n_162),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_2),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_2),
.B(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_2),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_2),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_3),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_3),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_3),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_3),
.B(n_198),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_507),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_4),
.B(n_508),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_8),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_8),
.B(n_137),
.Y(n_136)
);

NAND2x1_ASAP7_75t_L g161 ( 
.A(n_8),
.B(n_162),
.Y(n_161)
);

NAND2x1p5_ASAP7_75t_L g194 ( 
.A(n_8),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_9),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_9),
.B(n_50),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_9),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_9),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_9),
.B(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_9),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_9),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_10),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_10),
.B(n_104),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_10),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_10),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_10),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_10),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_10),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_11),
.B(n_87),
.Y(n_236)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_11),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_11),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_11),
.B(n_378),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_11),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_12),
.Y(n_309)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_15),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_16),
.Y(n_246)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_16),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_17),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_17),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_17),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_17),
.B(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_17),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_17),
.B(n_499),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_473),
.Y(n_19)
);

OAI21x1_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_201),
.B(n_471),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_167),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_23),
.B(n_167),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_95),
.C(n_128),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_25),
.B(n_96),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_66),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_26),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_40),
.B(n_65),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_27),
.B(n_41),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_36),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_30),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_35),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_35),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_35),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_36),
.B(n_100),
.C(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_36),
.A2(n_37),
.B1(n_235),
.B2(n_236),
.Y(n_338)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_37),
.B(n_194),
.C(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_39),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_39),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_54),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_54),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B(n_53),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_43),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_43),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_43),
.A2(n_146),
.B1(n_274),
.B2(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_45),
.Y(n_366)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_45),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_46),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_92),
.C(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_64),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g447 ( 
.A1(n_46),
.A2(n_64),
.B1(n_364),
.B2(n_448),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_47),
.Y(n_437)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_52),
.Y(n_502)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_53),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_54),
.Y(n_253)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_61),
.B(n_155),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_63),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_64),
.B(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_84),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_67),
.B(n_169),
.C(n_170),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.C(n_80),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_68),
.B(n_165),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.C(n_75),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_69),
.A2(n_75),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_69),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_69),
.A2(n_133),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_69),
.B(n_183),
.C(n_489),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_71),
.B(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_73),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_78),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_78),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_89),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_80),
.A2(n_81),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_81),
.B(n_86),
.C(n_90),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_92),
.B(n_119),
.C(n_122),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_116),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_115),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_98),
.B(n_115),
.C(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_103),
.B(n_106),
.C(n_109),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_114),
.Y(n_105)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_136),
.C(n_140),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_106),
.A2(n_114),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_113),
.Y(n_285)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_119),
.A2(n_192),
.B1(n_193),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_119),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_119),
.B(n_278),
.C(n_281),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_119),
.A2(n_196),
.B1(n_281),
.B2(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_120),
.Y(n_384)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_121),
.Y(n_241)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_121),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_124),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_128),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_147),
.C(n_163),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_130),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.C(n_143),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_131),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_135),
.A2(n_143),
.B1(n_144),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_135),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_136),
.B(n_140),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_136),
.A2(n_192),
.B1(n_193),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_136),
.Y(n_504)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_147),
.A2(n_148),
.B1(n_163),
.B2(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_157),
.C(n_161),
.Y(n_148)
);

XOR2x2_ASAP7_75t_L g249 ( 
.A(n_149),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_155),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_152),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_155),
.B(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx4_ASAP7_75t_SL g276 ( 
.A(n_156),
.Y(n_276)
);

INVx8_ASAP7_75t_L g405 ( 
.A(n_156),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_158),
.B(n_161),
.Y(n_250)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_168),
.B(n_186),
.C(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_172),
.Y(n_476)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_185),
.Y(n_172)
);

XOR2x1_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_184),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_174),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g489 ( 
.A(n_175),
.Y(n_489)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_184),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_185),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_197),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_192),
.B(n_196),
.C(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_193),
.B(n_338),
.Y(n_337)
);

BUFx4f_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_197),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_465),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_294),
.C(n_459),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_257),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g465 ( 
.A1(n_205),
.A2(n_258),
.B(n_466),
.C(n_469),
.D(n_470),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_255),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_206),
.B(n_255),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.C(n_251),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_208),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_252),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_231),
.C(n_247),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_266),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_221),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g342 ( 
.A(n_213),
.B(n_343),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_215),
.A2(n_216),
.B1(n_221),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_216),
.A2(n_217),
.B(n_218),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_221),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.C(n_228),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_222),
.A2(n_223),
.B1(n_228),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AO22x2_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_233),
.B1(n_248),
.B2(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_242),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_234),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_237),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_291)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_241),
.Y(n_413)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_292),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_259),
.B(n_292),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.C(n_267),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g464 ( 
.A(n_261),
.B(n_265),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_267),
.B(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_286),
.C(n_290),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_268),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.C(n_277),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_272),
.A2(n_273),
.B1(n_277),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2x1p5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_350),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_340),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_296),
.B(n_340),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.C(n_323),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_324),
.Y(n_353)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.C(n_320),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_302),
.B(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_320),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.C(n_317),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_306),
.B(n_388),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_309),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_310),
.A2(n_311),
.B1(n_317),
.B2(n_318),
.Y(n_388)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_312),
.B(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_336),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_346),
.C(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.C(n_332),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_333),
.Y(n_369)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_348),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_342),
.B(n_348),
.C(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_345),
.Y(n_462)
);

AOI21x1_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_370),
.B(n_458),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_352),
.B(n_354),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.C(n_367),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_368),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.C(n_363),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_359),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_405),
.Y(n_416)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

BUFx4f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_391),
.B(n_457),
.Y(n_370)
);

NOR2x1_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_389),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_372),
.B(n_389),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.C(n_385),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_374),
.B(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_376),
.A2(n_386),
.B1(n_387),
.B2(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_376),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_380),
.C(n_382),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_377),
.B(n_380),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_382),
.B(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_451),
.B(n_456),
.Y(n_391)
);

OAI21x1_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_439),
.B(n_450),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_420),
.B(n_438),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_406),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_406),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_397),
.A2(n_398),
.B1(n_402),
.B2(n_403),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_397),
.B(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_414),
.B2(n_415),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_412),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_412),
.C(n_414),
.Y(n_449)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_417),
.Y(n_445)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_432),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_431),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_423),
.A2(n_431),
.B(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_449),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_449),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_444),
.C(n_447),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_453),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

AOI21x1_ASAP7_75t_L g466 ( 
.A1(n_460),
.A2(n_467),
.B(n_468),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_463),
.Y(n_467)
);

HB1xp67_ASAP7_75t_SL g471 ( 
.A(n_472),
.Y(n_471)
);

OAI21xp33_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_477),
.B(n_505),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_475),
.B(n_478),
.Y(n_506)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_483),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.C(n_482),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_494),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_488),
.B1(n_490),
.B2(n_493),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_490),
.Y(n_493)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_497),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_503),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);


endmodule