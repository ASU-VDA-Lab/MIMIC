module real_jpeg_13879_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_32),
.B1(n_36),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_4),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_4),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_40),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_55),
.C(n_58),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_56),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_32),
.C(n_67),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_23),
.C(n_35),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_4),
.B(n_191),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_32),
.B1(n_36),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_42),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_6),
.A2(n_42),
.B1(n_57),
.B2(n_58),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_27),
.B1(n_32),
.B2(n_36),
.Y(n_74)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_102),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_100),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_86),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_14),
.B(n_86),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_62),
.C(n_76),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_44),
.B2(n_61),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_16),
.A2(n_45),
.B(n_60),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_28),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_18),
.A2(n_45),
.B1(n_46),
.B2(n_60),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_18),
.A2(n_28),
.B1(n_60),
.B2(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_21),
.A2(n_22),
.B1(n_80),
.B2(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_21),
.B(n_40),
.Y(n_199)
);

AO22x1_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_24),
.B1(n_33),
.B2(n_35),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_24),
.B(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_30),
.A2(n_37),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OA21x2_ASAP7_75t_L g81 ( 
.A1(n_30),
.A2(n_37),
.B(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_37),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OA22x2_ASAP7_75t_SL g69 ( 
.A1(n_32),
.A2(n_36),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_32),
.B(n_186),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_40),
.B(n_43),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_46),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_45),
.A2(n_46),
.B1(n_64),
.B2(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_45),
.A2(n_46),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

AOI211xp5_ASAP7_75t_SL g155 ( 
.A1(n_45),
.A2(n_81),
.B(n_85),
.C(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_64),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_49),
.B(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_56),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_58),
.B(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_75),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_64),
.A2(n_81),
.B1(n_83),
.B2(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_64),
.B(n_131),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_64),
.A2(n_131),
.B(n_168),
.C(n_173),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_64),
.A2(n_83),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_69),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_88),
.B1(n_89),
.B2(n_98),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_77),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_82),
.B(n_84),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_81),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_81),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_81),
.A2(n_114),
.B1(n_131),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_81),
.A2(n_131),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_81),
.A2(n_131),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_81),
.A2(n_131),
.B1(n_185),
.B2(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_81),
.B(n_139),
.C(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_81),
.B(n_175),
.C(n_179),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_84),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_82),
.A2(n_84),
.B(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_139),
.C(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_99),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_121),
.B(n_222),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_117),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_105),
.B(n_117),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_110),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_107),
.A2(n_108),
.B1(n_135),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_141),
.B(n_221),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_123),
.B(n_125),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_133),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_219)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_133),
.A2(n_134),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_140),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_140),
.B1(n_150),
.B2(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_139),
.B(n_170),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_139),
.A2(n_140),
.B1(n_188),
.B2(n_192),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_139),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_140),
.B(n_201),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_162),
.B(n_215),
.C(n_220),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_152),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_144),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_145),
.A2(n_146),
.B1(n_168),
.B2(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_154),
.B(n_158),
.C(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_209),
.B(n_214),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_181),
.B(n_208),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_204),
.B(n_207),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_193),
.B(n_203),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_213),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);


endmodule