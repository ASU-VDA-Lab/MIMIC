module fake_jpeg_18920_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_32),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_33),
.B1(n_22),
.B2(n_19),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_33),
.B1(n_23),
.B2(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_57),
.B1(n_42),
.B2(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_51),
.Y(n_64)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_2),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_33),
.B1(n_21),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_58),
.B1(n_41),
.B2(n_24),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_21),
.B1(n_16),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_56),
.B1(n_37),
.B2(n_40),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_26),
.B1(n_31),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_37),
.B1(n_38),
.B2(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_70),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_40),
.C(n_42),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_54),
.C(n_5),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_93),
.B1(n_4),
.B2(n_5),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_42),
.B1(n_37),
.B2(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_73),
.B1(n_78),
.B2(n_80),
.Y(n_104)
);

XNOR2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_5),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_75),
.Y(n_118)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_41),
.B(n_35),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_87),
.B(n_89),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_39),
.B1(n_36),
.B2(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_39),
.B1(n_30),
.B2(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_84),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_36),
.A3(n_16),
.B1(n_25),
.B2(n_29),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_3),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_25),
.B1(n_28),
.B2(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_28),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_20),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_41),
.B1(n_32),
.B2(n_20),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_10),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_47),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_86),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_82),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_76),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_111),
.B1(n_114),
.B2(n_117),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_10),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_6),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_9),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_9),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_72),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_93),
.B1(n_69),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_130),
.B1(n_100),
.B2(n_107),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_63),
.B1(n_66),
.B2(n_78),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_72),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_134),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_140),
.B1(n_144),
.B2(n_102),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_112),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_108),
.C(n_101),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_103),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_145),
.B(n_120),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_141),
.B(n_116),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_74),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_92),
.B1(n_95),
.B2(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_119),
.B(n_118),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_68),
.B1(n_91),
.B2(n_79),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_68),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_61),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_118),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_143),
.B(n_120),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_156),
.B(n_163),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_157),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_155),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_170),
.B1(n_169),
.B2(n_153),
.C(n_156),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_116),
.C(n_115),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_115),
.C(n_98),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_111),
.C(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_167),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_144),
.B1(n_133),
.B2(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

XOR2x2_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_102),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_85),
.B(n_87),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_165),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_128),
.A2(n_136),
.B(n_147),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_125),
.B1(n_123),
.B2(n_128),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_124),
.B1(n_170),
.B2(n_165),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_161),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_188),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_146),
.A3(n_124),
.B1(n_126),
.B2(n_113),
.C1(n_14),
.C2(n_10),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_70),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_163),
.B(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_159),
.C(n_168),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_160),
.C(n_181),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_163),
.B(n_149),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_203),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_162),
.B1(n_155),
.B2(n_157),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_174),
.B1(n_176),
.B2(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_168),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_204),
.B(n_186),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_172),
.B(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_212),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_204),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_213),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_175),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_182),
.C(n_171),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_217),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_203),
.C(n_197),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_187),
.B1(n_180),
.B2(n_173),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_210),
.C(n_223),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_202),
.C(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_222),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_208),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_190),
.B(n_191),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_190),
.B(n_195),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_212),
.C(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_210),
.C(n_211),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_233),
.Y(n_238)
);

OAI321xp33_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_196),
.A3(n_221),
.B1(n_214),
.B2(n_195),
.C(n_180),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_181),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_221),
.B(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_236),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_194),
.B1(n_184),
.B2(n_13),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_11),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_235),
.B(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_238),
.B(n_13),
.C(n_14),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_12),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_75),
.C(n_71),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_245),
.B1(n_12),
.B2(n_71),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_12),
.Y(n_247)
);


endmodule