module fake_jpeg_21435_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_22),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_21),
.B1(n_10),
.B2(n_4),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_10),
.B(n_11),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_20),
.B(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_40),
.B1(n_19),
.B2(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_29),
.B(n_25),
.Y(n_42)
);

NAND5xp2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_24),
.C(n_14),
.D(n_17),
.E(n_11),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_32),
.C(n_27),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_39),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_36),
.C(n_34),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_36),
.B1(n_38),
.B2(n_35),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_19),
.C(n_26),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_26),
.C(n_17),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_45),
.B(n_6),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_45),
.Y(n_51)
);

AOI322xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.A3(n_0),
.B1(n_8),
.B2(n_14),
.C1(n_46),
.C2(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_52),
.B(n_8),
.Y(n_53)
);


endmodule