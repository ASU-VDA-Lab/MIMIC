module fake_jpeg_12120_n_65 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_65);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_65;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_8),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_1),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_28)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_24),
.A2(n_12),
.B1(n_17),
.B2(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_14),
.B(n_13),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_28),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_17),
.B1(n_11),
.B2(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_16),
.B1(n_22),
.B2(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_20),
.C(n_19),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_1),
.C(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_22),
.B1(n_18),
.B2(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_39),
.B1(n_26),
.B2(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_37),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_43),
.B1(n_34),
.B2(n_36),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_18),
.C(n_3),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.C(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_52),
.B1(n_43),
.B2(n_42),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_38),
.B(n_34),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_46),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_56),
.C(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_4),
.Y(n_58)
);

XNOR2x1_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_50),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_48),
.B(n_50),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.C(n_59),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_54),
.C(n_56),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_8),
.C(n_6),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B(n_6),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

BUFx24_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);


endmodule