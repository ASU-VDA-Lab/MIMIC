module fake_jpeg_25117_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_35),
.B1(n_33),
.B2(n_17),
.Y(n_58)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_34),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_55),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_50),
.B(n_51),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_38),
.B1(n_33),
.B2(n_35),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_29),
.B1(n_44),
.B2(n_39),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_102),
.B1(n_35),
.B2(n_33),
.Y(n_111)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_70),
.Y(n_116)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_72),
.B(n_96),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_95),
.Y(n_108)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_26),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_88),
.Y(n_121)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_91),
.B1(n_33),
.B2(n_23),
.Y(n_112)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_26),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_28),
.B1(n_23),
.B2(n_29),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_103),
.Y(n_124)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_97),
.B1(n_87),
.B2(n_77),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_115),
.B1(n_123),
.B2(n_27),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_44),
.B1(n_39),
.B2(n_45),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_55),
.C(n_36),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_126),
.C(n_65),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_46),
.B1(n_28),
.B2(n_27),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_36),
.C(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_36),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_36),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_0),
.B(n_1),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_36),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_136),
.B(n_142),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_86),
.B1(n_69),
.B2(n_94),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_139),
.B1(n_149),
.B2(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_21),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_143),
.Y(n_169)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_151),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_126),
.B1(n_115),
.B2(n_116),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_71),
.B1(n_82),
.B2(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_41),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_158),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_155),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_43),
.C(n_80),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_27),
.B1(n_78),
.B2(n_76),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_166),
.B1(n_21),
.B2(n_122),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_88),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_157),
.B(n_22),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_42),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_42),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_163),
.B1(n_120),
.B2(n_125),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_165),
.B(n_21),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_105),
.B(n_75),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_107),
.A2(n_134),
.B1(n_84),
.B2(n_106),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_43),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_15),
.C(n_14),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_112),
.A2(n_59),
.B1(n_34),
.B2(n_17),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_106),
.B1(n_120),
.B2(n_125),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_175),
.B1(n_140),
.B2(n_148),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_134),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_198),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_179),
.B1(n_183),
.B2(n_186),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_1),
.B(n_2),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_166),
.B(n_3),
.Y(n_209)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_185),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_133),
.B1(n_129),
.B2(n_113),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_113),
.B1(n_133),
.B2(n_122),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_182),
.B(n_13),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_136),
.B1(n_145),
.B2(n_151),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_67),
.B1(n_99),
.B2(n_34),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_109),
.B1(n_17),
.B2(n_16),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_194),
.B1(n_196),
.B2(n_142),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_199),
.Y(n_205)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_24),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_141),
.A2(n_16),
.B1(n_25),
.B2(n_20),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_25),
.B1(n_20),
.B2(n_18),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_31),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_31),
.C(n_22),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_200),
.B(n_138),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_153),
.C(n_159),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_199),
.C(n_178),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_219),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_161),
.B1(n_158),
.B2(n_147),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_208),
.B1(n_211),
.B2(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_210),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_209),
.B(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_152),
.B1(n_31),
.B2(n_22),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_214),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_31),
.B(n_22),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_215),
.B(n_221),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_15),
.B(n_13),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_32),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_15),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_31),
.B(n_22),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_223),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_168),
.A2(n_189),
.B1(n_193),
.B2(n_181),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_193),
.A2(n_24),
.B1(n_32),
.B2(n_7),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_187),
.B1(n_191),
.B2(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_32),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_238),
.C(n_239),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_235),
.A2(n_245),
.B1(n_203),
.B2(n_231),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_236),
.B(n_244),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_178),
.C(n_190),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_198),
.C(n_181),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_169),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_201),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_185),
.B1(n_180),
.B2(n_194),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_173),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_177),
.C(n_196),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_251),
.C(n_253),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_180),
.C(n_32),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_32),
.C(n_24),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_243),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_256),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_206),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_261),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_252),
.B1(n_250),
.B2(n_210),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_259),
.B(n_11),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_202),
.B(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_204),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_221),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_213),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_269),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_272),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_231),
.A2(n_208),
.B1(n_216),
.B2(n_203),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_275),
.B1(n_258),
.B2(n_247),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_211),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_209),
.B1(n_227),
.B2(n_24),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_238),
.C(n_230),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_261),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_246),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_257),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_251),
.C(n_236),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_273),
.C(n_255),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_233),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_264),
.A2(n_11),
.B(n_13),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_290),
.A2(n_6),
.B(n_8),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_282),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_299),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_303),
.Y(n_309)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_273),
.B1(n_269),
.B2(n_263),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_306),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_263),
.C(n_8),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_276),
.C(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_279),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_6),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_292),
.B(n_291),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_308),
.B(n_310),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_288),
.B(n_281),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_281),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_277),
.C(n_282),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_318),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_302),
.B1(n_294),
.B2(n_283),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_317),
.B(n_293),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_307),
.B(n_305),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_315),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_322),
.B(n_296),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_296),
.B1(n_277),
.B2(n_9),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_310),
.B1(n_316),
.B2(n_314),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_327),
.A2(n_331),
.B(n_324),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.C(n_329),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_325),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_321),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_323),
.B(n_308),
.C(n_9),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_6),
.C(n_8),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_9),
.C(n_10),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_10),
.B(n_243),
.Y(n_339)
);


endmodule