module fake_jpeg_3658_n_493 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_493);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_493;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_16),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_63),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_9),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_67),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g154 ( 
.A(n_66),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_68),
.B(n_69),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_82),
.B(n_85),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_0),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_30),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_89),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_26),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_92),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_29),
.B(n_10),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_10),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g140 ( 
.A(n_97),
.Y(n_140)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_38),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_116),
.B(n_119),
.Y(n_178)
);

INVx2_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_118),
.B(n_90),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_86),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_121),
.A2(n_129),
.B(n_0),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_59),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_126),
.B(n_127),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_61),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_45),
.B(n_38),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_50),
.B(n_30),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_66),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_60),
.A2(n_80),
.B1(n_76),
.B2(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_171)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_55),
.A2(n_37),
.B1(n_35),
.B2(n_45),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_33),
.B1(n_40),
.B2(n_84),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_56),
.Y(n_151)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_157),
.B(n_145),
.Y(n_240)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_158),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_89),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_160),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_87),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_174),
.Y(n_222)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_54),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_188),
.Y(n_228)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_111),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_191),
.B1(n_204),
.B2(n_118),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_87),
.C(n_62),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_176),
.C(n_202),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_173),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_43),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_35),
.B(n_37),
.C(n_23),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_175),
.A2(n_197),
.B(n_208),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_106),
.B(n_64),
.C(n_98),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_33),
.B1(n_40),
.B2(n_43),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_179),
.A2(n_194),
.B1(n_200),
.B2(n_207),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_115),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_181),
.B(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_187),
.B1(n_199),
.B2(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_81),
.B1(n_27),
.B2(n_46),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_96),
.B1(n_32),
.B2(n_91),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_27),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_193),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_128),
.A2(n_46),
.B1(n_99),
.B2(n_18),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_140),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_201),
.Y(n_236)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_99),
.B1(n_32),
.B2(n_36),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_122),
.A2(n_36),
.B1(n_18),
.B2(n_49),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_119),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_101),
.B(n_96),
.C(n_83),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_104),
.A2(n_32),
.B1(n_36),
.B2(n_28),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_32),
.B1(n_28),
.B2(n_2),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_142),
.A2(n_32),
.B1(n_58),
.B2(n_28),
.Y(n_207)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_131),
.B(n_1),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_1),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_214),
.B(n_234),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_110),
.B1(n_104),
.B2(n_105),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_218),
.A2(n_241),
.B1(n_252),
.B2(n_255),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_221),
.B(n_206),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_238),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_174),
.A2(n_124),
.B1(n_102),
.B2(n_156),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_116),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_161),
.A2(n_117),
.B(n_152),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_251),
.B(n_202),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_246),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_184),
.A2(n_108),
.B1(n_143),
.B2(n_141),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_193),
.B(n_115),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_172),
.B(n_120),
.C(n_110),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_190),
.C(n_198),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_162),
.B(n_176),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_191),
.A2(n_153),
.B1(n_143),
.B2(n_141),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_108),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_175),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_189),
.A2(n_153),
.B1(n_138),
.B2(n_120),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_163),
.B(n_11),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_256),
.B(n_181),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_258),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_259),
.B(n_264),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_260),
.A2(n_285),
.B(n_295),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_226),
.A2(n_204),
.B(n_164),
.C(n_168),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_261),
.A2(n_216),
.B(n_244),
.C(n_230),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_262),
.Y(n_320)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_263),
.Y(n_331)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_169),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_177),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_269),
.B(n_279),
.Y(n_327)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_245),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_281),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_195),
.B1(n_190),
.B2(n_177),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_275),
.A2(n_212),
.B1(n_247),
.B2(n_254),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_188),
.Y(n_276)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_294),
.C(n_251),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_167),
.Y(n_279)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_280),
.Y(n_306)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_243),
.B(n_188),
.Y(n_281)
);

BUFx4f_ASAP7_75t_SL g282 ( 
.A(n_217),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_217),
.A2(n_225),
.B1(n_227),
.B2(n_242),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_220),
.B(n_170),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_210),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_289),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_235),
.B(n_209),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_288),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_180),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_239),
.A2(n_12),
.B1(n_17),
.B2(n_15),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_234),
.B1(n_242),
.B2(n_250),
.Y(n_308)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_223),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_1),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_228),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_182),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_246),
.B(n_11),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_214),
.A2(n_182),
.B1(n_5),
.B2(n_7),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_4),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_298),
.B(n_304),
.C(n_319),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_232),
.B1(n_252),
.B2(n_218),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_300),
.A2(n_307),
.B1(n_330),
.B2(n_291),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_301),
.B(n_328),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_238),
.C(n_235),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_305),
.B(n_294),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_240),
.B1(n_212),
.B2(n_215),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_315),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_272),
.A2(n_245),
.B(n_244),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_310),
.A2(n_321),
.B(n_329),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_249),
.C(n_247),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_260),
.A2(n_249),
.B(n_233),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_266),
.A2(n_233),
.B(n_230),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_270),
.A2(n_215),
.B1(n_11),
.B2(n_13),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_266),
.A2(n_17),
.B1(n_5),
.B2(n_7),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_333),
.A2(n_267),
.B1(n_282),
.B2(n_274),
.Y(n_362)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_359),
.Y(n_380)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_311),
.Y(n_339)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_279),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_340),
.B(n_341),
.C(n_342),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_269),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_259),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_265),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_344),
.B(n_348),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_SL g345 ( 
.A(n_303),
.B(n_287),
.C(n_264),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_346),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_277),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_293),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_351),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_271),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_303),
.A2(n_261),
.B(n_296),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_350),
.A2(n_321),
.B(n_315),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_322),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_352),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_282),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_358),
.Y(n_375)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_297),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_355),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_357),
.B(n_318),
.Y(n_392)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_302),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_361),
.Y(n_368)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_363),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_292),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_334),
.B(n_278),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_332),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_267),
.B1(n_297),
.B2(n_281),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_365),
.A2(n_300),
.B1(n_330),
.B2(n_326),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_298),
.C(n_319),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_340),
.C(n_337),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_338),
.B1(n_349),
.B2(n_366),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_379),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_304),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_389),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_351),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_320),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_387),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_384),
.A2(n_355),
.B1(n_366),
.B2(n_362),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_350),
.B(n_338),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_385),
.A2(n_328),
.B(n_297),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_263),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_326),
.Y(n_389)
);

NOR4xp25_ASAP7_75t_L g390 ( 
.A(n_346),
.B(n_326),
.C(n_329),
.D(n_310),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_390),
.B(n_336),
.CI(n_365),
.CON(n_395),
.SN(n_395)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_392),
.B(n_352),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_318),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_348),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_395),
.A2(n_396),
.B1(n_397),
.B2(n_398),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_308),
.B1(n_344),
.B2(n_355),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_380),
.Y(n_399)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_399),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_384),
.A2(n_366),
.B1(n_360),
.B2(n_328),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_409),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_411),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_403),
.C(n_408),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_358),
.C(n_354),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_372),
.B(n_339),
.Y(n_404)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_404),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_331),
.Y(n_405)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_405),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_353),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_414),
.Y(n_435)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_361),
.C(n_359),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_372),
.A2(n_295),
.B1(n_301),
.B2(n_343),
.Y(n_412)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_412),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_335),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_299),
.C(n_313),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_418),
.C(n_374),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_373),
.B(n_299),
.Y(n_417)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_417),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_380),
.C(n_385),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_413),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_431),
.B1(n_368),
.B2(n_386),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_426),
.B(n_433),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_377),
.Y(n_428)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_428),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_380),
.B1(n_394),
.B2(n_375),
.Y(n_429)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_429),
.Y(n_442)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_377),
.Y(n_432)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_416),
.C(n_415),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_SL g434 ( 
.A(n_418),
.B(n_394),
.C(n_333),
.Y(n_434)
);

FAx1_ASAP7_75t_SL g438 ( 
.A(n_434),
.B(n_426),
.CI(n_427),
.CON(n_438),
.SN(n_438)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_451),
.Y(n_465)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_427),
.A2(n_396),
.B(n_395),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_441),
.A2(n_409),
.B(n_430),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_416),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_445),
.Y(n_456)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_400),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_369),
.Y(n_446)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_411),
.C(n_386),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_450),
.B(n_452),
.Y(n_455)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_433),
.B(n_367),
.Y(n_452)
);

AOI22x1_ASAP7_75t_L g453 ( 
.A1(n_442),
.A2(n_436),
.B1(n_429),
.B2(n_421),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_454),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_435),
.C(n_434),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_464),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_437),
.B1(n_420),
.B2(n_409),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_461),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_424),
.C(n_386),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_424),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_449),
.C(n_450),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_467),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_441),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_448),
.C(n_442),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_472),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_465),
.B(n_444),
.Y(n_471)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_438),
.C(n_391),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_438),
.C(n_391),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_473),
.B(n_475),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_383),
.C(n_381),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_468),
.A2(n_459),
.B1(n_453),
.B2(n_457),
.Y(n_476)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_476),
.Y(n_485)
);

OAI321xp33_ASAP7_75t_L g478 ( 
.A1(n_471),
.A2(n_463),
.A3(n_453),
.B1(n_367),
.B2(n_383),
.C(n_381),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_478),
.A2(n_474),
.B(n_469),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_481),
.Y(n_482)
);

O2A1O1Ixp33_ASAP7_75t_L g487 ( 
.A1(n_482),
.A2(n_483),
.B(n_484),
.C(n_476),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_474),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_479),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_486),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_487),
.C(n_456),
.Y(n_489)
);

AOI322xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_456),
.A3(n_331),
.B1(n_464),
.B2(n_313),
.C1(n_280),
.C2(n_7),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_4),
.B(n_5),
.Y(n_491)
);

AOI21x1_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_4),
.B(n_5),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_7),
.Y(n_493)
);


endmodule