module fake_jpeg_187_n_232 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_232);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_10),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_22),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_35),
.B(n_17),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_85),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_95),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_70),
.B1(n_56),
.B2(n_79),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_98),
.B(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_58),
.B1(n_77),
.B2(n_74),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_58),
.B1(n_77),
.B2(n_56),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_88),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_R g129 ( 
.A(n_103),
.B(n_61),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_SL g105 ( 
.A(n_89),
.Y(n_105)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_120),
.Y(n_135)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_112),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_83),
.C(n_60),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_119),
.B1(n_111),
.B2(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_118),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_88),
.B1(n_87),
.B2(n_86),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_63),
.C(n_68),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_71),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_88),
.B1(n_87),
.B2(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_133),
.B1(n_80),
.B2(n_73),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_87),
.B1(n_79),
.B2(n_59),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_134),
.B1(n_4),
.B2(n_6),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_79),
.B1(n_80),
.B2(n_75),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_81),
.B1(n_90),
.B2(n_55),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_27),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_141),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_78),
.B1(n_65),
.B2(n_75),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_9),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_67),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_72),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_24),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_146),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_150),
.B1(n_159),
.B2(n_164),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_80),
.B(n_73),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_165),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_59),
.B1(n_62),
.B2(n_3),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_2),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_2),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_155),
.A2(n_163),
.B1(n_13),
.B2(n_14),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_7),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_168),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_23),
.C(n_50),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_167),
.C(n_32),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_11),
.Y(n_165)
);

HAxp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_12),
.CON(n_166),
.SN(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_26),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_12),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_171),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_33),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_20),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_140),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_176),
.C(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_177),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_128),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_166),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_128),
.B1(n_15),
.B2(n_16),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_183),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_186),
.B1(n_187),
.B2(n_19),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_37),
.B1(n_49),
.B2(n_47),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_198),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_21),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_199),
.B(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_183),
.B1(n_176),
.B2(n_181),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_38),
.C(n_25),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_169),
.C(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_211),
.C(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_189),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_202),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_187),
.C(n_180),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_208),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_193),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_207),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_212),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_221),
.B(n_223),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_218),
.A2(n_213),
.B(n_200),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_200),
.B1(n_191),
.B2(n_204),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_198),
.B(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_179),
.C(n_31),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_36),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_41),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_43),
.C(n_45),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_231),
.Y(n_232)
);


endmodule