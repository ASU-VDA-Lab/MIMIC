module fake_netlist_1_4998_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_L g13 ( .A(n_1), .B(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
AND2x2_ASAP7_75t_SL g15 ( .A(n_9), .B(n_1), .Y(n_15) );
OAI22xp5_ASAP7_75t_SL g16 ( .A1(n_6), .A2(n_2), .B1(n_10), .B2(n_11), .Y(n_16) );
OAI22xp5_ASAP7_75t_SL g17 ( .A1(n_2), .A2(n_0), .B1(n_5), .B2(n_12), .Y(n_17) );
O2A1O1Ixp5_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_3), .B(n_4), .C(n_5), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_14), .B(n_3), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_15), .B(n_17), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g21 ( .A(n_19), .B(n_14), .Y(n_21) );
OA21x2_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_19), .B(n_15), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_21), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_22), .Y(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_16), .B1(n_23), .B2(n_20), .C(n_8), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AO22x2_ASAP7_75t_SL g28 ( .A1(n_27), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_28) );
AOI21x1_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_27), .B(n_20), .Y(n_29) );
AOI221xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_8), .B1(n_9), .B2(n_10), .C(n_11), .Y(n_30) );
endmodule