module fake_netlist_1_12604_n_736 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_736);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_736;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_10), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_17), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_50), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_96), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_57), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_103), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_102), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_79), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_65), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_39), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_73), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_56), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_29), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_8), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_78), .Y(n_124) );
BUFx10_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
INVxp33_ASAP7_75t_SL g126 ( .A(n_45), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_13), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_71), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_62), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_108), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_59), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_93), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_47), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_7), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_6), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_53), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_7), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_64), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_43), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_21), .Y(n_145) );
INVx1_ASAP7_75t_SL g146 ( .A(n_54), .Y(n_146) );
BUFx5_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_5), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_34), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_26), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_0), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_66), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_21), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_145), .B(n_0), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_123), .B(n_1), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_111), .B(n_1), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g160 ( .A1(n_127), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_136), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_123), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_117), .B(n_22), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_136), .B(n_23), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_110), .B(n_2), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_125), .B(n_3), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_116), .Y(n_168) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_118), .B(n_24), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_125), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_119), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_120), .Y(n_172) );
BUFx12f_ASAP7_75t_L g173 ( .A(n_125), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_158), .A2(n_153), .B1(n_151), .B2(n_140), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_170), .B(n_148), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_170), .B(n_121), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_154), .Y(n_179) );
OR2x6_ASAP7_75t_L g180 ( .A(n_167), .B(n_124), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_161), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_170), .B(n_114), .Y(n_183) );
NAND2xp33_ASAP7_75t_L g184 ( .A(n_164), .B(n_147), .Y(n_184) );
XNOR2xp5_ASAP7_75t_L g185 ( .A(n_160), .B(n_127), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_170), .B(n_147), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_173), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_169), .B(n_128), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_161), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_156), .Y(n_191) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_164), .B(n_166), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_173), .B(n_166), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_173), .B(n_126), .Y(n_194) );
INVxp67_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_158), .A2(n_152), .B1(n_129), .B2(n_149), .Y(n_196) );
NAND3xp33_ASAP7_75t_L g197 ( .A(n_154), .B(n_135), .C(n_130), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_167), .Y(n_198) );
INVx4_ASAP7_75t_SL g199 ( .A(n_164), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_157), .B(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_198), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_186), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_200), .B(n_171), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_189), .A2(n_169), .B1(n_163), .B2(n_157), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_189), .A2(n_169), .B1(n_163), .B2(n_157), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_200), .B(n_171), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
NAND3xp33_ASAP7_75t_SL g208 ( .A(n_195), .B(n_112), .C(n_137), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_193), .B(n_159), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_189), .A2(n_158), .B1(n_154), .B2(n_164), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_179), .B(n_154), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_179), .B(n_158), .Y(n_212) );
INVxp33_ASAP7_75t_L g213 ( .A(n_187), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_177), .B(n_165), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_178), .B(n_165), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_180), .B(n_138), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_178), .B(n_162), .Y(n_217) );
OR2x6_ASAP7_75t_L g218 ( .A(n_180), .B(n_160), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_180), .A2(n_112), .B1(n_137), .B2(n_138), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_178), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_178), .B(n_162), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_186), .Y(n_222) );
OAI22xp5_ASAP7_75t_SL g223 ( .A1(n_185), .A2(n_142), .B1(n_109), .B2(n_139), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_192), .A2(n_156), .B(n_144), .Y(n_224) );
INVx5_ASAP7_75t_L g225 ( .A(n_175), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_180), .B(n_142), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_183), .B(n_131), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_180), .B(n_133), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_176), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_182), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_196), .B(n_115), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_194), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g233 ( .A1(n_185), .A2(n_134), .B1(n_146), .B2(n_122), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_174), .B(n_132), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_182), .Y(n_235) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_197), .B(n_164), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_213), .B(n_197), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_214), .B(n_188), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_212), .A2(n_184), .B(n_191), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_214), .B(n_188), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_207), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_219), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_201), .A2(n_191), .B(n_156), .C(n_181), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_215), .B(n_199), .Y(n_244) );
NOR2xp67_ASAP7_75t_L g245 ( .A(n_208), .B(n_4), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_204), .A2(n_168), .B1(n_172), .B2(n_141), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_212), .A2(n_181), .B(n_190), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
AO21x1_ASAP7_75t_L g249 ( .A1(n_236), .A2(n_181), .B(n_161), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_203), .B(n_199), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_229), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_205), .A2(n_168), .B1(n_172), .B2(n_143), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_235), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g255 ( .A(n_210), .B(n_25), .Y(n_255) );
OAI21x1_ASAP7_75t_SL g256 ( .A1(n_210), .A2(n_199), .B(n_164), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_220), .B(n_199), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_232), .B(n_150), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_225), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_202), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_209), .A2(n_227), .B(n_217), .C(n_222), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_209), .B(n_168), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_220), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_211), .A2(n_190), .B(n_175), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_227), .A2(n_172), .B(n_168), .C(n_161), .Y(n_265) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_224), .A2(n_164), .B(n_147), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_225), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_228), .A2(n_218), .B1(n_217), .B2(n_206), .Y(n_268) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_249), .A2(n_228), .A3(n_221), .B(n_231), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_250), .A2(n_234), .B(n_225), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_261), .A2(n_218), .B(n_216), .C(n_226), .Y(n_271) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_249), .A2(n_161), .A3(n_168), .B(n_172), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_255), .A2(n_168), .B(n_172), .C(n_225), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_238), .A2(n_190), .B(n_175), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_268), .A2(n_218), .B1(n_233), .B2(n_223), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_240), .Y(n_276) );
OAI222xp33_ASAP7_75t_L g277 ( .A1(n_242), .A2(n_5), .B1(n_6), .B2(n_8), .C1(n_9), .C2(n_10), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_264), .A2(n_164), .B(n_175), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_259), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_260), .B(n_172), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_241), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_242), .B(n_9), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g283 ( .A1(n_245), .A2(n_190), .B1(n_175), .B2(n_13), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_SL g285 ( .A1(n_265), .A2(n_60), .B(n_107), .C(n_106), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_255), .A2(n_190), .B(n_12), .C(n_14), .Y(n_286) );
AO31x2_ASAP7_75t_L g287 ( .A1(n_246), .A2(n_11), .A3(n_14), .B(n_15), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_259), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_260), .B(n_11), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_241), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_239), .A2(n_58), .B(n_104), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_263), .B(n_15), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_258), .B(n_16), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_276), .B(n_251), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_290), .Y(n_295) );
OAI322xp33_ASAP7_75t_L g296 ( .A1(n_275), .A2(n_237), .A3(n_262), .B1(n_252), .B2(n_251), .C1(n_253), .C2(n_254), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_271), .B(n_252), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_281), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_271), .B(n_263), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_281), .B(n_254), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_293), .B(n_248), .Y(n_301) );
AOI21x1_ASAP7_75t_L g302 ( .A1(n_274), .A2(n_256), .B(n_247), .Y(n_302) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_278), .A2(n_256), .B(n_248), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_288), .B(n_267), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_289), .B(n_267), .Y(n_305) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_273), .A2(n_244), .B(n_257), .Y(n_306) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_286), .A2(n_266), .B(n_243), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_270), .A2(n_266), .B(n_259), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_280), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_291), .A2(n_266), .B(n_259), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_280), .Y(n_311) );
OAI332xp33_ASAP7_75t_L g312 ( .A1(n_282), .A2(n_16), .A3(n_17), .B1(n_18), .B2(n_19), .B3(n_20), .C1(n_27), .C2(n_28), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_292), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_292), .B(n_18), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_303), .Y(n_316) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_308), .A2(n_297), .B(n_302), .Y(n_317) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_302), .A2(n_283), .B(n_285), .Y(n_318) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_307), .A2(n_283), .B(n_277), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_298), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_310), .A2(n_277), .B(n_269), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_303), .Y(n_322) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_307), .A2(n_269), .B(n_272), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_299), .B(n_269), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_298), .B(n_269), .Y(n_325) );
NOR2xp33_ASAP7_75t_R g326 ( .A(n_300), .B(n_279), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_298), .B(n_272), .Y(n_327) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_310), .A2(n_272), .B(n_287), .Y(n_328) );
OA21x2_ASAP7_75t_L g329 ( .A1(n_309), .A2(n_272), .B(n_287), .Y(n_329) );
OA21x2_ASAP7_75t_L g330 ( .A1(n_309), .A2(n_287), .B(n_279), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_315), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_315), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_287), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_315), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_300), .B(n_284), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_295), .B(n_19), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_312), .A2(n_20), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_315), .B(n_33), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_35), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_305), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_303), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_338), .A2(n_296), .B1(n_313), .B2(n_314), .Y(n_343) );
AO21x2_ASAP7_75t_L g344 ( .A1(n_318), .A2(n_307), .B(n_311), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_316), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_316), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_325), .B(n_307), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_316), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_320), .Y(n_353) );
INVx5_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_322), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_332), .B(n_315), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_332), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_338), .A2(n_296), .B1(n_294), .B2(n_301), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_332), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_341), .B(n_311), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_341), .B(n_301), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_341), .B(n_312), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_322), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_325), .B(n_305), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_334), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_325), .B(n_303), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_325), .B(n_304), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_338), .A2(n_306), .B1(n_315), .B2(n_38), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_326), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_319), .A2(n_306), .B1(n_37), .B2(n_40), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_324), .B(n_306), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_334), .B(n_306), .Y(n_380) );
INVx4_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_324), .B(n_105), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_334), .B(n_36), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_333), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_323), .B(n_101), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_333), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_324), .B(n_41), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_384), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_365), .B(n_323), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_365), .B(n_323), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_381), .B(n_323), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_375), .A2(n_337), .B(n_340), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_384), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_345), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_360), .B(n_329), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_367), .B(n_337), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_371), .B(n_323), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_372), .B(n_323), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_371), .B(n_329), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_386), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_372), .B(n_329), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_350), .B(n_329), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_349), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_350), .B(n_380), .Y(n_404) );
NOR3xp33_ASAP7_75t_SL g405 ( .A(n_368), .B(n_330), .C(n_319), .Y(n_405) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_354), .B(n_342), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_386), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_350), .B(n_329), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_380), .B(n_329), .Y(n_409) );
NAND2x1_ASAP7_75t_SL g410 ( .A(n_381), .B(n_337), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_381), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_360), .B(n_329), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_376), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_371), .B(n_330), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_380), .B(n_328), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_345), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_347), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_373), .B(n_328), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_374), .B(n_330), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_349), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_373), .B(n_328), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_361), .B(n_330), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_354), .B(n_337), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_346), .Y(n_426) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_367), .B(n_339), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_373), .B(n_328), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_361), .B(n_328), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_346), .Y(n_430) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_381), .B(n_342), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_363), .B(n_328), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_363), .B(n_330), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_353), .B(n_328), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_346), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_348), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_362), .B(n_330), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_362), .B(n_330), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_348), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_348), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_353), .B(n_321), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_377), .B(n_340), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_351), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_351), .Y(n_444) );
NOR2x1_ASAP7_75t_L g445 ( .A(n_377), .B(n_339), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_351), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_381), .B(n_332), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_374), .B(n_321), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_355), .B(n_321), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_355), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_347), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_366), .B(n_332), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_355), .B(n_369), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_369), .B(n_321), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_369), .B(n_321), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_388), .Y(n_456) );
BUFx2_ASAP7_75t_SL g457 ( .A(n_406), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_388), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_389), .B(n_379), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_404), .B(n_347), .Y(n_460) );
NAND2xp33_ASAP7_75t_L g461 ( .A(n_427), .B(n_354), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_404), .B(n_352), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_389), .B(n_379), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_394), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_409), .B(n_352), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_409), .B(n_352), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_405), .B(n_368), .C(n_375), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_393), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_390), .B(n_379), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_452), .B(n_357), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_427), .B(n_357), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_393), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_420), .B(n_374), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_400), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_400), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_394), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_397), .B(n_364), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_390), .B(n_344), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_420), .B(n_357), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_407), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_407), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_398), .B(n_344), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_453), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_414), .B(n_370), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_398), .B(n_344), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_402), .B(n_344), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_452), .Y(n_487) );
NOR2x1_ASAP7_75t_L g488 ( .A(n_445), .B(n_366), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_423), .B(n_383), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_402), .B(n_344), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_423), .B(n_383), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_428), .B(n_383), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_428), .B(n_359), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_415), .B(n_359), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_452), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_408), .B(n_370), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_414), .B(n_370), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_415), .B(n_359), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_408), .B(n_366), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_413), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_452), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_453), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_403), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_421), .B(n_366), .Y(n_504) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_394), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_413), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_418), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_401), .B(n_366), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_419), .Y(n_509) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_445), .B(n_339), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_421), .B(n_364), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_405), .B(n_378), .C(n_385), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_401), .B(n_321), .Y(n_513) );
AND2x4_ASAP7_75t_SL g514 ( .A(n_447), .B(n_356), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_422), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_451), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_392), .A2(n_343), .B(n_358), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_397), .B(n_385), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_399), .B(n_382), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_442), .B(n_387), .C(n_385), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_429), .B(n_321), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_399), .B(n_382), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_437), .B(n_382), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_436), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_416), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_437), .B(n_336), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_436), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_429), .B(n_432), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_438), .B(n_336), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_406), .B(n_447), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_432), .B(n_356), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_395), .B(n_319), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_440), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_451), .B(n_356), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_440), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_391), .B(n_356), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_391), .B(n_356), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_416), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_424), .Y(n_540) );
NOR2x1p5_ASAP7_75t_L g541 ( .A(n_531), .B(n_411), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_500), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_506), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_529), .B(n_431), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_484), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_509), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_473), .B(n_431), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_479), .B(n_431), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_516), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_456), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_507), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_468), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_517), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_438), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_510), .B(n_354), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_472), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_540), .B(n_395), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_518), .A2(n_343), .B1(n_358), .B2(n_411), .C(n_392), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_540), .B(n_412), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_493), .B(n_391), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_460), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_503), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_477), .B(n_434), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_531), .A2(n_410), .B(n_411), .C(n_418), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_474), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_486), .B(n_412), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_461), .A2(n_396), .B(n_447), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_475), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_504), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_480), .Y(n_572) );
OA21x2_ASAP7_75t_SL g573 ( .A1(n_501), .A2(n_391), .B(n_447), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_481), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_503), .Y(n_575) );
OAI32xp33_ASAP7_75t_L g576 ( .A1(n_521), .A2(n_411), .A3(n_425), .B1(n_418), .B2(n_424), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_515), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_494), .B(n_434), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_457), .B(n_410), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_477), .B(n_441), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_515), .B(n_448), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_461), .A2(n_433), .B(n_387), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_498), .B(n_441), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_486), .B(n_433), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_467), .A2(n_425), .A3(n_340), .B(n_448), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_464), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_496), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_490), .B(n_450), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_490), .B(n_450), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_525), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_488), .B(n_354), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_528), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_518), .A2(n_340), .B(n_378), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_534), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_459), .B(n_455), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_499), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g597 ( .A(n_512), .B(n_455), .C(n_454), .D(n_449), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_536), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_459), .B(n_454), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_464), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_463), .B(n_449), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_463), .B(n_446), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_462), .B(n_425), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_532), .B(n_446), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_465), .B(n_446), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_478), .B(n_430), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_466), .B(n_430), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_478), .A2(n_444), .B(n_443), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_482), .B(n_430), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_537), .B(n_444), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_476), .Y(n_611) );
OAI32xp33_ASAP7_75t_L g612 ( .A1(n_521), .A2(n_444), .A3(n_443), .B1(n_439), .B2(n_435), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_471), .A2(n_339), .B(n_354), .Y(n_613) );
AOI21xp33_ASAP7_75t_SL g614 ( .A1(n_471), .A2(n_339), .B(n_319), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_482), .B(n_439), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_SL g616 ( .A1(n_487), .A2(n_336), .B(n_439), .C(n_435), .Y(n_616) );
NOR2xp67_ASAP7_75t_SL g617 ( .A(n_520), .B(n_354), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_469), .B(n_443), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_485), .B(n_469), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_563), .B(n_487), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_564), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_578), .B(n_538), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_560), .A2(n_471), .B1(n_523), .B2(n_511), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_605), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_575), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_581), .B(n_485), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_555), .Y(n_627) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_559), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_577), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_541), .B(n_495), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_619), .B(n_519), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_542), .Y(n_632) );
AOI21xp33_ASAP7_75t_L g633 ( .A1(n_576), .A2(n_533), .B(n_319), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_543), .Y(n_634) );
OAI21xp33_ASAP7_75t_SL g635 ( .A1(n_573), .A2(n_489), .B(n_492), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_619), .B(n_491), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_568), .B(n_533), .Y(n_637) );
OA211x2_ASAP7_75t_L g638 ( .A1(n_585), .A2(n_513), .B(n_522), .C(n_514), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_546), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_597), .A2(n_495), .B1(n_508), .B2(n_470), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_566), .A2(n_513), .B(n_522), .C(n_535), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_549), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_562), .B(n_514), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_555), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_568), .B(n_483), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_590), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_592), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_594), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_556), .B(n_502), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_614), .B(n_470), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_593), .A2(n_524), .B1(n_530), .B2(n_527), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_553), .A2(n_505), .B1(n_319), .B2(n_476), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_612), .A2(n_505), .B(n_339), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_617), .B(n_354), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_584), .A2(n_539), .B1(n_526), .B2(n_435), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_587), .B(n_426), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_559), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_607), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_561), .B(n_426), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_561), .B(n_426), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_596), .B(n_417), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_598), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_550), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_552), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_584), .B(n_417), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_583), .B(n_417), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_554), .Y(n_667) );
AOI21xp33_ASAP7_75t_SL g668 ( .A1(n_579), .A2(n_416), .B(n_336), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_558), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_608), .A2(n_317), .B(n_335), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_623), .A2(n_627), .B(n_644), .C(n_635), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_623), .A2(n_548), .B1(n_565), .B2(n_544), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_641), .A2(n_603), .B1(n_557), .B2(n_569), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_638), .A2(n_580), .B1(n_547), .B2(n_571), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_650), .A2(n_668), .B1(n_579), .B2(n_654), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_628), .B(n_588), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_640), .A2(n_588), .B1(n_589), .B2(n_615), .Y(n_677) );
AO22x2_ASAP7_75t_L g678 ( .A1(n_621), .A2(n_613), .B1(n_591), .B2(n_567), .Y(n_678) );
OAI22xp33_ASAP7_75t_SL g679 ( .A1(n_620), .A2(n_579), .B1(n_557), .B2(n_589), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_651), .A2(n_609), .B1(n_615), .B2(n_606), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_632), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_657), .B(n_545), .Y(n_682) );
NOR2x1_ASAP7_75t_SL g683 ( .A(n_643), .B(n_618), .Y(n_683) );
OAI211xp5_ASAP7_75t_SL g684 ( .A1(n_633), .A2(n_593), .B(n_609), .C(n_606), .Y(n_684) );
AOI322xp5_ASAP7_75t_L g685 ( .A1(n_631), .A2(n_595), .A3(n_601), .B1(n_599), .B2(n_604), .C1(n_551), .C2(n_610), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_633), .A2(n_616), .B1(n_572), .B2(n_570), .C(n_574), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g687 ( .A1(n_653), .A2(n_582), .B(n_602), .C(n_600), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_634), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_639), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_630), .A2(n_611), .B(n_586), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_652), .A2(n_653), .B(n_637), .C(n_629), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_661), .Y(n_692) );
OAI322xp33_ASAP7_75t_SL g693 ( .A1(n_636), .A2(n_342), .A3(n_322), .B1(n_317), .B2(n_318), .C1(n_49), .C2(n_51), .Y(n_693) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_626), .A2(n_342), .A3(n_335), .B1(n_331), .B2(n_317), .C1(n_318), .C2(n_55), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_630), .A2(n_335), .B1(n_331), .B2(n_317), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_642), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g697 ( .A1(n_670), .A2(n_335), .B(n_331), .C(n_317), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_637), .B(n_317), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_671), .A2(n_670), .B(n_625), .C(n_667), .Y(n_699) );
AOI322xp5_ASAP7_75t_L g700 ( .A1(n_686), .A2(n_624), .A3(n_658), .B1(n_645), .B2(n_666), .C1(n_622), .C2(n_662), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_673), .A2(n_645), .B(n_659), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_684), .A2(n_669), .B1(n_648), .B2(n_664), .C(n_663), .Y(n_702) );
NOR2x1p5_ASAP7_75t_L g703 ( .A(n_676), .B(n_646), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_691), .A2(n_647), .B1(n_665), .B2(n_660), .C(n_656), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_681), .Y(n_705) );
AOI311xp33_ASAP7_75t_L g706 ( .A1(n_679), .A2(n_655), .A3(n_649), .B(n_654), .C(n_48), .Y(n_706) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_672), .A2(n_331), .B(n_318), .C(n_46), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_675), .A2(n_318), .B(n_44), .C(n_52), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g709 ( .A1(n_678), .A2(n_318), .B1(n_61), .B2(n_63), .C1(n_67), .C2(n_68), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_674), .A2(n_42), .B1(n_69), .B2(n_70), .Y(n_710) );
NOR2x1_ASAP7_75t_SL g711 ( .A(n_683), .B(n_72), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_677), .B(n_74), .Y(n_712) );
AOI222xp33_ASAP7_75t_L g713 ( .A1(n_678), .A2(n_75), .B1(n_76), .B2(n_77), .C1(n_80), .C2(n_81), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_706), .B(n_687), .C(n_694), .D(n_697), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_710), .A2(n_685), .B(n_690), .C(n_680), .Y(n_715) );
AOI211x1_ASAP7_75t_SL g716 ( .A1(n_699), .A2(n_695), .B(n_698), .C(n_693), .Y(n_716) );
OAI211xp5_ASAP7_75t_SL g717 ( .A1(n_700), .A2(n_689), .B(n_688), .C(n_696), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_702), .B(n_692), .Y(n_718) );
NOR3xp33_ASAP7_75t_L g719 ( .A(n_712), .B(n_682), .C(n_87), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_713), .B(n_85), .Y(n_720) );
AND2x4_ASAP7_75t_SL g721 ( .A(n_719), .B(n_705), .Y(n_721) );
XOR2xp5_ASAP7_75t_L g722 ( .A(n_716), .B(n_711), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_718), .Y(n_723) );
NOR3xp33_ASAP7_75t_SL g724 ( .A(n_720), .B(n_714), .C(n_717), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_723), .A2(n_715), .B1(n_701), .B2(n_703), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_724), .B(n_704), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_722), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_727), .B(n_721), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_726), .A2(n_709), .B1(n_708), .B2(n_707), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_728), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_729), .Y(n_731) );
OAI21x1_ASAP7_75t_L g732 ( .A1(n_730), .A2(n_725), .B(n_707), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_731), .B(n_89), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_733), .A2(n_90), .B1(n_92), .B2(n_95), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_734), .Y(n_735) );
AOI222xp33_ASAP7_75t_L g736 ( .A1(n_735), .A2(n_732), .B1(n_98), .B2(n_99), .C1(n_100), .C2(n_97), .Y(n_736) );
endmodule