module fake_jpeg_29350_n_391 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_391);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_391;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx2_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_48),
.Y(n_90)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_17),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_67),
.Y(n_93)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_12),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx2_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_63),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_12),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_66),
.Y(n_108)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_21),
.B(n_11),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_76),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_37),
.B(n_0),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_22),
.B(n_33),
.C(n_32),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_11),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_80),
.Y(n_127)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_11),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_81),
.B(n_1),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_16),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_88),
.A2(n_100),
.B1(n_105),
.B2(n_111),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_96),
.B(n_134),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_29),
.B1(n_38),
.B2(n_34),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_98),
.A2(n_102),
.B1(n_123),
.B2(n_132),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_46),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_29),
.B1(n_38),
.B2(n_34),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_40),
.B1(n_35),
.B2(n_28),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_16),
.B1(n_20),
.B2(n_85),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_69),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_20),
.B1(n_22),
.B2(n_33),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_49),
.A2(n_32),
.B(n_26),
.C(n_40),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_82),
.B(n_80),
.C(n_48),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_59),
.A2(n_35),
.B1(n_28),
.B2(n_23),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_119),
.A2(n_128),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_28),
.B1(n_23),
.B2(n_2),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_45),
.A2(n_58),
.B1(n_82),
.B2(n_65),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_77),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_56),
.A2(n_79),
.B1(n_51),
.B2(n_68),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_52),
.A2(n_28),
.B1(n_23),
.B2(n_4),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_82),
.B1(n_62),
.B2(n_60),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_80),
.Y(n_147)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_57),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_84),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_93),
.B(n_83),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_146),
.B(n_165),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_169),
.B1(n_100),
.B2(n_119),
.Y(n_195)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_94),
.B(n_50),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_156),
.Y(n_205)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_161),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_113),
.B(n_64),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_160),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_86),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_114),
.B(n_1),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_170),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_96),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_90),
.B(n_116),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_135),
.B1(n_99),
.B2(n_97),
.Y(n_197)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_6),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_172),
.B(n_105),
.Y(n_214)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_6),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_176),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_7),
.C(n_8),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_182),
.Y(n_210)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_95),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_139),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_88),
.B(n_7),
.Y(n_180)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

CKINVDCx10_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_188),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_203),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_131),
.B1(n_138),
.B2(n_92),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_201),
.B1(n_208),
.B2(n_99),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_195),
.A2(n_217),
.B1(n_208),
.B2(n_151),
.Y(n_245)
);

OAI22x1_ASAP7_75t_L g246 ( 
.A1(n_197),
.A2(n_124),
.B1(n_140),
.B2(n_165),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_138),
.B1(n_91),
.B2(n_92),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_207),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

AO21x2_ASAP7_75t_L g208 ( 
.A1(n_146),
.A2(n_128),
.B(n_124),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_211),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_143),
.B(n_118),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_142),
.B(n_103),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_103),
.B1(n_106),
.B2(n_115),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_222),
.A2(n_246),
.B1(n_247),
.B2(n_251),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_174),
.B1(n_157),
.B2(n_106),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_174),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_241),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_195),
.B1(n_189),
.B2(n_208),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_250),
.B(n_208),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_216),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_237),
.B(n_242),
.Y(n_271)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_180),
.C(n_168),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_187),
.C(n_186),
.Y(n_264)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_243),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_163),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_244),
.B(n_248),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_208),
.B1(n_187),
.B2(n_214),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_203),
.A2(n_177),
.B1(n_172),
.B2(n_115),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_153),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_206),
.B(n_209),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_164),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_173),
.B1(n_176),
.B2(n_167),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_199),
.B(n_182),
.CI(n_178),
.CON(n_252),
.SN(n_252)
);

OA21x2_ASAP7_75t_SL g265 ( 
.A1(n_252),
.A2(n_187),
.B(n_208),
.Y(n_265)
);

AOI32xp33_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_97),
.A3(n_121),
.B1(n_107),
.B2(n_150),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_211),
.B(n_209),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_263),
.C(n_264),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_257),
.A2(n_191),
.B1(n_198),
.B2(n_221),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_276),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_186),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_265),
.B(n_267),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_226),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_266),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_233),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_251),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_223),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_277),
.C(n_228),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_210),
.B(n_205),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_223),
.B(n_217),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_278),
.B(n_279),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_246),
.B1(n_238),
.B2(n_253),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_281),
.A2(n_286),
.B1(n_289),
.B2(n_277),
.Y(n_324)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_245),
.B1(n_231),
.B2(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_234),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_296),
.C(n_294),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_288),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_222),
.B1(n_235),
.B2(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_266),
.B(n_252),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_256),
.A2(n_247),
.B1(n_252),
.B2(n_225),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_196),
.B1(n_243),
.B2(n_192),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_261),
.B1(n_192),
.B2(n_243),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_293),
.B(n_294),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_232),
.B1(n_242),
.B2(n_241),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_239),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_270),
.B1(n_275),
.B2(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_307),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_257),
.B1(n_279),
.B2(n_278),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_308),
.A2(n_324),
.B1(n_313),
.B2(n_312),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_309),
.A2(n_316),
.B(n_319),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_264),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_287),
.C(n_296),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_262),
.B(n_267),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_271),
.Y(n_318)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_299),
.A2(n_304),
.B1(n_292),
.B2(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_280),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_290),
.A2(n_262),
.B(n_271),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_288),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_275),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_326),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_314),
.B1(n_305),
.B2(n_269),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_333),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_287),
.C(n_290),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_336),
.C(n_341),
.Y(n_345)
);

AOI322xp5_ASAP7_75t_SL g330 ( 
.A1(n_320),
.A2(n_303),
.A3(n_289),
.B1(n_280),
.B2(n_272),
.C1(n_293),
.C2(n_274),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_330),
.B(n_315),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_318),
.A2(n_306),
.B(n_316),
.Y(n_332)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_332),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_322),
.C(n_311),
.Y(n_336)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_337),
.Y(n_350)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_302),
.B1(n_301),
.B2(n_300),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_314),
.B(n_305),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_321),
.B(n_308),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_298),
.C(n_191),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_202),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_339),
.A2(n_324),
.B1(n_323),
.B2(n_315),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_343),
.A2(n_339),
.B1(n_327),
.B2(n_340),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_348),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_354),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_269),
.B1(n_198),
.B2(n_196),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_352),
.B(n_353),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_230),
.C(n_221),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_335),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_331),
.A2(n_196),
.B1(n_149),
.B2(n_202),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_190),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_334),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_359),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_350),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_338),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_360),
.B(n_364),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_363),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_346),
.A2(n_329),
.B(n_341),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_362),
.A2(n_166),
.B(n_126),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_349),
.A2(n_336),
.B1(n_333),
.B2(n_107),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_141),
.B1(n_166),
.B2(n_179),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_366),
.A2(n_345),
.B(n_353),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_370),
.A2(n_373),
.B(n_376),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_364),
.A2(n_347),
.B1(n_355),
.B2(n_345),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_372),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_358),
.B(n_351),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_351),
.C(n_218),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_373),
.A2(n_375),
.B(n_367),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_365),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_357),
.Y(n_380)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

AOI21x1_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_382),
.B(n_374),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_121),
.C(n_190),
.Y(n_382)
);

AOI21x1_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_368),
.B(n_190),
.Y(n_388)
);

NOR3xp33_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_379),
.C(n_380),
.Y(n_387)
);

OAI321xp33_ASAP7_75t_L g389 ( 
.A1(n_387),
.A2(n_388),
.A3(n_385),
.B1(n_383),
.B2(n_368),
.C(n_181),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_120),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_9),
.Y(n_391)
);


endmodule