module fake_netlist_5_829_n_2305 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2305);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2305;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_339;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_2248;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2213;
wire n_2023;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_138),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_157),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_75),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_67),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_87),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_154),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_201),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_112),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_175),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_62),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_78),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_41),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_105),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_142),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_38),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_152),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_27),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_184),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_6),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_203),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_168),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_34),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_43),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_177),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_136),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_183),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_12),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_106),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_72),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_26),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_187),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_44),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_146),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_119),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_206),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_76),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_81),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_46),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_71),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_20),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_179),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_9),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_160),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_111),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_95),
.Y(n_281)
);

BUFx8_ASAP7_75t_SL g282 ( 
.A(n_204),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_18),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_75),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_82),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_135),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_9),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_63),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_97),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_41),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_208),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_64),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_10),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_23),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_107),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_47),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_166),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_214),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_14),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_192),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_61),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_42),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_86),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_37),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_131),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_84),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_176),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_4),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_82),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_210),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_19),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_86),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_76),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_158),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_79),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_66),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_81),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_212),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_0),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_98),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_62),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_25),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_182),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_7),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_31),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_218),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_39),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_22),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_178),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_172),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_150),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_84),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_115),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_34),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_16),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_10),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_61),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_90),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_68),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_53),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_200),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_73),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_100),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_110),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_173),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_54),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_170),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_51),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_38),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_79),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_85),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_19),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_20),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_193),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_197),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_104),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_7),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_14),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_148),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_89),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_188),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_42),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_69),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_128),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_171),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_58),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_72),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_102),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_33),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_147),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_50),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_83),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_120),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_5),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_27),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_40),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_35),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_73),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_216),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_39),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_0),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_199),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_33),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_66),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_69),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_181),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_67),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_85),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_63),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_185),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_202),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_125),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_167),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_22),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_215),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_12),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_134),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_162),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_17),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_96),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_217),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_117),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_15),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_23),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_169),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_198),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_92),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_141),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_165),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_94),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_24),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_56),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_196),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_59),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_123),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_77),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_74),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_47),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_140),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_43),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_114),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_51),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_57),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_55),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_116),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_70),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_149),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_70),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_262),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_262),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_308),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_282),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_262),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_398),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_316),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_250),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_250),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_219),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_220),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_225),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_262),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_262),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_262),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_229),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_231),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_262),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_234),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_223),
.B(n_1),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_255),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_262),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_223),
.B(n_1),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_242),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_262),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_319),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_244),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_245),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_319),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_319),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_319),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_253),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_319),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_319),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_2),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_257),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_261),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_330),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_268),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_276),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_316),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_410),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_330),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_330),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_330),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_330),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_347),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_255),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_278),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_330),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_280),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_287),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_291),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_292),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_331),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_331),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_331),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_300),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_301),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_303),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_401),
.B(n_2),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_228),
.B(n_3),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_310),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_390),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_313),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_351),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_351),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_256),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_317),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_312),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_256),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_321),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_323),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_326),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_329),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_256),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_333),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_344),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_285),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_285),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_224),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_241),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_357),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_224),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_285),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_227),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_232),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_358),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_359),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_367),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_368),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_241),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_373),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_221),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_376),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_232),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_239),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_239),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_228),
.B(n_3),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_222),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_235),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_241),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_243),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_382),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_243),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_237),
.B(n_4),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_385),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_273),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_443),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_502),
.B(n_227),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_531),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_237),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_433),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_R g552 ( 
.A(n_435),
.B(n_400),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_457),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_502),
.B(n_505),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_447),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_444),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_448),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

INVxp33_ASAP7_75t_L g561 ( 
.A(n_537),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_460),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_538),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_504),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_450),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_461),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_520),
.B(n_422),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_461),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_505),
.B(n_227),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_462),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_459),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_464),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_451),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_463),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_468),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_464),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_465),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_465),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_469),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_469),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_439),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_510),
.B(n_334),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_475),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_438),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_470),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_475),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_482),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_520),
.B(n_422),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_510),
.B(n_334),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_432),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_476),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_513),
.B(n_334),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_R g599 ( 
.A(n_454),
.B(n_431),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_434),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_436),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_495),
.B(n_403),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_436),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_R g604 ( 
.A(n_483),
.B(n_404),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_445),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_445),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_477),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_481),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_536),
.B(n_543),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_481),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_513),
.B(n_408),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_514),
.B(n_281),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_533),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_446),
.B(n_449),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_440),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_484),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_485),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_533),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_472),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_437),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_534),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_446),
.Y(n_624)
);

BUFx8_ASAP7_75t_L g625 ( 
.A(n_514),
.Y(n_625)
);

BUFx8_ASAP7_75t_L g626 ( 
.A(n_519),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_489),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_535),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_441),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_442),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_540),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_497),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_499),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_506),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_555),
.B(n_519),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_551),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_610),
.B(n_507),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_603),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_551),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_600),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_610),
.B(n_508),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_615),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g644 ( 
.A(n_569),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_576),
.A2(n_494),
.B1(n_466),
.B2(n_478),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_602),
.B(n_509),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_603),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_576),
.B(n_511),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_615),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_555),
.B(n_548),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_569),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_602),
.B(n_512),
.Y(n_652)
);

CKINVDCx8_ASAP7_75t_R g653 ( 
.A(n_547),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_615),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_551),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_552),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_615),
.A2(n_548),
.B1(n_587),
.B2(n_571),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_603),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_615),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_560),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_560),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_549),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_589),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_555),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_604),
.B(n_517),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_551),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_560),
.B(n_281),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_548),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_589),
.B(n_452),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_551),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_571),
.A2(n_493),
.B1(n_290),
.B2(n_299),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_604),
.B(n_526),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_561),
.B(n_527),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_546),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_612),
.B(n_530),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_556),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_612),
.B(n_544),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_552),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_551),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_560),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_559),
.B(n_516),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_635),
.B(n_529),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_565),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_571),
.B(n_587),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_596),
.B(n_281),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_596),
.B(n_362),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_613),
.B(n_226),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_596),
.Y(n_689)
);

AND2x2_ASAP7_75t_SL g690 ( 
.A(n_550),
.B(n_362),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_587),
.B(n_522),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_566),
.B(n_455),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_573),
.B(n_539),
.Y(n_694)
);

XOR2xp5_ASAP7_75t_L g695 ( 
.A(n_622),
.B(n_630),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_596),
.B(n_428),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_596),
.B(n_449),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_601),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_601),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_603),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_577),
.B(n_479),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_546),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_601),
.B(n_453),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_546),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_578),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_590),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_557),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_601),
.B(n_453),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_593),
.B(n_458),
.Y(n_709)
);

BUFx4_ASAP7_75t_L g710 ( 
.A(n_631),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_617),
.B(n_467),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_595),
.B(n_522),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_595),
.B(n_525),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_558),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_599),
.A2(n_318),
.B1(n_391),
.B2(n_233),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_601),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_558),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_618),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_595),
.B(n_525),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_558),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_627),
.B(n_471),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_598),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_633),
.B(n_273),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_634),
.B(n_480),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_598),
.B(n_528),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_598),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_557),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_624),
.B(n_456),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_613),
.B(n_614),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_624),
.Y(n_731)
);

BUFx4f_ASAP7_75t_L g732 ( 
.A(n_603),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_557),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_563),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_549),
.B(n_490),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_624),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_558),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_624),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_620),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_586),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_624),
.B(n_456),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_558),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_603),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_613),
.B(n_528),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_564),
.B(n_492),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_563),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_SL g748 ( 
.A1(n_564),
.A2(n_293),
.B1(n_341),
.B2(n_288),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_565),
.B(n_503),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_553),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_620),
.B(n_523),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_550),
.B(n_240),
.Y(n_752)
);

OAI21xp33_ASAP7_75t_SL g753 ( 
.A1(n_568),
.A2(n_594),
.B(n_275),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_568),
.A2(n_487),
.B(n_486),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_594),
.B(n_332),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_553),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_614),
.B(n_226),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_619),
.B(n_621),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_599),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_603),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_606),
.B(n_230),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_619),
.B(n_621),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_623),
.B(n_230),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_606),
.B(n_405),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_586),
.B(n_515),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_570),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_554),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_606),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_623),
.B(n_524),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_558),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_554),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_606),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_570),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_606),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_562),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_625),
.A2(n_290),
.B1(n_299),
.B2(n_277),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_562),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_606),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_567),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_616),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_567),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_572),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_570),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_616),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_606),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_628),
.B(n_486),
.Y(n_786)
);

BUFx4f_ASAP7_75t_L g787 ( 
.A(n_607),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_588),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_572),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_607),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_638),
.B(n_642),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_648),
.B(n_532),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_643),
.Y(n_793)
);

NAND2x1p5_ASAP7_75t_L g794 ( 
.A(n_659),
.B(n_236),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_657),
.B(n_685),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_659),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_685),
.B(n_646),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_750),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_643),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_652),
.B(n_541),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_649),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_759),
.B(n_625),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_669),
.B(n_607),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_669),
.B(n_607),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_759),
.A2(n_626),
.B1(n_625),
.B2(n_411),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_722),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_784),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_SL g808 ( 
.A(n_748),
.B(n_423),
.C(n_415),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_676),
.B(n_625),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_750),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_678),
.B(n_625),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_651),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_739),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_649),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_756),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_722),
.A2(n_428),
.B1(n_238),
.B2(n_247),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_654),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_726),
.B(n_607),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_656),
.B(n_626),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_674),
.B(n_626),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_690),
.A2(n_626),
.B1(n_238),
.B2(n_247),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_706),
.Y(n_822)
);

AND2x4_ASAP7_75t_SL g823 ( 
.A(n_705),
.B(n_336),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_726),
.B(n_607),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_656),
.B(n_626),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_740),
.B(n_644),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_654),
.A2(n_249),
.B(n_251),
.C(n_236),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_729),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_650),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_769),
.B(n_246),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_650),
.Y(n_831)
);

OR2x6_ASAP7_75t_SL g832 ( 
.A(n_780),
.B(n_248),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_690),
.B(n_607),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_692),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_690),
.A2(n_249),
.B1(n_252),
.B2(n_251),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_692),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_729),
.A2(n_416),
.B1(n_424),
.B2(n_409),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_729),
.B(n_574),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_712),
.B(n_628),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_729),
.A2(n_645),
.B1(n_713),
.B2(n_712),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_756),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_765),
.B(n_258),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_752),
.B(n_574),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_755),
.B(n_575),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_765),
.B(n_259),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_665),
.B(n_575),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_751),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_679),
.B(n_336),
.Y(n_848)
);

INVx8_ASAP7_75t_L g849 ( 
.A(n_677),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_679),
.B(n_336),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_754),
.A2(n_580),
.B(n_579),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_684),
.B(n_263),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_665),
.B(n_579),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_767),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_776),
.A2(n_252),
.B1(n_260),
.B2(n_254),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_670),
.B(n_518),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_713),
.B(n_629),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_688),
.A2(n_254),
.B1(n_264),
.B2(n_260),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_684),
.B(n_266),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_688),
.A2(n_264),
.B1(n_267),
.B2(n_265),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_758),
.B(n_580),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_767),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_771),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_677),
.Y(n_864)
);

AND2x2_ASAP7_75t_SL g865 ( 
.A(n_688),
.B(n_265),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_715),
.B(n_336),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_SL g867 ( 
.A1(n_746),
.A2(n_780),
.B1(n_718),
.B2(n_706),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_758),
.B(n_581),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_651),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_758),
.B(n_581),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_771),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_739),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_775),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_775),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_777),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_719),
.A2(n_267),
.B1(n_279),
.B2(n_269),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_758),
.B(n_582),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_762),
.B(n_582),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_762),
.B(n_583),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_777),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_668),
.B(n_269),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_688),
.A2(n_286),
.B1(n_294),
.B2(n_279),
.Y(n_882)
);

AOI22x1_ASAP7_75t_L g883 ( 
.A1(n_660),
.A2(n_286),
.B1(n_298),
.B2(n_294),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_663),
.B(n_350),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_762),
.B(n_583),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_762),
.B(n_745),
.Y(n_886)
);

O2A1O1Ixp5_ASAP7_75t_L g887 ( 
.A1(n_660),
.A2(n_662),
.B(n_681),
.C(n_661),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_745),
.A2(n_430),
.B1(n_298),
.B2(n_394),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_663),
.B(n_719),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_653),
.B(n_350),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_725),
.A2(n_389),
.B1(n_346),
.B2(n_348),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_670),
.B(n_270),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_664),
.B(n_271),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_725),
.B(n_584),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_666),
.B(n_272),
.Y(n_895)
);

AND2x6_ASAP7_75t_SL g896 ( 
.A(n_693),
.B(n_274),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_779),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_673),
.B(n_350),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_784),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_779),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_636),
.B(n_584),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_636),
.B(n_629),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_781),
.B(n_585),
.Y(n_903)
);

O2A1O1Ixp5_ASAP7_75t_L g904 ( 
.A1(n_661),
.A2(n_585),
.B(n_611),
.C(n_592),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_757),
.A2(n_346),
.B1(n_394),
.B2(n_395),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_781),
.B(n_592),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_782),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_749),
.B(n_701),
.Y(n_908)
);

AND2x4_ASAP7_75t_SL g909 ( 
.A(n_705),
.B(n_350),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_782),
.B(n_597),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_757),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_739),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_789),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_753),
.B(n_705),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_754),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_789),
.B(n_597),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_662),
.B(n_605),
.Y(n_917)
);

BUFx5_ASAP7_75t_L g918 ( 
.A(n_668),
.Y(n_918)
);

OAI22xp33_ASAP7_75t_L g919 ( 
.A1(n_764),
.A2(n_364),
.B1(n_430),
.B2(n_396),
.Y(n_919)
);

AND2x6_ASAP7_75t_SL g920 ( 
.A(n_709),
.B(n_274),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_675),
.Y(n_921)
);

NOR3xp33_ASAP7_75t_L g922 ( 
.A(n_735),
.B(n_378),
.C(n_314),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_681),
.B(n_605),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_689),
.B(n_611),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_689),
.B(n_348),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_741),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_723),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_677),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_698),
.B(n_364),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_682),
.B(n_521),
.C(n_277),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_757),
.B(n_632),
.Y(n_931)
);

INVxp33_ASAP7_75t_L g932 ( 
.A(n_695),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_698),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_699),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_699),
.B(n_371),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_723),
.A2(n_396),
.B1(n_418),
.B2(n_413),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_757),
.B(n_632),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_668),
.B(n_686),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_716),
.B(n_371),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_716),
.B(n_389),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_731),
.B(n_393),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_763),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_683),
.B(n_283),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_753),
.B(n_393),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_731),
.B(n_736),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_736),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_763),
.B(n_395),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_705),
.B(n_412),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_763),
.B(n_412),
.Y(n_949)
);

AND2x6_ASAP7_75t_SL g950 ( 
.A(n_710),
.B(n_275),
.Y(n_950)
);

NAND2x1p5_ASAP7_75t_L g951 ( 
.A(n_744),
.B(n_413),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_732),
.A2(n_591),
.B(n_588),
.Y(n_952)
);

INVxp67_ASAP7_75t_SL g953 ( 
.A(n_637),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_675),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_763),
.B(n_418),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_668),
.A2(n_609),
.B1(n_608),
.B2(n_591),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_786),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_653),
.B(n_289),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_640),
.B(n_671),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_668),
.B(n_296),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_677),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_694),
.B(n_711),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_640),
.B(n_588),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_828),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_828),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_822),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_791),
.B(n_718),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_793),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_849),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_822),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_793),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_847),
.B(n_721),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_799),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_798),
.Y(n_974)
);

AND2x6_ASAP7_75t_SL g975 ( 
.A(n_792),
.B(n_284),
.Y(n_975)
);

BUFx10_ASAP7_75t_L g976 ( 
.A(n_820),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_799),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_801),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_926),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_798),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_797),
.B(n_640),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_812),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_856),
.B(n_724),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_829),
.B(n_831),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_795),
.A2(n_686),
.B1(n_668),
.B2(n_687),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_801),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_814),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_912),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_813),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_814),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_817),
.Y(n_991)
);

BUFx12f_ASAP7_75t_L g992 ( 
.A(n_807),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_817),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_849),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_806),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_856),
.B(n_695),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_796),
.B(n_786),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_865),
.B(n_640),
.Y(n_998)
);

INVx4_ASAP7_75t_L g999 ( 
.A(n_849),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_829),
.A2(n_668),
.B1(n_686),
.B2(n_687),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_SL g1001 ( 
.A(n_864),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_810),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_933),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_933),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_934),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_869),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_831),
.B(n_697),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_796),
.B(n_641),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_834),
.B(n_703),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_810),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_815),
.Y(n_1011)
);

NOR2xp67_ASAP7_75t_L g1012 ( 
.A(n_899),
.B(n_672),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_865),
.B(n_671),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_957),
.B(n_834),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_934),
.Y(n_1015)
);

NOR2x1p5_ASAP7_75t_L g1016 ( 
.A(n_808),
.B(n_710),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_806),
.B(n_760),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_912),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_815),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_813),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_918),
.B(n_671),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_902),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_946),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_836),
.B(n_708),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_864),
.B(n_744),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_836),
.B(n_728),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_928),
.B(n_744),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_946),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_912),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_800),
.B(n_677),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_813),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_931),
.B(n_760),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_872),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_871),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_928),
.B(n_774),
.Y(n_1035)
);

BUFx8_ASAP7_75t_L g1036 ( 
.A(n_961),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_872),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_931),
.B(n_768),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_871),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_830),
.A2(n_686),
.B1(n_696),
.B2(n_687),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_872),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_937),
.B(n_768),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_L g1043 ( 
.A(n_961),
.B(n_742),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_SL g1044 ( 
.A(n_890),
.B(n_241),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_807),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_912),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_826),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_875),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_875),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_880),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_880),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_912),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_902),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_843),
.B(n_671),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_844),
.B(n_691),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_849),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_842),
.B(n_658),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_915),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_803),
.A2(n_787),
.B(n_732),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_807),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_841),
.B(n_691),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_897),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_897),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_918),
.B(n_691),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_841),
.B(n_691),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_900),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_937),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_867),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_854),
.B(n_714),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_957),
.B(n_702),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_854),
.B(n_714),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_862),
.B(n_714),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_839),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_950),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_900),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_862),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_927),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_863),
.B(n_714),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_911),
.B(n_738),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_915),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_942),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_839),
.Y(n_1083)
);

BUFx4f_ASAP7_75t_SL g1084 ( 
.A(n_958),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_896),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_863),
.Y(n_1086)
);

AND3x1_ASAP7_75t_SL g1087 ( 
.A(n_920),
.B(n_295),
.C(n_284),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_886),
.B(n_761),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_942),
.B(n_738),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_918),
.B(n_738),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_873),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_873),
.B(n_738),
.Y(n_1092)
);

INVx5_ASAP7_75t_L g1093 ( 
.A(n_915),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_918),
.B(n_743),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_857),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_921),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_852),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_921),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_889),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_954),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_918),
.B(n_743),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_857),
.B(n_743),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_874),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_845),
.B(n_658),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_874),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_794),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_954),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_823),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_907),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_840),
.A2(n_304),
.B(n_295),
.C(n_325),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_907),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_794),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_913),
.B(n_743),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_913),
.Y(n_1114)
);

AND2x2_ASAP7_75t_SL g1115 ( 
.A(n_821),
.B(n_304),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_859),
.B(n_702),
.Y(n_1116)
);

OAI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_901),
.A2(n_761),
.B1(n_366),
.B2(n_429),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_794),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_832),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_851),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_851),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_894),
.B(n_835),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_951),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_846),
.B(n_790),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_945),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_838),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_892),
.B(n_704),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_918),
.B(n_774),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_861),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_832),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_914),
.B(n_658),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_853),
.B(n_790),
.Y(n_1132)
);

BUFx4f_ASAP7_75t_L g1133 ( 
.A(n_951),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_951),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_868),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_870),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_804),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_877),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_878),
.B(n_879),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_885),
.B(n_790),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_809),
.B(n_774),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_887),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_904),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_811),
.B(n_774),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_818),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_944),
.B(n_819),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_903),
.B(n_785),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_932),
.B(n_540),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_960),
.B(n_785),
.Y(n_1149)
);

AO21x2_ASAP7_75t_L g1150 ( 
.A1(n_833),
.A2(n_737),
.B(n_734),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_906),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_910),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_858),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_918),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_824),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_893),
.B(n_704),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_916),
.B(n_785),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1122),
.A2(n_1030),
.B1(n_1125),
.B2(n_1126),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1151),
.B(n_895),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1131),
.A2(n_959),
.B(n_963),
.Y(n_1160)
);

AO21x1_ASAP7_75t_L g1161 ( 
.A1(n_998),
.A2(n_929),
.B(n_925),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1074),
.A2(n_962),
.B1(n_908),
.B2(n_837),
.Y(n_1162)
);

OR2x4_ASAP7_75t_L g1163 ( 
.A(n_996),
.B(n_943),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_988),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1058),
.A2(n_787),
.B(n_732),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1059),
.A2(n_923),
.B(n_917),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1058),
.A2(n_787),
.B(n_938),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1152),
.B(n_860),
.Y(n_1168)
);

AOI31xp67_ASAP7_75t_L g1169 ( 
.A1(n_1143),
.A2(n_939),
.A3(n_940),
.B(n_935),
.Y(n_1169)
);

AOI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1097),
.A2(n_866),
.B(n_932),
.Y(n_1170)
);

AOI211x1_ASAP7_75t_L g1171 ( 
.A1(n_984),
.A2(n_882),
.B(n_855),
.C(n_816),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1111),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1058),
.A2(n_938),
.B(n_953),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1058),
.A2(n_700),
.B(n_658),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_967),
.A2(n_972),
.B1(n_1146),
.B2(n_983),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1022),
.B(n_891),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_L g1177 ( 
.A(n_979),
.B(n_966),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1061),
.A2(n_924),
.B(n_941),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1111),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_979),
.Y(n_1180)
);

AO21x1_ASAP7_75t_L g1181 ( 
.A1(n_998),
.A2(n_1013),
.B(n_1057),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1074),
.A2(n_888),
.B1(n_905),
.B2(n_802),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_982),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1131),
.A2(n_949),
.B(n_947),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1022),
.B(n_1053),
.Y(n_1185)
);

NOR2xp67_ASAP7_75t_L g1186 ( 
.A(n_966),
.B(n_948),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1053),
.B(n_955),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1045),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1142),
.A2(n_1143),
.B(n_1121),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1058),
.A2(n_772),
.B(n_700),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1110),
.A2(n_827),
.A3(n_952),
.B(n_737),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1110),
.A2(n_936),
.B(n_876),
.C(n_909),
.Y(n_1192)
);

OA22x2_ASAP7_75t_L g1193 ( 
.A1(n_1068),
.A2(n_823),
.B1(n_909),
.B2(n_884),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1114),
.Y(n_1194)
);

AO21x2_ASAP7_75t_L g1195 ( 
.A1(n_1141),
.A2(n_825),
.B(n_898),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1095),
.B(n_848),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1142),
.A2(n_790),
.B(n_785),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1095),
.B(n_1014),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_970),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1120),
.A2(n_883),
.B(n_761),
.Y(n_1200)
);

OAI21xp33_ASAP7_75t_L g1201 ( 
.A1(n_1044),
.A2(n_922),
.B(n_850),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1014),
.B(n_930),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1071),
.B(n_918),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1065),
.A2(n_883),
.B(n_956),
.Y(n_1204)
);

NAND2xp33_ASAP7_75t_L g1205 ( 
.A(n_1056),
.B(n_686),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1069),
.A2(n_727),
.B(n_707),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1120),
.A2(n_788),
.A3(n_747),
.B(n_773),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1129),
.B(n_919),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1135),
.B(n_707),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1081),
.A2(n_772),
.B(n_700),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_981),
.A2(n_1121),
.B(n_1073),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1114),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1072),
.A2(n_733),
.B(n_727),
.Y(n_1213)
);

BUFx2_ASAP7_75t_SL g1214 ( 
.A(n_1001),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_981),
.A2(n_733),
.B(n_734),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1006),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1083),
.A2(n_805),
.B1(n_655),
.B2(n_637),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1047),
.B(n_960),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1081),
.A2(n_772),
.B(n_700),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1056),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1081),
.A2(n_772),
.B(n_881),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1083),
.B(n_307),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1081),
.A2(n_881),
.B(n_655),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1139),
.A2(n_686),
.B(n_687),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1081),
.A2(n_655),
.B(n_637),
.Y(n_1225)
);

NOR2x1_ASAP7_75t_L g1226 ( 
.A(n_967),
.B(n_747),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1136),
.B(n_766),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_SL g1228 ( 
.A(n_1056),
.B(n_325),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1134),
.A2(n_773),
.B(n_766),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_970),
.B(n_93),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1093),
.A2(n_655),
.B(n_637),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1138),
.B(n_783),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1093),
.A2(n_655),
.B(n_637),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_974),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1036),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1116),
.B(n_783),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1093),
.A2(n_1154),
.B(n_1133),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_983),
.B(n_1148),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1134),
.A2(n_788),
.B(n_488),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1036),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1116),
.B(n_686),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1093),
.A2(n_770),
.B1(n_730),
.B2(n_720),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1104),
.A2(n_328),
.A3(n_335),
.B(n_342),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1156),
.B(n_687),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1134),
.A2(n_488),
.B(n_487),
.Y(n_1245)
);

NAND3x1_ASAP7_75t_L g1246 ( 
.A(n_1077),
.B(n_335),
.C(n_328),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1093),
.A2(n_1154),
.B(n_1133),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_L g1248 ( 
.A(n_1056),
.B(n_687),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_974),
.Y(n_1249)
);

INVx4_ASAP7_75t_SL g1250 ( 
.A(n_988),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1079),
.A2(n_496),
.B(n_491),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_996),
.B(n_302),
.C(n_297),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1092),
.A2(n_608),
.B(n_591),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1145),
.A2(n_342),
.A3(n_343),
.B(n_361),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1071),
.B(n_667),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1156),
.B(n_687),
.Y(n_1256)
);

OA22x2_ASAP7_75t_L g1257 ( 
.A1(n_1068),
.A2(n_429),
.B1(n_420),
.B2(n_419),
.Y(n_1257)
);

AOI221x1_ASAP7_75t_L g1258 ( 
.A1(n_1146),
.A2(n_542),
.B1(n_545),
.B2(n_366),
.C(n_370),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1113),
.A2(n_496),
.B(n_491),
.Y(n_1259)
);

OAI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1148),
.A2(n_306),
.B(n_305),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1021),
.A2(n_498),
.B(n_608),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_988),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_992),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_SL g1264 ( 
.A(n_969),
.B(n_778),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_988),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_SL g1266 ( 
.A1(n_1112),
.A2(n_361),
.B(n_343),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1067),
.B(n_309),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1127),
.B(n_696),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1008),
.B(n_542),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1127),
.B(n_696),
.Y(n_1270)
);

AOI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1013),
.A2(n_609),
.B(n_498),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1021),
.A2(n_609),
.B(n_545),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1115),
.A2(n_370),
.B(n_379),
.C(n_392),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_992),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_968),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_985),
.A2(n_696),
.B(n_647),
.Y(n_1276)
);

INVx8_ASAP7_75t_L g1277 ( 
.A(n_1001),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1067),
.B(n_311),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1140),
.A2(n_696),
.B(n_647),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_997),
.B(n_307),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1071),
.B(n_667),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1145),
.B(n_696),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1155),
.A2(n_379),
.A3(n_392),
.B(n_397),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1155),
.B(n_696),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1086),
.B(n_667),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1071),
.B(n_667),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1007),
.A2(n_647),
.B(n_639),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1078),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1102),
.A2(n_647),
.B(n_639),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_980),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1102),
.A2(n_647),
.B(n_639),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1064),
.A2(n_501),
.B(n_500),
.Y(n_1292)
);

CKINVDCx12_ASAP7_75t_R g1293 ( 
.A(n_1088),
.Y(n_1293)
);

AO21x1_ASAP7_75t_L g1294 ( 
.A1(n_1146),
.A2(n_407),
.B(n_397),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_971),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1064),
.A2(n_501),
.B(n_500),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1090),
.A2(n_419),
.B(n_407),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1012),
.B(n_383),
.C(n_337),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1154),
.A2(n_680),
.B(n_770),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1112),
.A2(n_770),
.B1(n_730),
.B2(n_720),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1153),
.A2(n_770),
.B1(n_730),
.B2(n_720),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1091),
.A2(n_420),
.A3(n_8),
.B(n_11),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1103),
.B(n_667),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1090),
.A2(n_717),
.B(n_770),
.Y(n_1304)
);

CKINVDCx6p67_ASAP7_75t_R g1305 ( 
.A(n_1060),
.Y(n_1305)
);

BUFx2_ASAP7_75t_SL g1306 ( 
.A(n_1001),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_973),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1105),
.B(n_680),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1094),
.A2(n_1101),
.B(n_1128),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_SL g1310 ( 
.A1(n_969),
.A2(n_129),
.B(n_213),
.Y(n_1310)
);

O2A1O1Ixp5_ASAP7_75t_L g1311 ( 
.A1(n_1133),
.A2(n_730),
.B(n_720),
.C(n_717),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_977),
.Y(n_1312)
);

BUFx4_ASAP7_75t_SL g1313 ( 
.A(n_1045),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_997),
.B(n_680),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1109),
.B(n_680),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1094),
.A2(n_778),
.B(n_730),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_980),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_997),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1144),
.A2(n_778),
.B(n_720),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1099),
.B(n_307),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1101),
.A2(n_778),
.B(n_717),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1128),
.A2(n_717),
.B(n_680),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1108),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_978),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1124),
.A2(n_778),
.B(n_717),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1189),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1197),
.A2(n_1132),
.B(n_1043),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1159),
.B(n_995),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1238),
.B(n_1102),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1251),
.A2(n_1157),
.B(n_1147),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1197),
.A2(n_1066),
.B(n_1010),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1201),
.A2(n_1115),
.B1(n_1016),
.B2(n_1084),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1277),
.B(n_1106),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1175),
.B(n_995),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1162),
.A2(n_1008),
.B1(n_1108),
.B2(n_1085),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1180),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1158),
.A2(n_1118),
.B1(n_987),
.B2(n_990),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1325),
.A2(n_1066),
.B(n_1010),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1275),
.Y(n_1340)
);

BUFx4f_ASAP7_75t_SL g1341 ( 
.A(n_1305),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1183),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1287),
.A2(n_1149),
.B(n_1150),
.Y(n_1343)
);

OR2x6_ASAP7_75t_L g1344 ( 
.A(n_1277),
.B(n_1214),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1234),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1163),
.A2(n_1008),
.B1(n_1085),
.B2(n_1130),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1295),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1170),
.B(n_975),
.Y(n_1348)
);

INVx4_ASAP7_75t_SL g1349 ( 
.A(n_1265),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1325),
.A2(n_1066),
.B(n_1011),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1239),
.A2(n_1011),
.B(n_1002),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1273),
.A2(n_991),
.B(n_993),
.C(n_986),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1234),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_SL g1354 ( 
.A1(n_1294),
.A2(n_1004),
.B(n_1003),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_SL g1355 ( 
.A1(n_1192),
.A2(n_1117),
.B(n_1039),
.C(n_1063),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1318),
.B(n_1314),
.Y(n_1356)
);

NAND2x1_ASAP7_75t_L g1357 ( 
.A(n_1220),
.B(n_969),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1218),
.A2(n_1168),
.B1(n_1118),
.B2(n_1196),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1249),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1307),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1198),
.B(n_1070),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1239),
.A2(n_1229),
.B(n_1245),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1318),
.B(n_1032),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1218),
.A2(n_1208),
.B1(n_1176),
.B2(n_1202),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1237),
.A2(n_999),
.B(n_994),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1181),
.A2(n_1150),
.B(n_1055),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1251),
.A2(n_1054),
.B(n_1050),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1312),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1161),
.A2(n_1048),
.A3(n_1049),
.B(n_1002),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1241),
.A2(n_1024),
.B(n_1009),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1187),
.B(n_1026),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1229),
.A2(n_1034),
.B(n_1019),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1262),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1273),
.A2(n_1005),
.B(n_1023),
.C(n_1028),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1236),
.B(n_964),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1245),
.A2(n_1034),
.B(n_1019),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1220),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1216),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1265),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1249),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1267),
.A2(n_1038),
.B1(n_1032),
.B2(n_1042),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1206),
.A2(n_1049),
.B(n_1048),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1324),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1259),
.A2(n_1076),
.B(n_1062),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1172),
.Y(n_1385)
);

NOR4xp25_ASAP7_75t_L g1386 ( 
.A(n_1192),
.B(n_1015),
.C(n_965),
.D(n_1051),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1179),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1290),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1258),
.A2(n_1051),
.A3(n_1062),
.B(n_1098),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1290),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1182),
.A2(n_1082),
.B1(n_1106),
.B2(n_1042),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1213),
.A2(n_1027),
.B(n_1025),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1262),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1199),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1288),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1199),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1194),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1269),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1188),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1212),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1265),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1304),
.A2(n_1322),
.B(n_1321),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1185),
.B(n_1227),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1220),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1271),
.A2(n_1088),
.B(n_1070),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1317),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1316),
.A2(n_1027),
.B(n_1025),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1207),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1262),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1232),
.B(n_1137),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1267),
.B(n_1137),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1165),
.A2(n_1088),
.B(n_1098),
.Y(n_1412)
);

INVx5_ASAP7_75t_L g1413 ( 
.A(n_1265),
.Y(n_1413)
);

NAND2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1262),
.B(n_994),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1314),
.B(n_1032),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1220),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1278),
.B(n_1137),
.Y(n_1417)
);

CKINVDCx16_ASAP7_75t_R g1418 ( 
.A(n_1188),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1313),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1316),
.A2(n_1020),
.B(n_989),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1244),
.A2(n_1040),
.B(n_1038),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1321),
.A2(n_1020),
.B(n_989),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1263),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1310),
.A2(n_999),
.B(n_994),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1160),
.A2(n_1020),
.B(n_989),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1163),
.B(n_976),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1207),
.Y(n_1427)
);

AOI222xp33_ASAP7_75t_L g1428 ( 
.A1(n_1260),
.A2(n_355),
.B1(n_307),
.B2(n_377),
.C1(n_1130),
.C2(n_1119),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1296),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_SL g1430 ( 
.A1(n_1203),
.A2(n_1107),
.B(n_1100),
.C(n_1033),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1259),
.A2(n_1150),
.B(n_1035),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1166),
.A2(n_1107),
.B(n_1100),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1292),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1278),
.A2(n_1038),
.B(n_1042),
.C(n_1088),
.Y(n_1434)
);

NAND2xp33_ASAP7_75t_R g1435 ( 
.A(n_1323),
.B(n_1119),
.Y(n_1435)
);

OAI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1252),
.A2(n_1075),
.B1(n_1060),
.B2(n_315),
.C(n_388),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1314),
.B(n_999),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1160),
.A2(n_1033),
.B(n_1031),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1164),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_SL g1440 ( 
.A(n_1306),
.B(n_1106),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1193),
.A2(n_1036),
.B1(n_976),
.B2(n_1075),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1313),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1177),
.A2(n_1017),
.B1(n_1106),
.B2(n_976),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1256),
.A2(n_1000),
.B(n_1080),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1280),
.B(n_1017),
.Y(n_1445)
);

NOR2x1_ASAP7_75t_L g1446 ( 
.A(n_1298),
.B(n_1052),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1215),
.A2(n_1031),
.B(n_1037),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1200),
.A2(n_1080),
.B(n_1089),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1222),
.A2(n_1137),
.B1(n_1017),
.B2(n_1082),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1323),
.Y(n_1450)
);

OAI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1320),
.A2(n_380),
.B(n_322),
.C(n_324),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1200),
.A2(n_1037),
.B(n_1041),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1247),
.A2(n_1123),
.B(n_1037),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1235),
.Y(n_1454)
);

NAND4xp25_ASAP7_75t_L g1455 ( 
.A(n_1186),
.B(n_1087),
.C(n_377),
.D(n_355),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1235),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1311),
.A2(n_1184),
.B(n_1261),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1207),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1184),
.A2(n_1041),
.B(n_1096),
.Y(n_1459)
);

NOR4xp25_ASAP7_75t_L g1460 ( 
.A(n_1246),
.B(n_1052),
.C(n_1096),
.D(n_1041),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1277),
.Y(n_1461)
);

AO31x2_ASAP7_75t_L g1462 ( 
.A1(n_1301),
.A2(n_1123),
.A3(n_1096),
.B(n_1052),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1193),
.A2(n_1082),
.B1(n_1089),
.B2(n_1080),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1207),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1261),
.A2(n_1123),
.B(n_1029),
.Y(n_1465)
);

AOI21xp33_ASAP7_75t_L g1466 ( 
.A1(n_1268),
.A2(n_1082),
.B(n_1089),
.Y(n_1466)
);

NOR2x1_ASAP7_75t_R g1467 ( 
.A(n_1263),
.B(n_1123),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1309),
.A2(n_1046),
.B(n_1029),
.Y(n_1468)
);

NOR2xp67_ASAP7_75t_L g1469 ( 
.A(n_1274),
.B(n_1018),
.Y(n_1469)
);

INVx4_ASAP7_75t_L g1470 ( 
.A(n_1250),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1178),
.A2(n_375),
.B(n_327),
.Y(n_1471)
);

BUFx10_ASAP7_75t_L g1472 ( 
.A(n_1274),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1211),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1211),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1309),
.A2(n_1046),
.B(n_1029),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1167),
.A2(n_1046),
.B(n_1029),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1292),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1204),
.A2(n_374),
.B(n_338),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1250),
.B(n_1018),
.Y(n_1479)
);

AOI222xp33_ASAP7_75t_L g1480 ( 
.A1(n_1230),
.A2(n_355),
.B1(n_377),
.B2(n_426),
.C1(n_425),
.C2(n_421),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1209),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1226),
.A2(n_1046),
.B1(n_1018),
.B2(n_355),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1297),
.A2(n_1018),
.B(n_647),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1195),
.B(n_320),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1272),
.A2(n_639),
.B(n_211),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1272),
.A2(n_639),
.B(n_207),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1240),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_L g1488 ( 
.A(n_1164),
.B(n_377),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1211),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1240),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1173),
.A2(n_639),
.B(n_205),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1299),
.A2(n_194),
.B(n_190),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1266),
.A2(n_417),
.B1(n_414),
.B2(n_406),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1171),
.B(n_339),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1253),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1224),
.A2(n_1279),
.B(n_1276),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1254),
.B(n_402),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1254),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1223),
.A2(n_163),
.B(n_159),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1253),
.Y(n_1500)
);

NAND2x1p5_ASAP7_75t_L g1501 ( 
.A(n_1228),
.B(n_99),
.Y(n_1501)
);

NOR2xp67_ASAP7_75t_L g1502 ( 
.A(n_1282),
.B(n_101),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1496),
.A2(n_1205),
.B(n_1248),
.C(n_1270),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1356),
.B(n_1250),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1356),
.B(n_1195),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1394),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1399),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1394),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1457),
.A2(n_1253),
.B(n_1221),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1337),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1413),
.B(n_1203),
.Y(n_1511)
);

AOI21xp33_ASAP7_75t_L g1512 ( 
.A1(n_1364),
.A2(n_1217),
.B(n_1284),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1398),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1337),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1395),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1356),
.B(n_1255),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1348),
.A2(n_1293),
.B1(n_365),
.B2(n_353),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1428),
.A2(n_1246),
.B1(n_1257),
.B2(n_1205),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1340),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1333),
.A2(n_340),
.B1(n_384),
.B2(n_386),
.C(n_387),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1480),
.A2(n_1257),
.B1(n_1484),
.B2(n_1361),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1330),
.B(n_1254),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1361),
.A2(n_345),
.B1(n_381),
.B2(n_372),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1363),
.B(n_1255),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1371),
.B(n_1330),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1347),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1381),
.A2(n_1291),
.B1(n_1289),
.B2(n_1308),
.Y(n_1527)
);

NAND2x1p5_ASAP7_75t_L g1528 ( 
.A(n_1413),
.B(n_1281),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1412),
.A2(n_1286),
.B(n_1281),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1360),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1368),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1453),
.A2(n_1248),
.B(n_1264),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1494),
.A2(n_349),
.B1(n_369),
.B2(n_363),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1411),
.B(n_1254),
.Y(n_1534)
);

BUFx4f_ASAP7_75t_SL g1535 ( 
.A(n_1423),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1426),
.A2(n_352),
.B1(n_399),
.B2(n_360),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1363),
.B(n_1286),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1383),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1342),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1329),
.B(n_1417),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1481),
.A2(n_1497),
.B1(n_1358),
.B2(n_1335),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1434),
.A2(n_1315),
.B(n_1303),
.C(n_1285),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1385),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1336),
.A2(n_1449),
.B1(n_1463),
.B2(n_1443),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1457),
.A2(n_1231),
.B(n_1233),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1387),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1413),
.B(n_1470),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1441),
.A2(n_1300),
.B1(n_1242),
.B2(n_1225),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1378),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1362),
.A2(n_1210),
.B(n_1174),
.Y(n_1550)
);

BUFx2_ASAP7_75t_R g1551 ( 
.A(n_1396),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1397),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1497),
.A2(n_354),
.B1(n_356),
.B2(n_1319),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1418),
.B(n_1283),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1400),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1445),
.Y(n_1556)
);

BUFx4_ASAP7_75t_SL g1557 ( 
.A(n_1399),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1433),
.A2(n_1319),
.B(n_1219),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1403),
.A2(n_1302),
.B1(n_1283),
.B2(n_1243),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1406),
.Y(n_1560)
);

AOI21xp33_ASAP7_75t_L g1561 ( 
.A1(n_1391),
.A2(n_1243),
.B(n_1190),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1461),
.Y(n_1562)
);

OAI211xp5_ASAP7_75t_L g1563 ( 
.A1(n_1493),
.A2(n_1302),
.B(n_1243),
.C(n_1283),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1470),
.A2(n_1414),
.B(n_1467),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1461),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1345),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1362),
.A2(n_1169),
.B(n_1191),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1403),
.A2(n_1302),
.B1(n_1243),
.B2(n_11),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1363),
.B(n_1191),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1346),
.A2(n_1191),
.B1(n_1302),
.B2(n_13),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1415),
.B(n_1191),
.Y(n_1571)
);

AOI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1405),
.A2(n_126),
.B(n_153),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1375),
.B(n_5),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1482),
.A2(n_8),
.B1(n_15),
.B2(n_16),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1396),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1415),
.B(n_17),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1344),
.B(n_156),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_R g1578 ( 
.A(n_1334),
.B(n_145),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1353),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1415),
.B(n_1375),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1341),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1370),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1353),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1488),
.A2(n_1498),
.B1(n_1354),
.B2(n_1455),
.Y(n_1584)
);

XOR2xp5_ASAP7_75t_L g1585 ( 
.A(n_1450),
.B(n_144),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1365),
.A2(n_143),
.B(n_133),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1359),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1410),
.B(n_21),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1450),
.B(n_25),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1410),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1436),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1355),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_1592)
);

OAI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1451),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.C(n_40),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1456),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1487),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1359),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1380),
.Y(n_1597)
);

BUFx8_ASAP7_75t_SL g1598 ( 
.A(n_1423),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1490),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1334),
.B(n_130),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1380),
.B(n_48),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1470),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_SL g1603 ( 
.A1(n_1352),
.A2(n_1374),
.B(n_1466),
.C(n_1421),
.Y(n_1603)
);

AND2x2_ASAP7_75t_SL g1604 ( 
.A(n_1460),
.B(n_49),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1388),
.B(n_50),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1388),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1390),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1456),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1419),
.B(n_52),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1442),
.B(n_52),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1334),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1334),
.B(n_124),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1344),
.B(n_1377),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1454),
.B(n_56),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1390),
.B(n_57),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1352),
.A2(n_1374),
.B1(n_1344),
.B2(n_1338),
.Y(n_1616)
);

NAND2x2_ASAP7_75t_L g1617 ( 
.A(n_1487),
.B(n_58),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1343),
.A2(n_122),
.B(n_121),
.Y(n_1618)
);

INVx8_ASAP7_75t_L g1619 ( 
.A(n_1413),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1472),
.Y(n_1620)
);

NOR2xp67_ASAP7_75t_L g1621 ( 
.A(n_1377),
.B(n_113),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1413),
.B(n_109),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1326),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_R g1624 ( 
.A(n_1435),
.B(n_108),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1490),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1389),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1373),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1472),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1327),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1369),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1446),
.A2(n_59),
.B(n_60),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1344),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1377),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1389),
.Y(n_1634)
);

AO21x2_ASAP7_75t_L g1635 ( 
.A1(n_1477),
.A2(n_103),
.B(n_68),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1479),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1469),
.B(n_1386),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1379),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1501),
.A2(n_1444),
.B1(n_1366),
.B2(n_1502),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1479),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1501),
.A2(n_65),
.B1(n_71),
.B2(n_74),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1472),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1369),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1366),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1369),
.Y(n_1645)
);

BUFx12f_ASAP7_75t_L g1646 ( 
.A(n_1416),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1343),
.A2(n_1355),
.B(n_1430),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1440),
.B(n_80),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1439),
.B(n_83),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1404),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1439),
.B(n_87),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1404),
.B(n_88),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1366),
.A2(n_92),
.B1(n_89),
.B2(n_90),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1404),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1389),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1437),
.A2(n_88),
.B1(n_91),
.B2(n_1393),
.Y(n_1656)
);

A2O1A1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1499),
.A2(n_1492),
.B(n_1491),
.C(n_1475),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1424),
.A2(n_91),
.B1(n_1478),
.B2(n_1427),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1401),
.B(n_1416),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1437),
.A2(n_1393),
.B1(n_1414),
.B2(n_1479),
.Y(n_1660)
);

BUFx2_ASAP7_75t_SL g1661 ( 
.A(n_1373),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1401),
.B(n_1416),
.Y(n_1662)
);

AO21x2_ASAP7_75t_L g1663 ( 
.A1(n_1339),
.A2(n_1350),
.B(n_1343),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1478),
.A2(n_1464),
.B1(n_1458),
.B2(n_1408),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1416),
.B(n_1369),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1373),
.B(n_1409),
.Y(n_1666)
);

OAI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1393),
.A2(n_1409),
.B1(n_1373),
.B2(n_1357),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1349),
.B(n_1478),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1393),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1499),
.A2(n_1409),
.B1(n_1492),
.B2(n_1471),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1430),
.A2(n_1331),
.B(n_1448),
.Y(n_1671)
);

NAND2x1_ASAP7_75t_L g1672 ( 
.A(n_1409),
.B(n_1429),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1471),
.A2(n_1431),
.B1(n_1349),
.B2(n_1491),
.Y(n_1673)
);

NOR2xp67_ASAP7_75t_SL g1674 ( 
.A(n_1471),
.B(n_1367),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1408),
.A2(n_1464),
.B1(n_1458),
.B2(n_1427),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1473),
.A2(n_1489),
.B1(n_1474),
.B2(n_1448),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1349),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1473),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1331),
.A2(n_1448),
.B(n_1432),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1489),
.A2(n_1500),
.B1(n_1495),
.B2(n_1331),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1495),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1462),
.B(n_1500),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1407),
.A2(n_1486),
.B1(n_1485),
.B2(n_1476),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1521),
.A2(n_1367),
.B1(n_1384),
.B2(n_1432),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1590),
.B(n_1554),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_1594),
.B2(n_1593),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1594),
.A2(n_1367),
.B1(n_1432),
.B2(n_1384),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1519),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1592),
.A2(n_1631),
.B(n_1582),
.C(n_1644),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1582),
.A2(n_1384),
.B1(n_1431),
.B2(n_1382),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1599),
.A2(n_1431),
.B1(n_1382),
.B2(n_1376),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1518),
.A2(n_1462),
.B1(n_1376),
.B2(n_1351),
.Y(n_1693)
);

OAI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1533),
.A2(n_1523),
.B(n_1536),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1544),
.A2(n_1392),
.B1(n_1476),
.B2(n_1407),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1526),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1644),
.A2(n_1328),
.B1(n_1351),
.B2(n_1459),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1523),
.A2(n_1462),
.B1(n_1475),
.B2(n_1468),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1533),
.A2(n_1486),
.B1(n_1485),
.B2(n_1392),
.C(n_1328),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1556),
.B(n_1459),
.Y(n_1700)
);

OAI211xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1536),
.A2(n_1425),
.B(n_1438),
.C(n_1452),
.Y(n_1701)
);

INVx4_ASAP7_75t_L g1702 ( 
.A(n_1619),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1530),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1539),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1531),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1513),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1538),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1507),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1543),
.Y(n_1709)
);

BUFx12f_ASAP7_75t_L g1710 ( 
.A(n_1625),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1653),
.A2(n_1372),
.B1(n_1438),
.B2(n_1447),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1517),
.A2(n_1465),
.B1(n_1483),
.B2(n_1447),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1520),
.A2(n_1574),
.B1(n_1653),
.B2(n_1641),
.C(n_1570),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1669),
.Y(n_1714)
);

AOI222xp33_ASAP7_75t_L g1715 ( 
.A1(n_1632),
.A2(n_1420),
.B1(n_1422),
.B2(n_1452),
.C1(n_1332),
.C2(n_1339),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1604),
.A2(n_1422),
.B1(n_1350),
.B2(n_1402),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1611),
.A2(n_1402),
.B1(n_1617),
.B2(n_1541),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_L g1718 ( 
.A(n_1656),
.B(n_1648),
.C(n_1563),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1546),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1552),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1514),
.B(n_1613),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1617),
.A2(n_1541),
.B1(n_1573),
.B2(n_1568),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1568),
.A2(n_1624),
.B1(n_1522),
.B2(n_1553),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1603),
.A2(n_1616),
.B1(n_1512),
.B2(n_1553),
.C(n_1588),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1514),
.B(n_1613),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1619),
.Y(n_1726)
);

BUFx12f_ASAP7_75t_L g1727 ( 
.A(n_1625),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1540),
.B(n_1534),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1510),
.B(n_1549),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1555),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1584),
.A2(n_1628),
.B1(n_1642),
.B2(n_1620),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1624),
.A2(n_1577),
.B1(n_1585),
.B2(n_1589),
.Y(n_1732)
);

BUFx4f_ASAP7_75t_L g1733 ( 
.A(n_1600),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1584),
.A2(n_1628),
.B1(n_1637),
.B2(n_1515),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1577),
.A2(n_1576),
.B1(n_1635),
.B2(n_1610),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1646),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1649),
.B(n_1659),
.Y(n_1737)
);

OAI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1639),
.A2(n_1578),
.B1(n_1658),
.B2(n_1577),
.C(n_1618),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1595),
.A2(n_1575),
.B1(n_1508),
.B2(n_1506),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_1614),
.B2(n_1639),
.C(n_1559),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1608),
.A2(n_1575),
.B1(n_1508),
.B2(n_1506),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1613),
.B(n_1504),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1635),
.A2(n_1600),
.B1(n_1612),
.B2(n_1608),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1559),
.A2(n_1658),
.B1(n_1548),
.B2(n_1651),
.C(n_1609),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1560),
.Y(n_1745)
);

AOI211xp5_ASAP7_75t_L g1746 ( 
.A1(n_1586),
.A2(n_1600),
.B(n_1612),
.C(n_1667),
.Y(n_1746)
);

AOI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1535),
.A2(n_1612),
.B1(n_1571),
.B2(n_1569),
.C1(n_1615),
.C2(n_1601),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1562),
.A2(n_1565),
.B1(n_1551),
.B2(n_1516),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_SL g1749 ( 
.A1(n_1578),
.A2(n_1622),
.B1(n_1505),
.B2(n_1527),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1652),
.B(n_1516),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1504),
.B(n_1636),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1681),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1569),
.A2(n_1605),
.B1(n_1537),
.B2(n_1524),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_L g1754 ( 
.A(n_1670),
.B(n_1673),
.C(n_1542),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1562),
.A2(n_1565),
.B1(n_1516),
.B2(n_1524),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1542),
.A2(n_1647),
.B1(n_1664),
.B2(n_1503),
.C(n_1505),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1638),
.B(n_1566),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1622),
.A2(n_1619),
.B1(n_1660),
.B2(n_1537),
.Y(n_1758)
);

AOI222xp33_ASAP7_75t_L g1759 ( 
.A1(n_1579),
.A2(n_1607),
.B1(n_1583),
.B2(n_1581),
.C1(n_1504),
.C2(n_1621),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1598),
.A2(n_1606),
.B1(n_1596),
.B2(n_1597),
.Y(n_1760)
);

AO21x2_ASAP7_75t_L g1761 ( 
.A1(n_1657),
.A2(n_1671),
.B(n_1679),
.Y(n_1761)
);

OAI211xp5_ASAP7_75t_L g1762 ( 
.A1(n_1664),
.A2(n_1564),
.B(n_1657),
.C(n_1633),
.Y(n_1762)
);

OAI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1681),
.A2(n_1636),
.B1(n_1640),
.B2(n_1677),
.Y(n_1763)
);

AOI22x1_ASAP7_75t_L g1764 ( 
.A1(n_1532),
.A2(n_1668),
.B1(n_1547),
.B2(n_1528),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1598),
.A2(n_1606),
.B1(n_1597),
.B2(n_1596),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1619),
.B(n_1672),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1587),
.A2(n_1654),
.B1(n_1650),
.B2(n_1602),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1503),
.A2(n_1666),
.B1(n_1683),
.B2(n_1511),
.C(n_1528),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1661),
.A2(n_1547),
.B1(n_1602),
.B2(n_1627),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1511),
.A2(n_1675),
.B1(n_1627),
.B2(n_1662),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1646),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1627),
.B(n_1665),
.Y(n_1772)
);

OAI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1627),
.A2(n_1682),
.B1(n_1678),
.B2(n_1557),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1684),
.B(n_1629),
.Y(n_1774)
);

NAND2x1_ASAP7_75t_L g1775 ( 
.A(n_1623),
.B(n_1680),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1529),
.A2(n_1643),
.B1(n_1630),
.B2(n_1645),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1675),
.B(n_1572),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1529),
.A2(n_1634),
.B1(n_1655),
.B2(n_1626),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1676),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1680),
.B(n_1567),
.Y(n_1780)
);

OAI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1674),
.A2(n_1567),
.B1(n_1558),
.B2(n_1663),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1663),
.B(n_1558),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1509),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1545),
.A2(n_1509),
.B(n_1550),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1550),
.A2(n_1591),
.B1(n_1521),
.B2(n_808),
.Y(n_1785)
);

A2O1A1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1521),
.A2(n_1030),
.B(n_792),
.C(n_830),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1521),
.A2(n_1333),
.B1(n_792),
.B2(n_759),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1591),
.A2(n_645),
.B1(n_576),
.B2(n_808),
.C(n_830),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1521),
.A2(n_792),
.B1(n_1348),
.B2(n_830),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1521),
.A2(n_1333),
.B1(n_792),
.B2(n_759),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1594),
.A2(n_1428),
.B(n_576),
.C(n_847),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1521),
.A2(n_792),
.B1(n_1348),
.B2(n_830),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_808),
.B2(n_1594),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1556),
.B(n_1580),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1525),
.B(n_1540),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1646),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1682),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_808),
.B2(n_1594),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_808),
.B2(n_1594),
.Y(n_1799)
);

OAI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1518),
.A2(n_1044),
.B1(n_1593),
.B2(n_1578),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1518),
.A2(n_1044),
.B1(n_1593),
.B2(n_1578),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1556),
.B(n_1580),
.Y(n_1802)
);

OAI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1518),
.A2(n_1044),
.B1(n_1593),
.B2(n_1578),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_808),
.B2(n_1594),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1556),
.B(n_1580),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1532),
.A2(n_1496),
.B(n_1030),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1631),
.A2(n_1044),
.B1(n_890),
.B2(n_792),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1592),
.A2(n_1030),
.B(n_1496),
.C(n_1631),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1521),
.A2(n_1333),
.B1(n_792),
.B2(n_759),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_808),
.B2(n_1594),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1556),
.B(n_1580),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1521),
.A2(n_1333),
.B1(n_792),
.B2(n_759),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_808),
.B2(n_1594),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1591),
.A2(n_645),
.B1(n_576),
.B2(n_808),
.C(n_830),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1521),
.A2(n_792),
.B1(n_830),
.B2(n_800),
.C(n_1044),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1519),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1521),
.A2(n_1333),
.B1(n_792),
.B2(n_759),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1525),
.B(n_1540),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1514),
.B(n_1613),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1521),
.A2(n_1333),
.B1(n_792),
.B2(n_759),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1682),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1519),
.Y(n_1822)
);

OAI211xp5_ASAP7_75t_L g1823 ( 
.A1(n_1594),
.A2(n_1428),
.B(n_830),
.C(n_1480),
.Y(n_1823)
);

AOI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1591),
.A2(n_645),
.B1(n_576),
.B2(n_808),
.C(n_830),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1591),
.A2(n_1521),
.B1(n_808),
.B2(n_1594),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1525),
.B(n_1540),
.Y(n_1826)
);

OAI221xp5_ASAP7_75t_SL g1827 ( 
.A1(n_1594),
.A2(n_1428),
.B1(n_1521),
.B2(n_792),
.C(n_847),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1556),
.B(n_1580),
.Y(n_1828)
);

NOR2xp67_ASAP7_75t_L g1829 ( 
.A(n_1513),
.B(n_1426),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1797),
.Y(n_1830)
);

OAI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1789),
.A2(n_1792),
.B(n_1823),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1774),
.B(n_1797),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1694),
.A2(n_1791),
.B1(n_1687),
.B2(n_1810),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1821),
.B(n_1782),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1783),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1827),
.A2(n_1690),
.B1(n_1687),
.B2(n_1804),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1775),
.Y(n_1837)
);

INVxp67_ASAP7_75t_SL g1838 ( 
.A(n_1821),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1721),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1779),
.B(n_1780),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1745),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1761),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1700),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1793),
.A2(n_1825),
.B1(n_1813),
.B2(n_1810),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1761),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1686),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1784),
.B(n_1695),
.Y(n_1847)
);

NAND2x1p5_ASAP7_75t_L g1848 ( 
.A(n_1806),
.B(n_1764),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1778),
.B(n_1776),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1728),
.B(n_1754),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1689),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1685),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1795),
.B(n_1818),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1696),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1703),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1705),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_SL g1857 ( 
.A1(n_1793),
.A2(n_1813),
.B1(n_1825),
.B2(n_1804),
.C(n_1799),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1757),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1716),
.B(n_1777),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1733),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1719),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1766),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1720),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1756),
.B(n_1772),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1730),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1816),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1707),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1826),
.B(n_1709),
.Y(n_1868)
);

BUFx4f_ASAP7_75t_SL g1869 ( 
.A(n_1708),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1822),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1697),
.B(n_1711),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1693),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1693),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1781),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1697),
.B(n_1711),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1699),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1781),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1691),
.B(n_1698),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1752),
.B(n_1734),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1750),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1766),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1691),
.B(n_1753),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1712),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1753),
.B(n_1688),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1688),
.B(n_1715),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1815),
.B(n_1800),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1740),
.B(n_1794),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1768),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1724),
.B(n_1722),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1725),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1755),
.B(n_1731),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1819),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1802),
.B(n_1805),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1770),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1722),
.B(n_1811),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1701),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1766),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1729),
.B(n_1828),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1706),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1692),
.B(n_1737),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1762),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1773),
.B(n_1744),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1763),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1763),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1773),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1735),
.B(n_1743),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1749),
.B(n_1717),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1717),
.B(n_1760),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1742),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1760),
.B(n_1765),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1765),
.B(n_1735),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1767),
.B(n_1690),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1742),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1723),
.B(n_1747),
.Y(n_1914)
);

INVx2_ASAP7_75t_SL g1915 ( 
.A(n_1796),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1843),
.B(n_1714),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1831),
.A2(n_1788),
.B1(n_1814),
.B2(n_1824),
.C(n_1790),
.Y(n_1917)
);

OAI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1831),
.A2(n_1807),
.B1(n_1799),
.B2(n_1798),
.C(n_1786),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1863),
.Y(n_1919)
);

AOI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1836),
.A2(n_1809),
.B1(n_1787),
.B2(n_1820),
.C(n_1812),
.Y(n_1920)
);

AOI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1836),
.A2(n_1817),
.B1(n_1801),
.B2(n_1803),
.C(n_1800),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1850),
.B(n_1801),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1863),
.Y(n_1923)
);

OAI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1889),
.A2(n_1803),
.B1(n_1738),
.B2(n_1713),
.Y(n_1924)
);

AOI222xp33_ASAP7_75t_L g1925 ( 
.A1(n_1833),
.A2(n_1798),
.B1(n_1785),
.B2(n_1723),
.C1(n_1808),
.C2(n_1732),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1867),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1886),
.B(n_1718),
.C(n_1785),
.Y(n_1927)
);

AOI221xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1833),
.A2(n_1889),
.B1(n_1844),
.B2(n_1914),
.C(n_1886),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1844),
.A2(n_1732),
.B1(n_1733),
.B2(n_1746),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1843),
.B(n_1704),
.Y(n_1930)
);

INVxp67_ASAP7_75t_SL g1931 ( 
.A(n_1830),
.Y(n_1931)
);

OAI31xp33_ASAP7_75t_L g1932 ( 
.A1(n_1857),
.A2(n_1914),
.A3(n_1901),
.B(n_1907),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1857),
.A2(n_1901),
.B1(n_1902),
.B2(n_1914),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1863),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1902),
.A2(n_1808),
.B1(n_1829),
.B2(n_1758),
.C(n_1748),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1865),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1869),
.Y(n_1937)
);

OAI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1912),
.A2(n_1739),
.B1(n_1702),
.B2(n_1726),
.Y(n_1938)
);

OR2x6_ASAP7_75t_L g1939 ( 
.A(n_1837),
.B(n_1796),
.Y(n_1939)
);

AOI21x1_ASAP7_75t_L g1940 ( 
.A1(n_1905),
.A2(n_1751),
.B(n_1759),
.Y(n_1940)
);

OAI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1912),
.A2(n_1796),
.B1(n_1727),
.B2(n_1710),
.Y(n_1941)
);

OAI322xp33_ASAP7_75t_L g1942 ( 
.A1(n_1850),
.A2(n_1741),
.A3(n_1736),
.B1(n_1771),
.B2(n_1796),
.C1(n_1769),
.C2(n_1767),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1899),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1865),
.Y(n_1944)
);

OAI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1888),
.A2(n_1736),
.B1(n_1771),
.B2(n_1751),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1865),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1907),
.A2(n_1888),
.B1(n_1908),
.B2(n_1911),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1866),
.Y(n_1948)
);

NAND4xp25_ASAP7_75t_L g1949 ( 
.A(n_1850),
.B(n_1895),
.C(n_1899),
.D(n_1879),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1851),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1839),
.Y(n_1951)
);

OAI33xp33_ASAP7_75t_L g1952 ( 
.A1(n_1895),
.A2(n_1879),
.A3(n_1846),
.B1(n_1834),
.B2(n_1872),
.B3(n_1873),
.Y(n_1952)
);

NAND4xp25_ASAP7_75t_SL g1953 ( 
.A(n_1907),
.B(n_1906),
.C(n_1888),
.D(n_1864),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1830),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1888),
.A2(n_1906),
.B1(n_1864),
.B2(n_1872),
.C(n_1885),
.Y(n_1955)
);

AND2x6_ASAP7_75t_SL g1956 ( 
.A(n_1869),
.B(n_1887),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1915),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1866),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1879),
.B(n_1864),
.Y(n_1959)
);

NOR2x1p5_ASAP7_75t_L g1960 ( 
.A(n_1910),
.B(n_1862),
.Y(n_1960)
);

NAND4xp25_ASAP7_75t_L g1961 ( 
.A(n_1894),
.B(n_1887),
.C(n_1885),
.D(n_1876),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1908),
.A2(n_1911),
.B(n_1905),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1905),
.A2(n_1910),
.B1(n_1891),
.B2(n_1908),
.Y(n_1963)
);

AOI221xp5_ASAP7_75t_L g1964 ( 
.A1(n_1885),
.A2(n_1873),
.B1(n_1876),
.B2(n_1852),
.C(n_1878),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1876),
.A2(n_1910),
.B1(n_1883),
.B2(n_1894),
.C(n_1852),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1897),
.B(n_1909),
.Y(n_1966)
);

OAI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1876),
.A2(n_1883),
.B1(n_1848),
.B2(n_1873),
.C(n_1911),
.Y(n_1967)
);

OA21x2_ASAP7_75t_L g1968 ( 
.A1(n_1842),
.A2(n_1845),
.B(n_1877),
.Y(n_1968)
);

BUFx4f_ASAP7_75t_L g1969 ( 
.A(n_1860),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1834),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1891),
.A2(n_1853),
.B1(n_1904),
.B2(n_1903),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1843),
.B(n_1898),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1853),
.B(n_1846),
.Y(n_1973)
);

AO21x2_ASAP7_75t_L g1974 ( 
.A1(n_1842),
.A2(n_1874),
.B(n_1877),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1880),
.B(n_1909),
.Y(n_1975)
);

OAI33xp33_ASAP7_75t_L g1976 ( 
.A1(n_1834),
.A2(n_1868),
.A3(n_1854),
.B1(n_1855),
.B2(n_1856),
.B3(n_1841),
.Y(n_1976)
);

NAND4xp25_ASAP7_75t_L g1977 ( 
.A(n_1887),
.B(n_1896),
.C(n_1840),
.D(n_1868),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1866),
.Y(n_1978)
);

OA21x2_ASAP7_75t_L g1979 ( 
.A1(n_1842),
.A2(n_1845),
.B(n_1874),
.Y(n_1979)
);

INVxp67_ASAP7_75t_L g1980 ( 
.A(n_1870),
.Y(n_1980)
);

AOI31xp33_ASAP7_75t_L g1981 ( 
.A1(n_1891),
.A2(n_1837),
.A3(n_1900),
.B(n_1878),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1835),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1839),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1897),
.B(n_1913),
.Y(n_1984)
);

AO21x2_ASAP7_75t_L g1985 ( 
.A1(n_1842),
.A2(n_1877),
.B(n_1874),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1861),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1982),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1982),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1975),
.B(n_1859),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1960),
.B(n_1837),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1966),
.B(n_1859),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1966),
.B(n_1859),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1984),
.B(n_1890),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1937),
.B(n_1898),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1970),
.B(n_1840),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1986),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1984),
.B(n_1972),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1939),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1970),
.B(n_1858),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1959),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1950),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1959),
.B(n_1840),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1954),
.B(n_1858),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1980),
.B(n_1838),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1951),
.B(n_1890),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1973),
.B(n_1893),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1919),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1923),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1934),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1954),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1936),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1980),
.B(n_1838),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1944),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1983),
.B(n_1892),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1968),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1943),
.B(n_1916),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1968),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1946),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1968),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1948),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1931),
.B(n_1883),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1930),
.B(n_1892),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1958),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1978),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1979),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_R g2026 ( 
.A(n_1956),
.B(n_1860),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1931),
.Y(n_2027)
);

OR2x6_ASAP7_75t_L g2028 ( 
.A(n_1939),
.B(n_1848),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1949),
.B(n_1883),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1979),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1971),
.B(n_1832),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1971),
.B(n_1832),
.Y(n_2032)
);

AND2x2_ASAP7_75t_SL g2033 ( 
.A(n_1922),
.B(n_1845),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1926),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1974),
.Y(n_2035)
);

AND2x4_ASAP7_75t_SL g2036 ( 
.A(n_1939),
.B(n_1860),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1974),
.B(n_1832),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1985),
.B(n_1892),
.Y(n_2038)
);

NAND4xp25_ASAP7_75t_L g2039 ( 
.A(n_2029),
.B(n_1917),
.C(n_1932),
.D(n_1927),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1996),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2030),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1996),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_2037),
.B(n_2031),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2007),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1991),
.B(n_1979),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_2026),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1991),
.B(n_1913),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_2000),
.B(n_1933),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2007),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2037),
.B(n_2031),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1992),
.B(n_1913),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2008),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2008),
.Y(n_2053)
);

INVxp67_ASAP7_75t_SL g2054 ( 
.A(n_2035),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1992),
.B(n_1913),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2000),
.B(n_1964),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2030),
.Y(n_2057)
);

OR2x2_ASAP7_75t_L g2058 ( 
.A(n_2032),
.B(n_1977),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1994),
.B(n_1961),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2030),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2033),
.B(n_1990),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2032),
.B(n_1985),
.Y(n_2062)
);

NOR5xp2_ASAP7_75t_L g2063 ( 
.A(n_2027),
.B(n_1918),
.C(n_1967),
.D(n_1942),
.E(n_1965),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2033),
.B(n_1847),
.Y(n_2064)
);

NOR2x1p5_ASAP7_75t_L g2065 ( 
.A(n_2029),
.B(n_1940),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2033),
.A2(n_1924),
.B1(n_1947),
.B2(n_1921),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2009),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2009),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2011),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2011),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2013),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2013),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1990),
.B(n_1847),
.Y(n_2073)
);

NOR2x1_ASAP7_75t_L g2074 ( 
.A(n_1998),
.B(n_2027),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1990),
.B(n_1847),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1990),
.B(n_1847),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1989),
.B(n_1847),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2018),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2015),
.Y(n_2079)
);

INVxp33_ASAP7_75t_L g2080 ( 
.A(n_2006),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1989),
.B(n_1847),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2018),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1997),
.B(n_1957),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1995),
.B(n_1981),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_2010),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_1995),
.B(n_1880),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1997),
.B(n_1957),
.Y(n_2087)
);

INVx1_ASAP7_75t_SL g2088 ( 
.A(n_2003),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2020),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2020),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_2028),
.B(n_1862),
.Y(n_2091)
);

NOR3xp33_ASAP7_75t_SL g2092 ( 
.A(n_2039),
.B(n_1941),
.C(n_1953),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2044),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2048),
.B(n_1962),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2061),
.B(n_1998),
.Y(n_2095)
);

INVx1_ASAP7_75t_SL g2096 ( 
.A(n_2046),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2041),
.Y(n_2097)
);

OAI31xp33_ASAP7_75t_L g2098 ( 
.A1(n_2066),
.A2(n_1924),
.A3(n_1929),
.B(n_1941),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2041),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2044),
.Y(n_2100)
);

AND2x4_ASAP7_75t_SL g2101 ( 
.A(n_2061),
.B(n_2028),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2049),
.Y(n_2102)
);

AOI31xp33_ASAP7_75t_L g2103 ( 
.A1(n_2066),
.A2(n_2063),
.A3(n_1928),
.B(n_2056),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2048),
.B(n_2002),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2056),
.B(n_2002),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2049),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_2039),
.B(n_1922),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2059),
.B(n_1955),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2041),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2088),
.B(n_1999),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2059),
.B(n_1963),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_2064),
.B(n_1938),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2057),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2073),
.B(n_2005),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2052),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2080),
.B(n_2058),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2052),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_2074),
.B(n_2028),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_2057),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2058),
.B(n_2065),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2053),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2053),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2074),
.B(n_2028),
.Y(n_2123)
);

OAI221xp5_ASAP7_75t_L g2124 ( 
.A1(n_2084),
.A2(n_2043),
.B1(n_2050),
.B2(n_1920),
.C(n_1925),
.Y(n_2124)
);

CKINVDCx16_ASAP7_75t_R g2125 ( 
.A(n_2064),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2067),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2073),
.B(n_2005),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2067),
.Y(n_2128)
);

NAND2xp33_ASAP7_75t_R g2129 ( 
.A(n_2063),
.B(n_1862),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2075),
.B(n_2014),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2088),
.B(n_1999),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2068),
.Y(n_2132)
);

BUFx2_ASAP7_75t_L g2133 ( 
.A(n_2085),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2065),
.B(n_2043),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2075),
.B(n_2014),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2076),
.B(n_2016),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2050),
.B(n_2022),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2076),
.B(n_2016),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2068),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2077),
.B(n_1993),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_2129),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2133),
.Y(n_2142)
);

AOI21xp33_ASAP7_75t_L g2143 ( 
.A1(n_2103),
.A2(n_2062),
.B(n_1938),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2093),
.Y(n_2144)
);

CKINVDCx14_ASAP7_75t_R g2145 ( 
.A(n_2107),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_2108),
.B(n_2096),
.Y(n_2146)
);

O2A1O1Ixp33_ASAP7_75t_SL g2147 ( 
.A1(n_2094),
.A2(n_2085),
.B(n_2084),
.C(n_2062),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2098),
.A2(n_1952),
.B(n_1935),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2125),
.A2(n_2028),
.B1(n_2036),
.B2(n_2091),
.Y(n_2149)
);

AOI221xp5_ASAP7_75t_L g2150 ( 
.A1(n_2124),
.A2(n_1976),
.B1(n_2054),
.B2(n_2045),
.C(n_2082),
.Y(n_2150)
);

INVxp67_ASAP7_75t_L g2151 ( 
.A(n_2116),
.Y(n_2151)
);

INVxp67_ASAP7_75t_L g2152 ( 
.A(n_2120),
.Y(n_2152)
);

INVx1_ASAP7_75t_SL g2153 ( 
.A(n_2095),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2093),
.Y(n_2154)
);

AO221x1_ASAP7_75t_L g2155 ( 
.A1(n_2133),
.A2(n_1945),
.B1(n_2057),
.B2(n_2060),
.C(n_2069),
.Y(n_2155)
);

AOI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2125),
.A2(n_2091),
.B1(n_1878),
.B2(n_1875),
.Y(n_2156)
);

INVx1_ASAP7_75t_SL g2157 ( 
.A(n_2095),
.Y(n_2157)
);

OAI22xp5_ASAP7_75t_SL g2158 ( 
.A1(n_2111),
.A2(n_2091),
.B1(n_1848),
.B2(n_1860),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2092),
.A2(n_2036),
.B1(n_2091),
.B2(n_1969),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2100),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_SL g2161 ( 
.A1(n_2098),
.A2(n_1875),
.B(n_1871),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2104),
.B(n_2105),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2136),
.B(n_2138),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2100),
.Y(n_2164)
);

OA21x2_ASAP7_75t_L g2165 ( 
.A1(n_2097),
.A2(n_2054),
.B(n_2079),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2102),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2134),
.B(n_2077),
.Y(n_2167)
);

OAI322xp33_ASAP7_75t_L g2168 ( 
.A1(n_2112),
.A2(n_2021),
.A3(n_2003),
.B1(n_2035),
.B2(n_2089),
.C1(n_2069),
.C2(n_2070),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2136),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2138),
.B(n_2081),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2102),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2106),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2106),
.Y(n_2173)
);

NOR2x1_ASAP7_75t_L g2174 ( 
.A(n_2118),
.B(n_2060),
.Y(n_2174)
);

OAI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_2110),
.A2(n_1896),
.B1(n_1904),
.B2(n_1903),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_R g2176 ( 
.A(n_2118),
.B(n_1915),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2115),
.Y(n_2177)
);

OAI32xp33_ASAP7_75t_L g2178 ( 
.A1(n_2110),
.A2(n_2019),
.A3(n_2025),
.B1(n_2015),
.B2(n_2017),
.Y(n_2178)
);

INVxp33_ASAP7_75t_L g2179 ( 
.A(n_2131),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2163),
.Y(n_2180)
);

OAI32xp33_ASAP7_75t_L g2181 ( 
.A1(n_2141),
.A2(n_2131),
.A3(n_2119),
.B1(n_2137),
.B2(n_2017),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_2145),
.A2(n_2123),
.B(n_2118),
.Y(n_2182)
);

OAI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_2145),
.A2(n_2123),
.B(n_2118),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_2146),
.A2(n_2148),
.B1(n_2143),
.B2(n_2151),
.Y(n_2184)
);

O2A1O1Ixp5_ASAP7_75t_L g2185 ( 
.A1(n_2168),
.A2(n_2123),
.B(n_2109),
.C(n_2099),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_2146),
.B(n_2152),
.Y(n_2186)
);

NOR4xp25_ASAP7_75t_L g2187 ( 
.A(n_2147),
.B(n_2113),
.C(n_2109),
.D(n_2099),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2144),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_2161),
.A2(n_2147),
.B(n_2162),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2153),
.B(n_2114),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2154),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_2179),
.B(n_2123),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2157),
.B(n_2114),
.Y(n_2193)
);

OAI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_2156),
.A2(n_2101),
.B1(n_2036),
.B2(n_2127),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2165),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2142),
.B(n_2127),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2169),
.B(n_2130),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2167),
.B(n_2130),
.Y(n_2198)
);

OAI221xp5_ASAP7_75t_L g2199 ( 
.A1(n_2150),
.A2(n_2122),
.B1(n_2139),
.B2(n_2128),
.C(n_2115),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2179),
.A2(n_2117),
.B(n_2139),
.Y(n_2200)
);

INVx2_ASAP7_75t_SL g2201 ( 
.A(n_2174),
.Y(n_2201)
);

AOI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_2155),
.A2(n_2101),
.B(n_2121),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2170),
.B(n_2135),
.Y(n_2203)
);

O2A1O1Ixp33_ASAP7_75t_SL g2204 ( 
.A1(n_2175),
.A2(n_2010),
.B(n_2117),
.C(n_2132),
.Y(n_2204)
);

AOI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_2159),
.A2(n_2101),
.B1(n_1871),
.B2(n_1875),
.Y(n_2205)
);

OAI22xp33_ASAP7_75t_SL g2206 ( 
.A1(n_2149),
.A2(n_2122),
.B1(n_2121),
.B2(n_2126),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_2160),
.B(n_2135),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2164),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_2201),
.Y(n_2209)
);

OAI32xp33_ASAP7_75t_L g2210 ( 
.A1(n_2184),
.A2(n_2172),
.A3(n_2177),
.B1(n_2166),
.B2(n_2171),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2183),
.B(n_2176),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_2182),
.B(n_2176),
.Y(n_2212)
);

INVx1_ASAP7_75t_SL g2213 ( 
.A(n_2192),
.Y(n_2213)
);

XOR2x2_ASAP7_75t_L g2214 ( 
.A(n_2186),
.B(n_2158),
.Y(n_2214)
);

CKINVDCx16_ASAP7_75t_R g2215 ( 
.A(n_2186),
.Y(n_2215)
);

AOI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_2184),
.A2(n_2175),
.B1(n_2173),
.B2(n_2126),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2195),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_2192),
.B(n_2081),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2197),
.B(n_2140),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2189),
.B(n_2140),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2195),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2190),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2188),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2180),
.B(n_2128),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2191),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_2199),
.B(n_2086),
.Y(n_2226)
);

INVxp67_ASAP7_75t_L g2227 ( 
.A(n_2196),
.Y(n_2227)
);

OAI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2187),
.A2(n_2132),
.B1(n_2165),
.B2(n_2099),
.C(n_2113),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_2200),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2193),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2207),
.B(n_2045),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2215),
.B(n_2207),
.Y(n_2232)
);

OAI211xp5_ASAP7_75t_L g2233 ( 
.A1(n_2216),
.A2(n_2229),
.B(n_2210),
.C(n_2213),
.Y(n_2233)
);

OAI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_2220),
.A2(n_2202),
.B1(n_2205),
.B2(n_2228),
.Y(n_2234)
);

NAND4xp25_ASAP7_75t_L g2235 ( 
.A(n_2227),
.B(n_2185),
.C(n_2194),
.D(n_2208),
.Y(n_2235)
);

NAND3xp33_ASAP7_75t_SL g2236 ( 
.A(n_2212),
.B(n_2185),
.C(n_2198),
.Y(n_2236)
);

NOR3xp33_ASAP7_75t_L g2237 ( 
.A(n_2210),
.B(n_2206),
.C(n_2181),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2217),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2209),
.B(n_2203),
.Y(n_2239)
);

AOI32xp33_ASAP7_75t_L g2240 ( 
.A1(n_2211),
.A2(n_2204),
.A3(n_2119),
.B1(n_2045),
.B2(n_2060),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2214),
.A2(n_2178),
.B(n_2113),
.Y(n_2241)
);

INVx1_ASAP7_75t_SL g2242 ( 
.A(n_2211),
.Y(n_2242)
);

NOR3xp33_ASAP7_75t_L g2243 ( 
.A(n_2222),
.B(n_2204),
.C(n_2119),
.Y(n_2243)
);

AND4x1_ASAP7_75t_L g2244 ( 
.A(n_2217),
.B(n_2083),
.C(n_2087),
.D(n_2078),
.Y(n_2244)
);

OAI21xp33_ASAP7_75t_L g2245 ( 
.A1(n_2214),
.A2(n_2109),
.B(n_2097),
.Y(n_2245)
);

OAI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_2226),
.A2(n_2165),
.B(n_2097),
.Y(n_2246)
);

NOR2xp67_ASAP7_75t_L g2247 ( 
.A(n_2209),
.B(n_2119),
.Y(n_2247)
);

OAI211xp5_ASAP7_75t_L g2248 ( 
.A1(n_2233),
.A2(n_2222),
.B(n_2230),
.C(n_2221),
.Y(n_2248)
);

NAND2x1_ASAP7_75t_L g2249 ( 
.A(n_2247),
.B(n_2230),
.Y(n_2249)
);

OAI221xp5_ASAP7_75t_SL g2250 ( 
.A1(n_2237),
.A2(n_2224),
.B1(n_2218),
.B2(n_2221),
.C(n_2223),
.Y(n_2250)
);

AOI322xp5_ASAP7_75t_L g2251 ( 
.A1(n_2234),
.A2(n_2225),
.A3(n_2223),
.B1(n_2219),
.B2(n_2231),
.C1(n_2025),
.C2(n_2019),
.Y(n_2251)
);

OAI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2236),
.A2(n_2225),
.B(n_2219),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_2246),
.A2(n_2243),
.B(n_2241),
.Y(n_2253)
);

AOI221xp5_ASAP7_75t_L g2254 ( 
.A1(n_2235),
.A2(n_2245),
.B1(n_2240),
.B2(n_2242),
.C(n_2232),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_R g2255 ( 
.A(n_2239),
.B(n_2231),
.Y(n_2255)
);

AOI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2238),
.A2(n_2079),
.B1(n_2015),
.B2(n_2025),
.C(n_2017),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2244),
.Y(n_2257)
);

AOI321xp33_ASAP7_75t_L g2258 ( 
.A1(n_2237),
.A2(n_1871),
.A3(n_1945),
.B1(n_1884),
.B2(n_1882),
.C(n_1849),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2233),
.A2(n_2010),
.B1(n_2089),
.B2(n_2071),
.Y(n_2259)
);

AOI222xp33_ASAP7_75t_L g2260 ( 
.A1(n_2236),
.A2(n_2019),
.B1(n_2079),
.B2(n_1896),
.C1(n_1884),
.C2(n_1849),
.Y(n_2260)
);

OAI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2236),
.A2(n_2021),
.B1(n_2012),
.B2(n_2004),
.Y(n_2261)
);

AOI221xp5_ASAP7_75t_L g2262 ( 
.A1(n_2237),
.A2(n_2090),
.B1(n_2082),
.B2(n_2070),
.C(n_2071),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2257),
.B(n_2072),
.Y(n_2263)
);

AOI211xp5_ASAP7_75t_SL g2264 ( 
.A1(n_2248),
.A2(n_1862),
.B(n_1881),
.C(n_2012),
.Y(n_2264)
);

NAND3xp33_ASAP7_75t_L g2265 ( 
.A(n_2262),
.B(n_2090),
.C(n_2078),
.Y(n_2265)
);

AOI222xp33_ASAP7_75t_L g2266 ( 
.A1(n_2253),
.A2(n_2004),
.B1(n_1884),
.B2(n_1849),
.C1(n_1882),
.C2(n_2038),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2249),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_2255),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2254),
.B(n_2252),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2250),
.A2(n_2072),
.B1(n_2042),
.B2(n_2040),
.Y(n_2270)
);

NOR3xp33_ASAP7_75t_L g2271 ( 
.A(n_2259),
.B(n_1915),
.C(n_1862),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2268),
.B(n_2261),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2267),
.B(n_2260),
.Y(n_2273)
);

OAI21xp5_ASAP7_75t_SL g2274 ( 
.A1(n_2269),
.A2(n_2251),
.B(n_2258),
.Y(n_2274)
);

AOI222xp33_ASAP7_75t_L g2275 ( 
.A1(n_2270),
.A2(n_2263),
.B1(n_2265),
.B2(n_2256),
.C1(n_2264),
.C2(n_2266),
.Y(n_2275)
);

O2A1O1Ixp33_ASAP7_75t_L g2276 ( 
.A1(n_2271),
.A2(n_1848),
.B(n_2040),
.C(n_2042),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2268),
.B(n_2083),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2268),
.B(n_2087),
.Y(n_2278)
);

INVx2_ASAP7_75t_SL g2279 ( 
.A(n_2267),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2279),
.Y(n_2280)
);

NOR3xp33_ASAP7_75t_L g2281 ( 
.A(n_2272),
.B(n_1881),
.C(n_1897),
.Y(n_2281)
);

AND2x4_ASAP7_75t_L g2282 ( 
.A(n_2277),
.B(n_2278),
.Y(n_2282)
);

INVx2_ASAP7_75t_SL g2283 ( 
.A(n_2273),
.Y(n_2283)
);

NAND3xp33_ASAP7_75t_SL g2284 ( 
.A(n_2274),
.B(n_1848),
.C(n_2038),
.Y(n_2284)
);

OAI211xp5_ASAP7_75t_SL g2285 ( 
.A1(n_2274),
.A2(n_1881),
.B(n_2086),
.C(n_1897),
.Y(n_2285)
);

AOI22xp33_ASAP7_75t_L g2286 ( 
.A1(n_2275),
.A2(n_1881),
.B1(n_1969),
.B2(n_1860),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2276),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2282),
.B(n_2047),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2283),
.B(n_2047),
.Y(n_2289)
);

AOI211xp5_ASAP7_75t_SL g2290 ( 
.A1(n_2280),
.A2(n_1881),
.B(n_1904),
.C(n_1903),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2282),
.B(n_2051),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2289),
.Y(n_2292)
);

BUFx2_ASAP7_75t_SL g2293 ( 
.A(n_2288),
.Y(n_2293)
);

OAI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2293),
.A2(n_2286),
.B1(n_2287),
.B2(n_2291),
.Y(n_2294)
);

XNOR2x2_ASAP7_75t_L g2295 ( 
.A(n_2292),
.B(n_2284),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2295),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2294),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_2295),
.B(n_2281),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2296),
.B(n_2293),
.Y(n_2299)
);

AOI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2297),
.A2(n_2285),
.B1(n_2290),
.B2(n_2051),
.Y(n_2300)
);

CKINVDCx14_ASAP7_75t_R g2301 ( 
.A(n_2299),
.Y(n_2301)
);

AOI222xp33_ASAP7_75t_SL g2302 ( 
.A1(n_2300),
.A2(n_2298),
.B1(n_1987),
.B2(n_1988),
.C1(n_2023),
.C2(n_2024),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_SL g2303 ( 
.A1(n_2301),
.A2(n_1860),
.B1(n_2001),
.B2(n_1988),
.Y(n_2303)
);

AOI221xp5_ASAP7_75t_L g2304 ( 
.A1(n_2303),
.A2(n_2302),
.B1(n_1987),
.B2(n_2023),
.C(n_2024),
.Y(n_2304)
);

AOI211xp5_ASAP7_75t_L g2305 ( 
.A1(n_2304),
.A2(n_1860),
.B(n_2034),
.C(n_2055),
.Y(n_2305)
);


endmodule