module fake_jpeg_18336_n_142 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_29),
.B1(n_17),
.B2(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_26),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_57),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_22),
.B(n_21),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_58),
.B1(n_39),
.B2(n_40),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.C(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_26),
.B1(n_18),
.B2(n_15),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_72),
.B1(n_55),
.B2(n_4),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_6),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_3),
.B1(n_9),
.B2(n_13),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_13),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_9),
.B(n_77),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_59),
.B(n_44),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_52),
.B1(n_51),
.B2(n_60),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_63),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_55),
.C(n_51),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_90),
.C(n_78),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_91),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_1),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_66),
.B1(n_63),
.B2(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_99),
.C(n_82),
.Y(n_113)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_84),
.B1(n_88),
.B2(n_93),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_80),
.C(n_71),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_110),
.C(n_98),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g106 ( 
.A(n_86),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_119),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_115),
.C(n_118),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_85),
.C(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_96),
.Y(n_119)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_105),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_123),
.B1(n_122),
.B2(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_93),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_100),
.B(n_103),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_110),
.C(n_108),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_108),
.C(n_88),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_129),
.Y(n_132)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_92),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_134),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_95),
.B(n_114),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_127),
.B(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_131),
.B(n_130),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_130),
.C(n_68),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_76),
.C(n_101),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_139),
.B(n_71),
.Y(n_142)
);


endmodule