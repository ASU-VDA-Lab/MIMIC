module fake_jpeg_4273_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_36),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_42),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_63),
.B1(n_57),
.B2(n_67),
.Y(n_95)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_51),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_32),
.C(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_67),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_62),
.B1(n_71),
.B2(n_26),
.Y(n_75)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_54),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_58),
.B1(n_20),
.B2(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_30),
.B1(n_18),
.B2(n_32),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_16),
.B1(n_17),
.B2(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_16),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_89),
.B1(n_97),
.B2(n_25),
.Y(n_127)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_80),
.Y(n_117)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_20),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_99),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_22),
.B1(n_25),
.B2(n_33),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_22),
.B1(n_33),
.B2(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_98),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_123),
.B1(n_125),
.B2(n_79),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_101),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_49),
.B1(n_73),
.B2(n_60),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_107),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_53),
.B1(n_61),
.B2(n_47),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_109),
.B1(n_118),
.B2(n_127),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_63),
.B1(n_52),
.B2(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_82),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_116),
.B(n_43),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_122),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_22),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_74),
.B1(n_66),
.B2(n_54),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_43),
.B(n_34),
.C(n_41),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_73),
.B1(n_49),
.B2(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_88),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_72),
.B1(n_23),
.B2(n_31),
.Y(n_125)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_94),
.B1(n_92),
.B2(n_77),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_129),
.A2(n_140),
.B1(n_143),
.B2(n_145),
.Y(n_185)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_136),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_101),
.B1(n_103),
.B2(n_107),
.Y(n_162)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_50),
.B(n_34),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_21),
.B(n_43),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_39),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_154),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_39),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_119),
.B1(n_114),
.B2(n_116),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_187),
.B(n_152),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_114),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_164),
.C(n_165),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_186),
.B1(n_132),
.B2(n_157),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_125),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_43),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_104),
.B1(n_124),
.B2(n_111),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_169),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_112),
.B1(n_120),
.B2(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_126),
.B1(n_122),
.B2(n_110),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_173),
.B1(n_176),
.B2(n_183),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_34),
.C(n_41),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_151),
.C(n_148),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_138),
.B1(n_136),
.B2(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_179),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_126),
.B1(n_35),
.B2(n_41),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_35),
.C(n_39),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_181),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_131),
.B(n_39),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_35),
.A3(n_45),
.B1(n_31),
.B2(n_23),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_137),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_45),
.B1(n_31),
.B2(n_23),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_143),
.B1(n_135),
.B2(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_31),
.B1(n_33),
.B2(n_25),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_105),
.B1(n_33),
.B2(n_24),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_213),
.B(n_190),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_194),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_196),
.C(n_214),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_195),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_132),
.B1(n_105),
.B2(n_133),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_197),
.A2(n_211),
.B1(n_15),
.B2(n_14),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_204),
.B1(n_208),
.B2(n_166),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_155),
.B(n_157),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_205),
.B(n_209),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_184),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_152),
.B(n_24),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_210),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_24),
.B1(n_15),
.B2(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_0),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_180),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_3),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_238),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_230),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_172),
.B1(n_185),
.B2(n_158),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_229),
.B(n_207),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_165),
.C(n_159),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_235),
.C(n_239),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_181),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_193),
.B(n_164),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_183),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_232),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_201),
.B(n_186),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_191),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_187),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_24),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_194),
.C(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_198),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_192),
.C(n_202),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_250),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_248),
.A2(n_249),
.B(n_252),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_210),
.B1(n_212),
.B2(n_206),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_219),
.A2(n_195),
.B(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_195),
.B1(n_211),
.B2(n_2),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_256),
.B1(n_221),
.B2(n_222),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

XOR2x2_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_232),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_0),
.C(n_3),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_266),
.C(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_3),
.C(n_4),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_260),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_233),
.Y(n_272)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_217),
.C(n_229),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_280),
.C(n_283),
.Y(n_287)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_281),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_231),
.C(n_238),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_225),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_282),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_235),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_254),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_267),
.A2(n_251),
.B1(n_247),
.B2(n_234),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_268),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_243),
.B(n_245),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_291),
.B(n_292),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_242),
.B1(n_255),
.B2(n_249),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_293),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_270),
.B(n_274),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_262),
.B1(n_266),
.B2(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_300),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_12),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_6),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_12),
.B(n_11),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_10),
.Y(n_312)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_275),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_308),
.B(n_287),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_314),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_273),
.B1(n_277),
.B2(n_280),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_309),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_307),
.B(n_311),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_301),
.C(n_288),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_283),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_5),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_6),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_322),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_320),
.B(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_292),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_6),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_296),
.B(n_7),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_324),
.A2(n_312),
.B(n_304),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_6),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_328),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_313),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_332),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_SL g333 ( 
.A(n_317),
.B(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_315),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_336),
.B(n_7),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_327),
.A2(n_330),
.B(n_331),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_8),
.B(n_9),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_340),
.B(n_335),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_337),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_334),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_8),
.B1(n_9),
.B2(n_316),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_9),
.Y(n_345)
);


endmodule