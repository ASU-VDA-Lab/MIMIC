module fake_jpeg_16966_n_210 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_210);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_39),
.B1(n_30),
.B2(n_4),
.Y(n_52)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_20),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_31),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_59),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_21),
.C(n_23),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_17),
.C(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_21),
.B(n_28),
.C(n_19),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_20),
.A3(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_5),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_19),
.B1(n_32),
.B2(n_26),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_0),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_43),
.B(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_42),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_41),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_71),
.B1(n_87),
.B2(n_9),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_52),
.B(n_54),
.C(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_76),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_5),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_79),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_5),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_81),
.B(n_9),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_6),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_7),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_88),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_9),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_104),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_33),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_86),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_82),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_37),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_78),
.C(n_89),
.Y(n_118)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_35),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_15),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_13),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_35),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_61),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_122),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_114),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_123),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_73),
.C(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_107),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_75),
.C(n_84),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_62),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_90),
.C(n_86),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_106),
.B1(n_104),
.B2(n_99),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_70),
.B1(n_81),
.B2(n_79),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_96),
.B1(n_95),
.B2(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_85),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_97),
.C(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_139),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_142),
.C(n_153),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_117),
.C(n_118),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_96),
.C(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_157),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_115),
.C(n_109),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_128),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_116),
.A3(n_111),
.B1(n_92),
.B2(n_71),
.C(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_158),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_106),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_106),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_137),
.B1(n_87),
.B2(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_166),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.C(n_167),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_146),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_136),
.C(n_130),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_156),
.C(n_158),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_105),
.C(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_171),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_143),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_105),
.A3(n_152),
.B1(n_81),
.B2(n_124),
.C1(n_82),
.C2(n_143),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_136),
.B(n_157),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_175),
.A2(n_185),
.B(n_24),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_171),
.C(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_182),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_165),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_183),
.C(n_175),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_65),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_126),
.B(n_119),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_177),
.C(n_185),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_167),
.B1(n_180),
.B2(n_181),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_183),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_161),
.B(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_193),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_164),
.B1(n_119),
.B2(n_90),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_35),
.B1(n_80),
.B2(n_12),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_18),
.B(n_25),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_184),
.B(n_80),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_24),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_201),
.B1(n_10),
.B2(n_11),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_200),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_12),
.B(n_16),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_195),
.B(n_192),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_198),
.Y(n_208)
);

AO31x2_ASAP7_75t_SL g209 ( 
.A1(n_207),
.A2(n_206),
.A3(n_205),
.B(n_198),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_208),
.Y(n_210)
);


endmodule