module fake_jpeg_8689_n_311 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_62),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_34),
.B1(n_22),
.B2(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_56),
.B1(n_30),
.B2(n_42),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_65),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_22),
.B1(n_20),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_61),
.B1(n_44),
.B2(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_30),
.B1(n_20),
.B2(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_71),
.Y(n_105)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_76),
.Y(n_118)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_83),
.B(n_85),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_80),
.B1(n_41),
.B2(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_82),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_81),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_41),
.B1(n_42),
.B2(n_52),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_17),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_43),
.B(n_40),
.C(n_28),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_38),
.B1(n_42),
.B2(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_88),
.Y(n_130)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_17),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_98),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_103),
.Y(n_114)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_43),
.C(n_37),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_37),
.C(n_26),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_113),
.B1(n_119),
.B2(n_124),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_38),
.B1(n_36),
.B2(n_28),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_93),
.B1(n_98),
.B2(n_103),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_38),
.B1(n_29),
.B2(n_35),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_26),
.C(n_76),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_80),
.B1(n_71),
.B2(n_100),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_95),
.B1(n_26),
.B2(n_35),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_114),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_123),
.B1(n_122),
.B2(n_106),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_138),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_83),
.B(n_97),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_137),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_139),
.B1(n_141),
.B2(n_149),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_97),
.B(n_102),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_101),
.B1(n_83),
.B2(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_79),
.B1(n_87),
.B2(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_81),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_148),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_79),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_88),
.B1(n_86),
.B2(n_89),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_70),
.B1(n_73),
.B2(n_18),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_158),
.B1(n_162),
.B2(n_116),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_29),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_152),
.B(n_154),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_122),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_130),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_24),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_159),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_90),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_35),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_26),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_161),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_107),
.A2(n_95),
.B1(n_35),
.B2(n_33),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_163),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

XOR2x1_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_127),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_168),
.A2(n_175),
.B(n_178),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_171),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_115),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_112),
.B(n_129),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_108),
.B(n_112),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_120),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_184),
.B(n_185),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_192),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_115),
.A3(n_120),
.B1(n_108),
.B2(n_123),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_123),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_131),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_109),
.B1(n_106),
.B2(n_131),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_147),
.B1(n_116),
.B2(n_33),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_177),
.A2(n_152),
.B1(n_154),
.B2(n_109),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_176),
.B1(n_179),
.B2(n_173),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_146),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_161),
.B1(n_139),
.B2(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_217),
.B1(n_163),
.B2(n_190),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_151),
.C(n_142),
.Y(n_207)
);

OAI322xp33_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_168),
.A3(n_181),
.B1(n_190),
.B2(n_166),
.C1(n_175),
.C2(n_189),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_153),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_210),
.B(n_214),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_213),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_134),
.Y(n_216)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_145),
.B1(n_158),
.B2(n_147),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_219),
.B1(n_176),
.B2(n_192),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_75),
.B1(n_33),
.B2(n_29),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_221),
.A2(n_229),
.B1(n_232),
.B2(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_170),
.C(n_169),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_227),
.C(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_169),
.C(n_171),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_164),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_237),
.B1(n_218),
.B2(n_203),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_212),
.B(n_164),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_178),
.B(n_182),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_75),
.B1(n_33),
.B2(n_24),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_9),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_26),
.C(n_1),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_0),
.C(n_1),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_201),
.B(n_9),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_7),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_10),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_206),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_240),
.C(n_215),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_259),
.B1(n_7),
.B2(n_14),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_206),
.B1(n_201),
.B2(n_205),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_246),
.A2(n_223),
.B1(n_237),
.B2(n_239),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_214),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_260),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_256),
.B(n_257),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_204),
.B1(n_220),
.B2(n_195),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_230),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_224),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_208),
.B1(n_219),
.B2(n_215),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_225),
.C(n_227),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_270),
.B1(n_246),
.B2(n_245),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_242),
.C(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_233),
.C(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_268),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_1),
.C(n_2),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_260),
.C(n_247),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_10),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_247),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_248),
.B(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_275),
.B(n_279),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_274),
.A2(n_256),
.B(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_282),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_255),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_285),
.C(n_276),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_7),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_286),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_272),
.B(n_263),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_11),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_288),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_261),
.B1(n_3),
.B2(n_2),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_11),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_276),
.B1(n_282),
.B2(n_281),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_5),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_3),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_300),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_3),
.C(n_4),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_5),
.C(n_6),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_288),
.A3(n_289),
.B1(n_6),
.B2(n_13),
.C1(n_14),
.C2(n_16),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_306),
.A3(n_296),
.B1(n_6),
.B2(n_13),
.C1(n_14),
.C2(n_3),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_299),
.B(n_297),
.C(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_303),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_13),
.Y(n_311)
);


endmodule