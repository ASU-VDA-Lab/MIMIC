module real_aes_7044_n_255 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_255);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_255;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_461;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_755;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_769;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_756;
wire n_598;
wire n_404;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_472;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_0), .A2(n_190), .B1(n_296), .B2(n_301), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_1), .Y(n_383) );
XOR2x2_ASAP7_75t_L g520 ( .A(n_2), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_3), .A2(n_17), .B1(n_397), .B2(n_400), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_4), .Y(n_593) );
INVx1_ASAP7_75t_L g796 ( .A(n_5), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_6), .A2(n_167), .B1(n_469), .B2(n_515), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_7), .A2(n_60), .B1(n_524), .B2(n_636), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_8), .A2(n_373), .B1(n_416), .B2(n_417), .Y(n_372) );
INVx1_ASAP7_75t_L g416 ( .A(n_8), .Y(n_416) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_9), .A2(n_29), .B1(n_202), .B2(n_382), .C1(n_542), .C2(n_544), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_10), .A2(n_227), .B1(n_459), .B2(n_462), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_11), .A2(n_107), .B1(n_683), .B2(n_804), .C(n_805), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_12), .A2(n_159), .B1(n_272), .B2(n_530), .Y(n_662) );
INVx1_ASAP7_75t_L g586 ( .A(n_13), .Y(n_586) );
OA22x2_ASAP7_75t_L g551 ( .A1(n_14), .A2(n_552), .B1(n_553), .B2(n_587), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_14), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_15), .A2(n_133), .B1(n_455), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_16), .A2(n_69), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_18), .A2(n_204), .B1(n_612), .B2(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_19), .A2(n_219), .B1(n_403), .B2(n_459), .C(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g806 ( .A(n_20), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_21), .A2(n_68), .B1(n_532), .B2(n_630), .C(n_792), .Y(n_791) );
AOI222xp33_ASAP7_75t_L g808 ( .A1(n_22), .A2(n_33), .B1(n_230), .B2(n_382), .C1(n_386), .C2(n_483), .Y(n_808) );
XOR2x2_ASAP7_75t_L g486 ( .A(n_23), .B(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_24), .A2(n_71), .B1(n_398), .B2(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g640 ( .A(n_25), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_26), .A2(n_87), .B1(n_544), .B2(n_716), .Y(n_715) );
AO22x2_ASAP7_75t_L g285 ( .A1(n_27), .A2(n_77), .B1(n_277), .B2(n_282), .Y(n_285) );
INVx1_ASAP7_75t_L g786 ( .A(n_27), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_28), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_30), .A2(n_32), .B1(n_397), .B2(n_539), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_31), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_34), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_35), .A2(n_168), .B1(n_430), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_36), .A2(n_63), .B1(n_478), .B2(n_651), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_37), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_38), .A2(n_39), .B1(n_524), .B2(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g584 ( .A(n_40), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_41), .A2(n_188), .B1(n_308), .B2(n_530), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_42), .A2(n_53), .B1(n_630), .B2(n_631), .Y(n_629) );
AO22x2_ASAP7_75t_L g287 ( .A1(n_43), .A2(n_81), .B1(n_277), .B2(n_278), .Y(n_287) );
INVx1_ASAP7_75t_L g787 ( .A(n_43), .Y(n_787) );
INVx1_ASAP7_75t_L g573 ( .A(n_44), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_45), .A2(n_110), .B1(n_532), .B2(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_46), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_47), .A2(n_48), .B1(n_508), .B2(n_569), .Y(n_723) );
INVx1_ASAP7_75t_L g564 ( .A(n_49), .Y(n_564) );
INVx1_ASAP7_75t_L g572 ( .A(n_50), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_51), .A2(n_244), .B1(n_385), .B2(n_542), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_52), .A2(n_138), .B1(n_412), .B2(n_414), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_54), .B(n_524), .Y(n_653) );
INVx1_ASAP7_75t_L g446 ( .A(n_55), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_56), .B(n_349), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_57), .A2(n_213), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp5_ASAP7_75t_SL g626 ( .A1(n_58), .A2(n_239), .B1(n_469), .B2(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_59), .A2(n_111), .B1(n_409), .B2(n_410), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_61), .A2(n_180), .B1(n_414), .B2(n_721), .Y(n_720) );
XOR2x2_ASAP7_75t_L g706 ( .A(n_62), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_64), .B(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_65), .A2(n_82), .B1(n_403), .B2(n_405), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_66), .A2(n_187), .B1(n_272), .B2(n_440), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_67), .A2(n_232), .B1(n_494), .B2(n_502), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_70), .A2(n_169), .B1(n_438), .B2(n_633), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_72), .A2(n_144), .B1(n_403), .B2(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_73), .A2(n_92), .B1(n_410), .B2(n_465), .Y(n_464) );
AO22x1_ASAP7_75t_L g450 ( .A1(n_74), .A2(n_451), .B1(n_452), .B2(n_484), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_74), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_75), .A2(n_142), .B1(n_350), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_76), .A2(n_236), .B1(n_475), .B2(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_78), .A2(n_163), .B1(n_401), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_79), .A2(n_135), .B1(n_415), .B2(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_80), .A2(n_83), .B1(n_481), .B2(n_575), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_84), .A2(n_186), .B1(n_301), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_85), .A2(n_194), .B1(n_413), .B2(n_538), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_86), .Y(n_762) );
INVx1_ASAP7_75t_L g262 ( .A(n_88), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_89), .B(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_90), .A2(n_125), .B1(n_608), .B2(n_609), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_91), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_93), .A2(n_170), .B1(n_539), .B2(n_606), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_94), .Y(n_596) );
INVx1_ASAP7_75t_L g259 ( .A(n_95), .Y(n_259) );
INVx1_ASAP7_75t_L g643 ( .A(n_96), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_97), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_98), .A2(n_166), .B1(n_322), .B2(n_515), .Y(n_763) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_99), .A2(n_241), .B1(n_606), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_100), .A2(n_214), .B1(n_415), .B2(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_101), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_102), .A2(n_175), .B1(n_506), .B2(n_507), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_103), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_104), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_105), .A2(n_134), .B1(n_242), .B2(n_342), .C1(n_382), .C2(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_106), .B(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_108), .A2(n_151), .B1(n_386), .B2(n_430), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_109), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_112), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_113), .A2(n_118), .B1(n_386), .B2(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_114), .A2(n_162), .B1(n_469), .B2(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g820 ( .A(n_115), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_115), .A2(n_790), .B1(n_810), .B2(n_820), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_116), .A2(n_191), .B1(n_318), .B2(n_322), .Y(n_317) );
INVx1_ASAP7_75t_L g807 ( .A(n_117), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_119), .A2(n_249), .B1(n_538), .B2(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g555 ( .A(n_120), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_121), .A2(n_229), .B1(n_318), .B2(n_469), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_122), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_123), .A2(n_158), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_124), .A2(n_155), .B1(n_519), .B2(n_721), .Y(n_729) );
INVx1_ASAP7_75t_L g799 ( .A(n_126), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_127), .A2(n_152), .B1(n_468), .B2(n_469), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_128), .A2(n_228), .B1(n_501), .B2(n_502), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_129), .A2(n_179), .B1(n_510), .B2(n_512), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_130), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g738 ( .A1(n_131), .A2(n_160), .B1(n_193), .B2(n_338), .C1(n_342), .C2(n_483), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_132), .Y(n_288) );
INVx1_ASAP7_75t_L g793 ( .A(n_136), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_137), .Y(n_310) );
INVx2_ASAP7_75t_L g263 ( .A(n_139), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_140), .A2(n_221), .B1(n_350), .B2(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_141), .A2(n_254), .B1(n_507), .B2(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_143), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_145), .Y(n_332) );
INVx1_ASAP7_75t_L g801 ( .A(n_146), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_147), .A2(n_222), .B1(n_651), .B2(n_716), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_148), .A2(n_201), .B1(n_405), .B2(n_515), .Y(n_514) );
AND2x6_ASAP7_75t_L g258 ( .A(n_149), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_149), .Y(n_780) );
AO22x2_ASAP7_75t_L g276 ( .A1(n_150), .A2(n_209), .B1(n_277), .B2(n_278), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_153), .A2(n_206), .B1(n_472), .B2(n_475), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_154), .Y(n_327) );
INVx1_ASAP7_75t_L g664 ( .A(n_156), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_157), .A2(n_208), .B1(n_291), .B2(n_445), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_161), .A2(n_790), .B1(n_809), .B2(n_810), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_161), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_164), .A2(n_247), .B1(n_457), .B2(n_462), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_165), .A2(n_215), .B1(n_307), .B2(n_538), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_171), .A2(n_198), .B1(n_409), .B2(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_172), .A2(n_203), .B1(n_532), .B2(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_173), .B(n_525), .Y(n_654) );
AO22x2_ASAP7_75t_L g281 ( .A1(n_174), .A2(n_223), .B1(n_277), .B2(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_176), .B(n_636), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_177), .Y(n_391) );
XOR2x2_ASAP7_75t_L g725 ( .A(n_178), .B(n_726), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_181), .A2(n_740), .B1(n_769), .B2(n_770), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_181), .Y(n_769) );
INVx1_ASAP7_75t_L g582 ( .A(n_182), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_183), .Y(n_392) );
INVx1_ASAP7_75t_L g434 ( .A(n_184), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_185), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_189), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_192), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_195), .Y(n_294) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_196), .A2(n_250), .B1(n_342), .B2(n_479), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_197), .Y(n_757) );
INVx1_ASAP7_75t_L g558 ( .A(n_199), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_200), .A2(n_246), .B1(n_461), .B2(n_608), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_205), .A2(n_218), .B1(n_478), .B2(n_481), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_207), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_209), .B(n_785), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_210), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_211), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_212), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_216), .A2(n_225), .B1(n_405), .B2(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_217), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_220), .Y(n_750) );
INVx1_ASAP7_75t_L g783 ( .A(n_223), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_224), .A2(n_251), .B1(n_636), .B2(n_732), .Y(n_731) );
OA22x2_ASAP7_75t_L g669 ( .A1(n_226), .A2(n_670), .B1(n_671), .B2(n_693), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_226), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_231), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_233), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_234), .B(n_472), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_235), .A2(n_589), .B1(n_615), .B2(n_616), .Y(n_588) );
INVx1_ASAP7_75t_L g615 ( .A(n_235), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_237), .Y(n_376) );
INVx1_ASAP7_75t_L g277 ( .A(n_238), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_238), .Y(n_279) );
AOI211xp5_ASAP7_75t_L g255 ( .A1(n_240), .A2(n_256), .B(n_264), .C(n_788), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_243), .B(n_350), .Y(n_598) );
INVx1_ASAP7_75t_L g567 ( .A(n_245), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_248), .A2(n_268), .B1(n_366), .B2(n_367), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_248), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_252), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_253), .Y(n_424) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_258), .B(n_260), .Y(n_257) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_259), .Y(n_779) );
OA21x2_ASAP7_75t_L g818 ( .A1(n_260), .A2(n_778), .B(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_547), .B1(n_773), .B2(n_774), .C(n_775), .Y(n_264) );
INVx1_ASAP7_75t_L g773 ( .A(n_265), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_368), .B1(n_545), .B2(n_546), .Y(n_265) );
INVx2_ASAP7_75t_L g545 ( .A(n_266), .Y(n_545) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g367 ( .A(n_268), .Y(n_367) );
AND2x2_ASAP7_75t_SL g268 ( .A(n_269), .B(n_325), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_305), .Y(n_269) );
OAI221xp5_ASAP7_75t_SL g270 ( .A1(n_271), .A2(n_288), .B1(n_289), .B2(n_294), .C(n_295), .Y(n_270) );
OAI221xp5_ASAP7_75t_SL g554 ( .A1(n_271), .A2(n_555), .B1(n_556), .B2(n_558), .C(n_559), .Y(n_554) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx3_ASAP7_75t_L g409 ( .A(n_272), .Y(n_409) );
BUFx3_ASAP7_75t_L g612 ( .A(n_272), .Y(n_612) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_272), .Y(n_630) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_SL g438 ( .A(n_273), .Y(n_438) );
INVx2_ASAP7_75t_L g511 ( .A(n_273), .Y(n_511) );
BUFx2_ASAP7_75t_SL g719 ( .A(n_273), .Y(n_719) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_283), .Y(n_273) );
AND2x6_ASAP7_75t_L g298 ( .A(n_274), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g308 ( .A(n_274), .B(n_309), .Y(n_308) );
AND2x6_ASAP7_75t_L g338 ( .A(n_274), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_280), .Y(n_274) );
AND2x2_ASAP7_75t_L g293 ( .A(n_275), .B(n_281), .Y(n_293) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_276), .B(n_281), .Y(n_304) );
AND2x2_ASAP7_75t_L g314 ( .A(n_276), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g346 ( .A(n_276), .B(n_285), .Y(n_346) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g282 ( .A(n_279), .Y(n_282) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g315 ( .A(n_281), .Y(n_315) );
INVx1_ASAP7_75t_L g345 ( .A(n_281), .Y(n_345) );
AND2x4_ASAP7_75t_L g292 ( .A(n_283), .B(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g302 ( .A(n_283), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_283), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g399 ( .A(n_283), .B(n_314), .Y(n_399) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
OR2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_287), .Y(n_300) );
AND2x2_ASAP7_75t_L g309 ( .A(n_284), .B(n_287), .Y(n_309) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g339 ( .A(n_285), .B(n_287), .Y(n_339) );
AND2x2_ASAP7_75t_L g344 ( .A(n_286), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g358 ( .A(n_286), .Y(n_358) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g410 ( .A(n_292), .Y(n_410) );
BUFx3_ASAP7_75t_L g518 ( .A(n_292), .Y(n_518) );
INVx2_ASAP7_75t_L g533 ( .A(n_292), .Y(n_533) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_292), .Y(n_557) );
INVx1_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_293), .B(n_309), .Y(n_335) );
AND2x4_ASAP7_75t_L g474 ( .A(n_293), .B(n_299), .Y(n_474) );
AND2x6_ASAP7_75t_L g476 ( .A(n_293), .B(n_309), .Y(n_476) );
INVx4_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx4_ASAP7_75t_L g538 ( .A(n_297), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g563 ( .A1(n_297), .A2(n_564), .B1(n_565), .B2(n_567), .C(n_568), .Y(n_563) );
INVx2_ASAP7_75t_SL g608 ( .A(n_297), .Y(n_608) );
INVx3_ASAP7_75t_L g689 ( .A(n_297), .Y(n_689) );
INVx11_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx11_ASAP7_75t_L g404 ( .A(n_298), .Y(n_404) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g330 ( .A(n_300), .B(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g401 ( .A(n_302), .Y(n_401) );
BUFx2_ASAP7_75t_L g445 ( .A(n_302), .Y(n_445) );
BUFx3_ASAP7_75t_L g462 ( .A(n_302), .Y(n_462) );
BUFx3_ASAP7_75t_L g512 ( .A(n_302), .Y(n_512) );
INVx1_ASAP7_75t_L g535 ( .A(n_302), .Y(n_535) );
BUFx2_ASAP7_75t_SL g569 ( .A(n_302), .Y(n_569) );
BUFx3_ASAP7_75t_L g606 ( .A(n_302), .Y(n_606) );
AND2x2_ASAP7_75t_L g660 ( .A(n_303), .B(n_358), .Y(n_660) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x6_ASAP7_75t_L g323 ( .A(n_304), .B(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_310), .B1(n_311), .B2(n_316), .C(n_317), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx6_ASAP7_75t_L g406 ( .A(n_308), .Y(n_406) );
BUFx3_ASAP7_75t_L g461 ( .A(n_308), .Y(n_461) );
BUFx3_ASAP7_75t_L g539 ( .A(n_308), .Y(n_539) );
AND2x2_ASAP7_75t_L g321 ( .A(n_309), .B(n_314), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_309), .B(n_314), .Y(n_795) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g800 ( .A(n_312), .Y(n_800) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx5_ASAP7_75t_L g413 ( .A(n_320), .Y(n_413) );
INVx2_ASAP7_75t_L g440 ( .A(n_320), .Y(n_440) );
INVx3_ASAP7_75t_L g468 ( .A(n_320), .Y(n_468) );
BUFx3_ASAP7_75t_L g516 ( .A(n_320), .Y(n_516) );
INVx4_ASAP7_75t_L g562 ( .A(n_320), .Y(n_562) );
INVx8_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx6_ASAP7_75t_SL g415 ( .A(n_323), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_323), .A2(n_793), .B1(n_794), .B2(n_796), .Y(n_792) );
INVx1_ASAP7_75t_L g480 ( .A(n_324), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_336), .C(n_353), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_332), .B2(n_333), .Y(n_326) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g571 ( .A(n_329), .Y(n_571) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
BUFx3_ASAP7_75t_L g423 ( .A(n_330), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_333), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_333), .A2(n_571), .B1(n_572), .B2(n_573), .C(n_574), .Y(n_570) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g379 ( .A(n_334), .Y(n_379) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g747 ( .A(n_335), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B1(n_341), .B2(n_347), .C(n_348), .Y(n_336) );
OAI21xp5_ASAP7_75t_SL g489 ( .A1(n_337), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
BUFx3_ASAP7_75t_L g428 ( .A(n_338), .Y(n_428) );
INVx4_ASAP7_75t_L g583 ( .A(n_338), .Y(n_583) );
INVx2_ASAP7_75t_L g648 ( .A(n_338), .Y(n_648) );
INVx1_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
AND2x4_ASAP7_75t_L g481 ( .A(n_339), .B(n_365), .Y(n_481) );
OAI221xp5_ASAP7_75t_SL g594 ( .A1(n_341), .A2(n_595), .B1(n_596), .B2(n_597), .C(n_598), .Y(n_594) );
OAI222xp33_ASAP7_75t_L g673 ( .A1(n_341), .A2(n_674), .B1(n_676), .B2(n_677), .C1(n_678), .C2(n_679), .Y(n_673) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g749 ( .A(n_342), .Y(n_749) );
BUFx4f_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_343), .Y(n_386) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_343), .Y(n_501) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_343), .Y(n_581) );
BUFx2_ASAP7_75t_L g642 ( .A(n_343), .Y(n_642) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g352 ( .A(n_345), .Y(n_352) );
AND2x4_ASAP7_75t_L g351 ( .A(n_346), .B(n_352), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_346), .B(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g479 ( .A(n_346), .B(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g753 ( .A(n_350), .Y(n_753) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_351), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_359), .B2(n_360), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_355), .A2(n_360), .B1(n_756), .B2(n_757), .Y(n_755) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx3_ASAP7_75t_SL g601 ( .A(n_356), .Y(n_601) );
INVx4_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_357), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_390) );
BUFx3_ASAP7_75t_L g433 ( .A(n_357), .Y(n_433) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g393 ( .A(n_362), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_362), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_362), .A2(n_433), .B1(n_806), .B2(n_807), .Y(n_805) );
OR2x6_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g546 ( .A(n_368), .Y(n_546) );
XNOR2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_448), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_418), .B2(n_447), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_394), .Y(n_373) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_380), .C(n_390), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_378), .B2(n_379), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_377), .A2(n_379), .B1(n_592), .B2(n_593), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_377), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B1(n_384), .B2(n_387), .C(n_388), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_381), .A2(n_710), .B(n_711), .Y(n_709) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g751 ( .A(n_382), .Y(n_751) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g678 ( .A(n_389), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_393), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_407), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_402), .Y(n_395) );
BUFx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx3_ASAP7_75t_L g457 ( .A(n_399), .Y(n_457) );
BUFx3_ASAP7_75t_L g508 ( .A(n_399), .Y(n_508) );
BUFx3_ASAP7_75t_L g530 ( .A(n_399), .Y(n_530) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx4_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_404), .Y(n_466) );
INVx2_ASAP7_75t_SL g506 ( .A(n_404), .Y(n_506) );
INVx2_ASAP7_75t_L g631 ( .A(n_404), .Y(n_631) );
INVx1_ASAP7_75t_L g737 ( .A(n_404), .Y(n_737) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
INVx2_ASAP7_75t_L g566 ( .A(n_406), .Y(n_566) );
INVx2_ASAP7_75t_L g609 ( .A(n_406), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g692 ( .A(n_410), .Y(n_692) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_413), .Y(n_721) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g469 ( .A(n_415), .Y(n_469) );
BUFx2_ASAP7_75t_L g519 ( .A(n_415), .Y(n_519) );
INVx2_ASAP7_75t_SL g447 ( .A(n_418), .Y(n_447) );
XOR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_446), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_435), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_425), .C(n_431), .Y(n_420) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B(n_429), .Y(n_425) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx4f_ASAP7_75t_SL g483 ( .A(n_430), .Y(n_483) );
INVx2_ASAP7_75t_L g543 ( .A(n_430), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_441), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g760 ( .A(n_438), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
XNOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_485), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
NAND4xp75_ASAP7_75t_SL g452 ( .A(n_453), .B(n_463), .C(n_470), .D(n_482), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_458), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_471), .B(n_477), .Y(n_470) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_472), .Y(n_497) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_472), .Y(n_732) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g524 ( .A(n_473), .Y(n_524) );
INVx2_ASAP7_75t_L g683 ( .A(n_473), .Y(n_683) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g499 ( .A(n_476), .Y(n_499) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_476), .Y(n_525) );
INVx1_ASAP7_75t_SL g637 ( .A(n_476), .Y(n_637) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g502 ( .A(n_479), .Y(n_502) );
BUFx3_ASAP7_75t_L g527 ( .A(n_479), .Y(n_527) );
INVx1_ASAP7_75t_L g576 ( .A(n_479), .Y(n_576) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_481), .Y(n_494) );
BUFx2_ASAP7_75t_SL g544 ( .A(n_481), .Y(n_544) );
BUFx2_ASAP7_75t_SL g651 ( .A(n_481), .Y(n_651) );
INVx1_ASAP7_75t_L g585 ( .A(n_483), .Y(n_585) );
XOR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_520), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_488), .B(n_503), .Y(n_487) );
NOR2xp33_ASAP7_75t_SL g488 ( .A(n_489), .B(n_495), .Y(n_488) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .C(n_500), .Y(n_495) );
NOR2x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
BUFx4f_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g768 ( .A(n_508), .Y(n_768) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_518), .Y(n_613) );
NAND4xp75_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .C(n_536), .D(n_541), .Y(n_521) );
AND2x2_ASAP7_75t_SL g522 ( .A(n_523), .B(n_526), .Y(n_522) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g774 ( .A(n_547), .Y(n_774) );
AOI22xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_700), .B1(n_701), .B2(n_772), .Y(n_547) );
INVx1_ASAP7_75t_L g772 ( .A(n_548), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_618), .B1(n_619), .B2(n_699), .Y(n_548) );
INVx1_ASAP7_75t_L g699 ( .A(n_549), .Y(n_699) );
OAI22xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_551), .B1(n_588), .B2(n_617), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g587 ( .A(n_553), .Y(n_587) );
OR4x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_563), .C(n_570), .D(n_577), .Y(n_553) );
INVx4_ASAP7_75t_L g633 ( .A(n_556), .Y(n_633) );
OAI221xp5_ASAP7_75t_SL g759 ( .A1(n_556), .A2(n_760), .B1(n_761), .B2(n_762), .C(n_763), .Y(n_759) );
INVx4_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_562), .Y(n_627) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_SL g802 ( .A(n_569), .Y(n_802) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g716 ( .A(n_576), .Y(n_716) );
OAI222xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_582), .B1(n_583), .B2(n_584), .C1(n_585), .C2(n_586), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx4_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g595 ( .A(n_583), .Y(n_595) );
INVx4_ASAP7_75t_L g675 ( .A(n_583), .Y(n_675) );
INVx1_ASAP7_75t_L g617 ( .A(n_588), .Y(n_617) );
INVx2_ASAP7_75t_L g616 ( .A(n_589), .Y(n_616) );
AND2x2_ASAP7_75t_SL g589 ( .A(n_590), .B(n_603), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .C(n_599), .Y(n_590) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_595), .A2(n_640), .B(n_641), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_610), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_621), .B1(n_667), .B2(n_668), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_644), .B1(n_665), .B2(n_666), .Y(n_621) );
INVx2_ASAP7_75t_SL g665 ( .A(n_622), .Y(n_665) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_643), .Y(n_622) );
NOR4xp75_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .C(n_634), .D(n_639), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_635), .B(n_638), .Y(n_634) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g804 ( .A(n_637), .Y(n_804) );
INVx1_ASAP7_75t_L g666 ( .A(n_644), .Y(n_666) );
INVx2_ASAP7_75t_L g695 ( .A(n_644), .Y(n_695) );
XOR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_664), .Y(n_644) );
NAND2x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_656), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_652), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_649), .B(n_650), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .C(n_655), .Y(n_652) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_661), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g698 ( .A(n_666), .Y(n_698) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_694), .B1(n_696), .B2(n_697), .Y(n_668) );
INVx1_ASAP7_75t_L g696 ( .A(n_669), .Y(n_696) );
INVx2_ASAP7_75t_L g693 ( .A(n_671), .Y(n_693) );
NAND3x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_684), .C(n_687), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_680), .Y(n_672) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_739), .B2(n_771), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
XNOR2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_725), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_717), .C(n_722), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_712), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .C(n_715), .Y(n_712) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
NAND4xp75_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .C(n_734), .D(n_738), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
AND2x2_ASAP7_75t_SL g730 ( .A(n_731), .B(n_733), .Y(n_730) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g771 ( .A(n_739), .Y(n_771) );
INVx1_ASAP7_75t_L g770 ( .A(n_740), .Y(n_770) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_758), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_748), .C(n_755), .Y(n_741) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI222xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_752), .C1(n_753), .C2(n_754), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_764), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
NOR2x1_ASAP7_75t_L g776 ( .A(n_777), .B(n_781), .Y(n_776) );
OR2x2_ASAP7_75t_SL g826 ( .A(n_777), .B(n_782), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_778), .Y(n_812) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_779), .B(n_815), .Y(n_819) );
CKINVDCx16_ASAP7_75t_R g815 ( .A(n_780), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
OAI322xp33_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_811), .A3(n_813), .B1(n_816), .B2(n_820), .C1(n_821), .C2(n_825), .Y(n_788) );
INVx1_ASAP7_75t_L g810 ( .A(n_790), .Y(n_810) );
AND4x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_797), .C(n_803), .D(n_808), .Y(n_790) );
BUFx2_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_798) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
CKINVDCx14_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
endmodule