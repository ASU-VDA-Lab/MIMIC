module fake_jpeg_14301_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_22),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_44),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_22),
.B(n_6),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_64),
.Y(n_90)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_6),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_70),
.Y(n_92)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_73),
.Y(n_91)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx9p33_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_29),
.B1(n_72),
.B2(n_71),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_78),
.A2(n_121),
.B1(n_92),
.B2(n_83),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_88),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_40),
.B1(n_18),
.B2(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_116),
.B1(n_118),
.B2(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_99),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_39),
.B1(n_19),
.B2(n_20),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_104),
.B1(n_120),
.B2(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_74),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_19),
.B1(n_34),
.B2(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_24),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_30),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_52),
.A2(n_16),
.B1(n_23),
.B2(n_30),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_119),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_16),
.B1(n_37),
.B2(n_27),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_7),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_56),
.A2(n_34),
.B1(n_37),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_34),
.B1(n_6),
.B2(n_7),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_61),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_3),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_147),
.C(n_149),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_68),
.B(n_42),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_161),
.B(n_147),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_128)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_128),
.A2(n_136),
.B1(n_140),
.B2(n_153),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_129),
.A2(n_163),
.B1(n_166),
.B2(n_126),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_8),
.B1(n_11),
.B2(n_86),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_134),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_86),
.A2(n_114),
.B1(n_77),
.B2(n_115),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_77),
.B1(n_115),
.B2(n_93),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_156),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_88),
.B1(n_97),
.B2(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_138),
.B1(n_164),
.B2(n_159),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_96),
.B1(n_110),
.B2(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

AO22x1_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_123),
.B1(n_85),
.B2(n_110),
.Y(n_140)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_154),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_91),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_108),
.C(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_76),
.A3(n_106),
.B1(n_94),
.B2(n_105),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_140),
.A3(n_127),
.B1(n_136),
.B2(n_129),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_105),
.A2(n_79),
.B(n_122),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_103),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_165),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_79),
.A2(n_122),
.B(n_80),
.C(n_84),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_161),
.B(n_167),
.Y(n_171)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_101),
.A2(n_83),
.B1(n_88),
.B2(n_93),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_101),
.A2(n_121),
.B1(n_47),
.B2(n_45),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_80),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_80),
.A2(n_87),
.B1(n_74),
.B2(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_152),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_184),
.B(n_194),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_190),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_128),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_128),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_142),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_149),
.B(n_141),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_155),
.B1(n_145),
.B2(n_148),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_130),
.A2(n_137),
.B(n_140),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_170),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_136),
.B(n_165),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_136),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_128),
.B(n_162),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_210),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_199),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_204),
.A2(n_224),
.B1(n_172),
.B2(n_177),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_220),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_171),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_185),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_222),
.C(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_184),
.B1(n_201),
.B2(n_187),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_229),
.B(n_195),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_182),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_225),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_173),
.B1(n_179),
.B2(n_171),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_176),
.B(n_170),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_177),
.Y(n_247)
);

AO22x1_ASAP7_75t_SL g229 ( 
.A1(n_179),
.A2(n_174),
.B1(n_175),
.B2(n_186),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_246),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_235),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_174),
.B(n_195),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_248),
.B(n_216),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_242),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_186),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_178),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_219),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_202),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_262),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_234),
.B(n_230),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_203),
.B1(n_204),
.B2(n_207),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_259),
.B1(n_261),
.B2(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_204),
.B1(n_213),
.B2(n_205),
.Y(n_259)
);

AOI211xp5_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_206),
.B(n_229),
.C(n_215),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_220),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_240),
.C(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_225),
.B1(n_206),
.B2(n_229),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_278),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_235),
.B1(n_248),
.B2(n_230),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_282),
.B1(n_244),
.B2(n_242),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_253),
.B(n_265),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_233),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_280),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_247),
.B1(n_229),
.B2(n_241),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_269),
.B1(n_267),
.B2(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_250),
.B1(n_240),
.B2(n_243),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_275),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_261),
.C(n_250),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_212),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_277),
.B(n_276),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_211),
.B(n_238),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_279),
.B(n_274),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_256),
.C(n_252),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_289),
.C(n_272),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_256),
.C(n_262),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_238),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_226),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_223),
.B1(n_218),
.B2(n_212),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_289),
.C(n_287),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_272),
.B1(n_274),
.B2(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_300),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_301),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_296),
.Y(n_307)
);

OAI221xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_291),
.B1(n_285),
.B2(n_290),
.C(n_293),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_295),
.B(n_299),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_294),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_305),
.B1(n_300),
.B2(n_286),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_311),
.B(n_286),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_306),
.CI(n_310),
.CON(n_313),
.SN(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_306),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_313),
.Y(n_315)
);


endmodule