module real_jpeg_11330_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_259;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_1),
.A2(n_28),
.B1(n_58),
.B2(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_1),
.A2(n_28),
.B1(n_53),
.B2(n_62),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_34),
.B1(n_53),
.B2(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_26),
.B1(n_29),
.B2(n_41),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_53),
.B1(n_62),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_5),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_102),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_5),
.A2(n_26),
.B1(n_29),
.B2(n_102),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_102),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_11),
.A2(n_53),
.B1(n_62),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_11),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_151),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_151),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_11),
.A2(n_26),
.B1(n_29),
.B2(n_151),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_13),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_13),
.A2(n_55),
.B(n_59),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_13),
.A2(n_53),
.B1(n_62),
.B2(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_13),
.B(n_66),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_13),
.A2(n_37),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_13),
.B(n_37),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_13),
.A2(n_82),
.B1(n_83),
.B2(n_231),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_14),
.A2(n_26),
.B1(n_29),
.B2(n_63),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_63),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_15),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_15),
.A2(n_26),
.B1(n_29),
.B2(n_48),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_15),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_19),
.B(n_106),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_79),
.C(n_90),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_20),
.A2(n_21),
.B1(n_79),
.B2(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_22),
.B(n_50),
.C(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_23),
.B(n_35),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_24),
.A2(n_83),
.B(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_26),
.A2(n_29),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_26),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_222)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_29),
.B(n_46),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_29),
.B(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_30),
.A2(n_31),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_31),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_32),
.A2(n_82),
.B(n_215),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_36),
.A2(n_45),
.B(n_96),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_43),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_38),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_37),
.B(n_70),
.Y(n_259)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_38),
.A2(n_75),
.B1(n_254),
.B2(n_259),
.Y(n_258)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_47),
.B(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_42),
.A2(n_45),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_42),
.A2(n_45),
.B1(n_221),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_42),
.A2(n_45),
.B1(n_244),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_42),
.A2(n_125),
.B(n_252),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_44),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_45),
.B(n_155),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_67),
.B2(n_78),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_61),
.B(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_57),
.B1(n_61),
.B2(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_52),
.A2(n_57),
.B1(n_101),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_52),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_53),
.A2(n_54),
.B(n_155),
.C(n_156),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.C(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_70),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g254 ( 
.A(n_59),
.B(n_155),
.CON(n_254),
.SN(n_254)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_66),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_73),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_77),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_68),
.A2(n_145),
.B1(n_146),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_68),
.A2(n_145),
.B1(n_176),
.B2(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_68),
.B(n_155),
.Y(n_242)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_74),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_69),
.B(n_104),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_69),
.A2(n_74),
.B1(n_199),
.B2(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_74),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_79),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_81),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_85),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_82),
.A2(n_83),
.B1(n_213),
.B2(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_82),
.A2(n_84),
.B(n_94),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_83),
.B(n_155),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_87),
.A2(n_98),
.B(n_127),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.C(n_103),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_95),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_130),
.B2(n_131),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_119),
.B1(n_120),
.B2(n_129),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B(n_128),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_130),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_162),
.B(n_285),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_159),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_136),
.B(n_159),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_141),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_140),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_141),
.A2(n_142),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.C(n_152),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B(n_147),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_204),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_185),
.B(n_203),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_205),
.C(n_284),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_182),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_182),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_181),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_175),
.B1(n_181),
.B2(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_186),
.B(n_188),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_189),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_192),
.A2(n_194),
.B1(n_195),
.B2(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_192),
.Y(n_282)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.C(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_196),
.A2(n_197),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_200),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_278),
.B(n_283),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_263),
.B(n_277),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_247),
.B(n_262),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_238),
.B(n_246),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_227),
.B(n_237),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_216),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_222),
.B2(n_226),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_226),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_222),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_232),
.B(n_236),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_248),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.CI(n_245),
.CON(n_241),
.SN(n_241)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_257),
.B2(n_261),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_256),
.C(n_261),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_257),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_260),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_271),
.B2(n_272),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_274),
.C(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_273),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);


endmodule