module fake_jpeg_87_n_543 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_150;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_46),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_51),
.Y(n_104)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_50),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_62),
.Y(n_114)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_19),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_12),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g99 ( 
.A(n_82),
.Y(n_99)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_87),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_26),
.B(n_13),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_95),
.B(n_22),
.Y(n_112)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_13),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_96),
.Y(n_118)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_101),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_19),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_42),
.B1(n_29),
.B2(n_34),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_102),
.A2(n_131),
.B1(n_145),
.B2(n_28),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_36),
.B1(n_42),
.B2(n_34),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_111),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_45),
.B(n_34),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_120),
.B(n_127),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_66),
.B(n_29),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_47),
.A2(n_42),
.B1(n_15),
.B2(n_29),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_36),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_135),
.B(n_139),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_36),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_15),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_158),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_15),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_42),
.B1(n_17),
.B2(n_16),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_82),
.B(n_16),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_86),
.B(n_38),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_93),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_53),
.B(n_16),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_20),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_17),
.B1(n_95),
.B2(n_38),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_161),
.A2(n_184),
.B1(n_197),
.B2(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_163),
.B(n_168),
.Y(n_227)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

BUFx4f_ASAP7_75t_SL g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_104),
.B(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_181),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_102),
.A2(n_88),
.B1(n_50),
.B2(n_55),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_193),
.B1(n_145),
.B2(n_39),
.Y(n_216)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_117),
.B(n_58),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_178),
.Y(n_231)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_100),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_192),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_17),
.B1(n_38),
.B2(n_39),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_107),
.B(n_21),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_146),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_189),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_136),
.C(n_152),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_134),
.A2(n_21),
.B(n_20),
.C(n_28),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_128),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_113),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_109),
.B(n_18),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_125),
.A2(n_17),
.B1(n_28),
.B2(n_39),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_109),
.B(n_18),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_0),
.Y(n_238)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_133),
.B1(n_56),
.B2(n_130),
.Y(n_240)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_78),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_116),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_212),
.B(n_215),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_170),
.B(n_128),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_216),
.A2(n_222),
.B1(n_204),
.B2(n_190),
.Y(n_274)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_188),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_195),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_133),
.B1(n_138),
.B2(n_147),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_196),
.B1(n_198),
.B2(n_174),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_167),
.A2(n_110),
.B1(n_147),
.B2(n_138),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_240),
.B1(n_201),
.B2(n_194),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_207),
.A3(n_213),
.B1(n_223),
.B2(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_260),
.Y(n_280)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_246),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_SL g247 ( 
.A1(n_208),
.A2(n_166),
.B(n_202),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_259),
.Y(n_299)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_167),
.B1(n_193),
.B2(n_199),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_253),
.B1(n_234),
.B2(n_218),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_202),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_250),
.B(n_255),
.Y(n_304)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_181),
.CI(n_183),
.CON(n_255),
.SN(n_255)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_230),
.B1(n_240),
.B2(n_176),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_166),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_258),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_162),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_262),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_165),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_212),
.A2(n_172),
.B(n_192),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_264),
.A2(n_236),
.B(n_233),
.Y(n_301)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_216),
.A2(n_160),
.B1(n_179),
.B2(n_205),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_274),
.B1(n_222),
.B2(n_210),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_224),
.B(n_208),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_224),
.B(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_218),
.B(n_204),
.CI(n_159),
.CON(n_270),
.SN(n_270)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_231),
.A3(n_236),
.B1(n_221),
.B2(n_220),
.Y(n_300)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_271),
.B(n_275),
.Y(n_298)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_L g337 ( 
.A1(n_276),
.A2(n_233),
.B(n_243),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_224),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_278),
.B(n_303),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_286),
.B1(n_267),
.B2(n_256),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_273),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_283),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_242),
.B(n_230),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_285),
.A2(n_288),
.B(n_301),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_264),
.B(n_260),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_290),
.A2(n_169),
.B1(n_251),
.B2(n_237),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_305),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_253),
.A2(n_231),
.B1(n_185),
.B2(n_110),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_307),
.B1(n_265),
.B2(n_210),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_261),
.B(n_220),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_221),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_249),
.B(n_214),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_248),
.C(n_244),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_259),
.A2(n_206),
.B1(n_164),
.B2(n_130),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_298),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_309),
.A2(n_311),
.B1(n_312),
.B2(n_325),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_285),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_310),
.B(n_336),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_298),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_259),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_313),
.B(n_329),
.C(n_299),
.Y(n_357)
);

XNOR2x2_ASAP7_75t_SL g315 ( 
.A(n_278),
.B(n_292),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_318),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_320),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_319),
.B1(n_323),
.B2(n_326),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_270),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_291),
.B(n_289),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_282),
.A2(n_252),
.B1(n_246),
.B2(n_255),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_302),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_305),
.A2(n_270),
.B1(n_262),
.B2(n_266),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_292),
.A2(n_273),
.B1(n_275),
.B2(n_271),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_327),
.A2(n_307),
.B1(n_290),
.B2(n_294),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_214),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_269),
.B1(n_254),
.B2(n_263),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_330),
.A2(n_334),
.B1(n_283),
.B2(n_279),
.Y(n_366)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

AO22x1_ASAP7_75t_SL g335 ( 
.A1(n_296),
.A2(n_251),
.B1(n_237),
.B2(n_241),
.Y(n_335)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_276),
.Y(n_355)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_237),
.Y(n_340)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_340),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_229),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_342),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_289),
.B(n_229),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_330),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_347),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_324),
.B(n_338),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_346),
.B(n_349),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_348),
.A2(n_366),
.B1(n_321),
.B2(n_333),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_324),
.B(n_280),
.Y(n_349)
);

OAI22x1_ASAP7_75t_L g351 ( 
.A1(n_310),
.A2(n_299),
.B1(n_300),
.B2(n_294),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_351),
.A2(n_375),
.B1(n_326),
.B2(n_327),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_331),
.A2(n_299),
.B(n_304),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_363),
.B(n_297),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_315),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_340),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_361),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_309),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_331),
.A2(n_277),
.B(n_308),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_279),
.Y(n_364)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_339),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_373),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_329),
.C(n_313),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_343),
.C(n_357),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_328),
.A2(n_308),
.B(n_287),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_371),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_287),
.Y(n_372)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_372),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_322),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_374),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_323),
.A2(n_328),
.B1(n_338),
.B2(n_317),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_379),
.B1(n_387),
.B2(n_395),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_344),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_392),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_390),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_354),
.A2(n_319),
.B1(n_315),
.B2(n_335),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_382),
.A2(n_384),
.B1(n_404),
.B2(n_356),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_345),
.A2(n_335),
.B1(n_336),
.B2(n_325),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_388),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_375),
.A2(n_297),
.B1(n_295),
.B2(n_302),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_295),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_239),
.C(n_243),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_393),
.C(n_407),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_228),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_347),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_228),
.C(n_241),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_367),
.A2(n_241),
.B1(n_203),
.B2(n_191),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_367),
.A2(n_177),
.B1(n_173),
.B2(n_182),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_396),
.A2(n_405),
.B1(n_391),
.B2(n_377),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_364),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_10),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_180),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_99),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_124),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_401),
.Y(n_416)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_403),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_361),
.A2(n_348),
.B1(n_369),
.B2(n_356),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_352),
.Y(n_405)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_156),
.C(n_150),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_409),
.A2(n_415),
.B1(n_394),
.B2(n_402),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_398),
.Y(n_411)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_SL g412 ( 
.A1(n_382),
.A2(n_371),
.B(n_369),
.C(n_363),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_412),
.A2(n_84),
.B(n_22),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_406),
.A2(n_350),
.B1(n_362),
.B2(n_373),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_423),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_417),
.A2(n_419),
.B1(n_422),
.B2(n_429),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_379),
.A2(n_374),
.B1(n_368),
.B2(n_360),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_388),
.B(n_360),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_420),
.B(n_123),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_387),
.A2(n_368),
.B1(n_359),
.B2(n_352),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_359),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_399),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_430),
.Y(n_454)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_426),
.Y(n_450)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_404),
.Y(n_428)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_385),
.A2(n_57),
.B1(n_63),
.B2(n_94),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_434),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_433),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_389),
.B(n_149),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_396),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_381),
.C(n_393),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_441),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_418),
.B(n_407),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_438),
.B(n_452),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_408),
.B(n_384),
.C(n_397),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_414),
.A2(n_395),
.B1(n_397),
.B2(n_90),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_442),
.A2(n_410),
.B1(n_416),
.B2(n_432),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_431),
.C(n_427),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_444),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_156),
.C(n_150),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_445),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g464 ( 
.A1(n_446),
.A2(n_412),
.B(n_43),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_123),
.C(n_121),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_449),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_123),
.C(n_121),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_79),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_40),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_121),
.C(n_129),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_0),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_89),
.Y(n_458)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_458),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_453),
.A2(n_409),
.B1(n_410),
.B2(n_412),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_461),
.A2(n_463),
.B1(n_445),
.B2(n_456),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_464),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_412),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_476),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_429),
.C(n_89),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_468),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_78),
.C(n_41),
.Y(n_468)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_40),
.C(n_27),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_474),
.B(n_477),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_475),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_43),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_43),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_40),
.C(n_27),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_479),
.C(n_455),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_27),
.C(n_1),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_490),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_456),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_486),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_467),
.A2(n_440),
.B1(n_458),
.B2(n_460),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_485),
.A2(n_488),
.B1(n_480),
.B2(n_476),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_461),
.A2(n_439),
.B(n_450),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_487),
.A2(n_495),
.B(n_471),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_469),
.A2(n_447),
.B1(n_457),
.B2(n_449),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_473),
.A2(n_452),
.B1(n_13),
.B2(n_11),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_11),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_494),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_10),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_462),
.A2(n_9),
.B(n_1),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_9),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_496),
.B(n_497),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_9),
.Y(n_497)
);

AO21x1_ASAP7_75t_L g519 ( 
.A1(n_500),
.A2(n_509),
.B(n_510),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_486),
.B(n_468),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_501),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_478),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_502),
.B(n_511),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_507),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_474),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_504),
.B(n_505),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_479),
.C(n_471),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_0),
.Y(n_507)
);

AOI21xp33_ASAP7_75t_L g508 ( 
.A1(n_487),
.A2(n_2),
.B(n_3),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_508),
.A2(n_499),
.B(n_506),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_2),
.Y(n_511)
);

INVx6_ASAP7_75t_L g512 ( 
.A(n_488),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_513),
.B(n_493),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_481),
.B(n_2),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_514),
.A2(n_516),
.B(n_520),
.Y(n_532)
);

AOI21x1_ASAP7_75t_L g516 ( 
.A1(n_512),
.A2(n_491),
.B(n_483),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_519),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_482),
.B1(n_490),
.B2(n_5),
.Y(n_521)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_521),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_504),
.A2(n_3),
.B(n_4),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_524),
.A2(n_5),
.B(n_6),
.Y(n_527)
);

OA21x2_ASAP7_75t_SL g525 ( 
.A1(n_518),
.A2(n_507),
.B(n_6),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_525),
.B(n_527),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_522),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_8),
.C(n_532),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_5),
.C(n_6),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_530),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_521),
.A2(n_5),
.B(n_7),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_531),
.A2(n_515),
.B(n_7),
.Y(n_534)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_534),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_526),
.A2(n_7),
.B(n_8),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_537),
.C(n_529),
.Y(n_539)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_536),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_538),
.A2(n_539),
.B(n_533),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_540),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_8),
.Y(n_543)
);


endmodule