module fake_netlist_1_11063_n_665 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_665);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_665;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g86 ( .A(n_9), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_41), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_24), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_0), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_65), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_18), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_67), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_38), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_12), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_10), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_45), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_29), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_18), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_7), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_73), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_40), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_23), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_49), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_82), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_80), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_19), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_11), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_43), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_28), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_26), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_31), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_37), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_57), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_46), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_35), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_68), .Y(n_123) );
BUFx8_ASAP7_75t_SL g124 ( .A(n_39), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_110), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_115), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_115), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_115), .B(n_1), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_87), .A2(n_42), .B(n_83), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_88), .B(n_1), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_86), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_107), .B(n_2), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_99), .B(n_3), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_93), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_91), .B(n_48), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_88), .B(n_5), .Y(n_140) );
AOI22x1_ASAP7_75t_SL g141 ( .A1(n_101), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_90), .B(n_8), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_92), .B(n_10), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_90), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_115), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_98), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_105), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_86), .B(n_11), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_109), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_96), .B(n_12), .Y(n_154) );
INVxp33_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_138), .B(n_89), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_145), .B(n_112), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_130), .B(n_95), .Y(n_159) );
BUFx8_ASAP7_75t_SL g160 ( .A(n_130), .Y(n_160) );
NAND2xp33_ASAP7_75t_L g161 ( .A(n_138), .B(n_102), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_131), .B(n_103), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_133), .B(n_96), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
NOR3xp33_ASAP7_75t_L g166 ( .A(n_134), .B(n_100), .C(n_111), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_154), .A2(n_113), .B1(n_109), .B2(n_111), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_131), .B(n_108), .Y(n_168) );
BUFx10_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_133), .B(n_114), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_135), .B(n_116), .Y(n_171) );
INVx11_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_153), .B(n_113), .Y(n_173) );
AO22x2_ASAP7_75t_L g174 ( .A1(n_141), .A2(n_119), .B1(n_105), .B2(n_106), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_126), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_133), .B(n_117), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_139), .B(n_112), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_125), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_126), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_125), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_135), .B(n_104), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_153), .B(n_97), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_126), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_127), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_139), .B(n_97), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_140), .B(n_121), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_144), .B(n_148), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_140), .A2(n_97), .B1(n_123), .B2(n_118), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_125), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_154), .A2(n_97), .B1(n_123), .B2(n_118), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_179), .B(n_171), .Y(n_192) );
AOI22xp5_ASAP7_75t_SL g193 ( .A1(n_179), .A2(n_136), .B1(n_141), .B2(n_154), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_182), .B(n_183), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_155), .B(n_136), .Y(n_195) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_174), .A2(n_134), .B1(n_140), .B2(n_142), .Y(n_196) );
AOI22xp33_ASAP7_75t_SL g197 ( .A1(n_174), .A2(n_140), .B1(n_142), .B2(n_152), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_170), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_183), .B(n_144), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_173), .B(n_148), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_173), .B(n_152), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_176), .B(n_149), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_156), .A2(n_132), .B(n_149), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_170), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_170), .A2(n_142), .B1(n_138), .B2(n_151), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_178), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_169), .B(n_142), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_178), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_189), .A2(n_137), .B1(n_151), .B2(n_129), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_181), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_160), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_165), .B(n_132), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_176), .B(n_143), .Y(n_219) );
AND3x2_ASAP7_75t_SL g220 ( .A(n_174), .B(n_137), .C(n_138), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_176), .B(n_129), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_169), .B(n_122), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_170), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_176), .B(n_120), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_187), .B(n_94), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_187), .B(n_129), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_187), .B(n_129), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_158), .B(n_13), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_159), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_187), .B(n_167), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_170), .B(n_138), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_165), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_162), .B(n_117), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_170), .A2(n_138), .B1(n_128), .B2(n_97), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_190), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_163), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g238 ( .A(n_189), .B(n_106), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_186), .B(n_97), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_209), .A2(n_161), .B(n_165), .Y(n_240) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_232), .A2(n_188), .B(n_164), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_233), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_204), .A2(n_165), .B(n_164), .Y(n_243) );
NOR3xp33_ASAP7_75t_SL g244 ( .A(n_229), .B(n_168), .C(n_174), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_217), .B(n_164), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_202), .A2(n_164), .B(n_163), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_201), .B(n_170), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_195), .B(n_172), .Y(n_248) );
OAI22xp5_ASAP7_75t_SL g249 ( .A1(n_215), .A2(n_174), .B1(n_166), .B2(n_191), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_233), .Y(n_250) );
BUFx2_ASAP7_75t_SL g251 ( .A(n_205), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_205), .B(n_186), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_201), .B(n_177), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_195), .B(n_138), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_200), .B(n_163), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_221), .A2(n_184), .B(n_180), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_228), .Y(n_257) );
NOR2xp33_ASAP7_75t_SL g258 ( .A(n_205), .B(n_124), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_233), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_226), .A2(n_184), .B(n_180), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_233), .Y(n_261) );
NAND3xp33_ASAP7_75t_SL g262 ( .A(n_197), .B(n_114), .C(n_119), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_192), .B(n_172), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_196), .A2(n_121), .B1(n_132), .B2(n_180), .Y(n_264) );
OAI21xp33_ASAP7_75t_L g265 ( .A1(n_207), .A2(n_184), .B(n_175), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_193), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_219), .A2(n_175), .B(n_150), .C(n_146), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_194), .B(n_175), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_199), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_217), .B(n_147), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_211), .A2(n_146), .B(n_150), .C(n_132), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g272 ( .A1(n_230), .A2(n_146), .B(n_150), .C(n_132), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_225), .B(n_13), .Y(n_273) );
AO21x1_ASAP7_75t_L g274 ( .A1(n_218), .A2(n_147), .B(n_127), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_SL g275 ( .A1(n_234), .A2(n_185), .B(n_147), .C(n_127), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_205), .B(n_14), .Y(n_276) );
AO21x1_ASAP7_75t_L g277 ( .A1(n_218), .A2(n_147), .B(n_127), .Y(n_277) );
OR2x6_ASAP7_75t_SL g278 ( .A(n_220), .B(n_193), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_203), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_224), .B(n_15), .Y(n_280) );
AND2x6_ASAP7_75t_L g281 ( .A(n_198), .B(n_147), .Y(n_281) );
O2A1O1Ixp5_ASAP7_75t_L g282 ( .A1(n_222), .A2(n_185), .B(n_56), .C(n_59), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_227), .A2(n_185), .B(n_147), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_238), .A2(n_210), .B(n_206), .C(n_236), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_228), .B(n_15), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_206), .A2(n_185), .B(n_127), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_243), .A2(n_238), .B(n_237), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_249), .A2(n_223), .B1(n_198), .B2(n_214), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_281), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_279), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_276), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_269), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_257), .A2(n_239), .B(n_210), .C(n_236), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_248), .A2(n_223), .B1(n_198), .B2(n_214), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_SL g295 ( .A1(n_267), .A2(n_203), .B(n_216), .C(n_208), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_253), .B(n_239), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_262), .A2(n_216), .B(n_208), .C(n_231), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_247), .A2(n_214), .B1(n_223), .B2(n_213), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_255), .Y(n_299) );
AO31x2_ASAP7_75t_L g300 ( .A1(n_264), .A2(n_216), .A3(n_203), .B(n_231), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_276), .B(n_213), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_255), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_240), .A2(n_237), .B(n_212), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_266), .B(n_213), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_254), .A2(n_237), .B(n_212), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_285), .A2(n_231), .B(n_208), .C(n_212), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_254), .A2(n_218), .B(n_213), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_256), .A2(n_235), .B(n_220), .Y(n_308) );
AO32x2_ASAP7_75t_L g309 ( .A1(n_264), .A2(n_220), .A3(n_127), .B1(n_19), .B2(n_17), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_252), .B(n_217), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_273), .A2(n_217), .B1(n_17), .B2(n_16), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_252), .A2(n_263), .B1(n_280), .B2(n_245), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_268), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g314 ( .A1(n_284), .A2(n_217), .B(n_20), .C(n_21), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_16), .B1(n_185), .B2(n_25), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_242), .B(n_22), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_268), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_250), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_SL g320 ( .A1(n_275), .A2(n_27), .B(n_30), .C(n_32), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_246), .A2(n_185), .B(n_34), .C(n_36), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_271), .A2(n_33), .B(n_44), .C(n_47), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_313), .B(n_244), .Y(n_323) );
OAI221xp5_ASAP7_75t_L g324 ( .A1(n_292), .A2(n_258), .B1(n_261), .B2(n_265), .C(n_259), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
OAI21x1_ASAP7_75t_L g326 ( .A1(n_303), .A2(n_274), .B(n_277), .Y(n_326) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_317), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_302), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_295), .A2(n_272), .B(n_283), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_307), .A2(n_286), .B(n_270), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_301), .B(n_241), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_291), .A2(n_251), .B1(n_260), .B2(n_281), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_304), .B(n_281), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g335 ( .A1(n_293), .A2(n_311), .B(n_297), .C(n_308), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_300), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_319), .Y(n_337) );
AOI222xp33_ASAP7_75t_L g338 ( .A1(n_288), .A2(n_281), .B1(n_282), .B2(n_53), .C1(n_54), .C2(n_55), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_296), .B(n_84), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_312), .B(n_50), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_301), .B(n_51), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_287), .A2(n_60), .B(n_61), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_305), .A2(n_62), .B(n_63), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_311), .A2(n_64), .B(n_66), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_306), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_314), .A2(n_69), .B(n_70), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_315), .A2(n_71), .B1(n_72), .B2(n_74), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_328), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_327), .B(n_300), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_335), .A2(n_322), .B(n_321), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_328), .Y(n_355) );
AO21x2_ASAP7_75t_L g356 ( .A1(n_329), .A2(n_320), .B(n_309), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_336), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_331), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_331), .B(n_300), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_326), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_325), .B(n_316), .Y(n_361) );
AO21x2_ASAP7_75t_L g362 ( .A1(n_345), .A2(n_316), .B(n_298), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_344), .A2(n_294), .B1(n_318), .B2(n_289), .C(n_79), .Y(n_363) );
AOI21x1_ASAP7_75t_L g364 ( .A1(n_345), .A2(n_289), .B(n_318), .Y(n_364) );
AO21x2_ASAP7_75t_L g365 ( .A1(n_326), .A2(n_289), .B(n_318), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_325), .B(n_75), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_347), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_347), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_331), .B(n_76), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_327), .A2(n_77), .B1(n_81), .B2(n_323), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_349), .A2(n_344), .B(n_346), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_349), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_338), .B(n_332), .Y(n_373) );
OAI21xp5_ASAP7_75t_L g374 ( .A1(n_338), .A2(n_350), .B(n_340), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_323), .B(n_348), .Y(n_375) );
AOI21xp5_ASAP7_75t_SL g376 ( .A1(n_333), .A2(n_341), .B(n_339), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_334), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_367), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_359), .B(n_331), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_354), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_354), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_352), .B(n_337), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_367), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_359), .B(n_337), .Y(n_385) );
INVx5_ASAP7_75t_SL g386 ( .A(n_369), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_367), .Y(n_387) );
INVx5_ASAP7_75t_L g388 ( .A(n_369), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_354), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_368), .Y(n_390) );
NOR2x1_ASAP7_75t_SL g391 ( .A(n_355), .B(n_341), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_355), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
OA21x2_ASAP7_75t_L g394 ( .A1(n_353), .A2(n_343), .B(n_330), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_352), .B(n_343), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_357), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_357), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
NAND2x1_ASAP7_75t_L g402 ( .A(n_369), .B(n_342), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_369), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
OAI321xp33_ASAP7_75t_L g405 ( .A1(n_373), .A2(n_352), .A3(n_374), .B1(n_363), .B2(n_375), .C(n_361), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_357), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_351), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_372), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_377), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_377), .B(n_324), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_378), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_359), .B(n_358), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_407), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_407), .B(n_359), .Y(n_417) );
INVx4_ASAP7_75t_L g418 ( .A(n_388), .Y(n_418) );
NAND2x1_ASAP7_75t_SL g419 ( .A(n_403), .B(n_369), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_408), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_385), .B(n_359), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_385), .B(n_358), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_408), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_379), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_388), .B(n_366), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_408), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_415), .B(n_358), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_415), .B(n_358), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_385), .B(n_415), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_379), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_409), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_401), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_383), .B(n_358), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_380), .B(n_360), .Y(n_435) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_403), .B(n_366), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_383), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_384), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_396), .B(n_375), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_380), .B(n_360), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_380), .B(n_360), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_396), .B(n_378), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_387), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_399), .B(n_365), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_387), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_390), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_390), .B(n_362), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_403), .A2(n_373), .B1(n_370), .B2(n_374), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_397), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_394), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_399), .B(n_365), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_414), .B(n_365), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_405), .B(n_376), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_414), .B(n_365), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_397), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_403), .Y(n_458) );
NOR2xp33_ASAP7_75t_R g459 ( .A(n_388), .B(n_366), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_386), .B(n_361), .Y(n_460) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_386), .B(n_370), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_409), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_414), .B(n_365), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_400), .B(n_404), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_400), .B(n_362), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_404), .B(n_362), .Y(n_466) );
OR2x6_ASAP7_75t_L g467 ( .A(n_393), .B(n_364), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_393), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_440), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_437), .B(n_413), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_461), .B(n_388), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_424), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_429), .B(n_395), .Y(n_475) );
INVxp67_ASAP7_75t_L g476 ( .A(n_416), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_461), .A2(n_386), .B1(n_388), .B2(n_392), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_429), .B(n_395), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_431), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_435), .B(n_382), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_459), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_434), .B(n_386), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_438), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_461), .A2(n_388), .B(n_405), .C(n_398), .Y(n_488) );
NOR2xp33_ASAP7_75t_SL g489 ( .A(n_436), .B(n_388), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_434), .B(n_417), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_421), .B(n_386), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_468), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_439), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_417), .B(n_413), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_430), .B(n_410), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_445), .B(n_410), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_430), .B(n_412), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_433), .B(n_412), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_433), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_420), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_435), .B(n_389), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_447), .B(n_412), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_442), .B(n_389), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_464), .B(n_389), .Y(n_506) );
INVx3_ASAP7_75t_SL g507 ( .A(n_436), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_458), .B(n_398), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_464), .B(n_381), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_420), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_447), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_421), .B(n_381), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_468), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_422), .B(n_398), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_448), .Y(n_515) );
OAI211xp5_ASAP7_75t_L g516 ( .A1(n_450), .A2(n_402), .B(n_393), .C(n_392), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_422), .B(n_392), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_442), .B(n_381), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_443), .B(n_382), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_448), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_455), .B(n_460), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_451), .B(n_382), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_420), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_443), .B(n_406), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_427), .B(n_391), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_427), .B(n_391), .Y(n_526) );
NAND2x1_ASAP7_75t_SL g527 ( .A(n_418), .B(n_406), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_427), .B(n_406), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_451), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_469), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_521), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_475), .B(n_428), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_484), .B(n_449), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_493), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_475), .B(n_428), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_479), .B(n_428), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_513), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_525), .B(n_418), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_472), .Y(n_539) );
AOI21x1_ASAP7_75t_L g540 ( .A1(n_471), .A2(n_402), .B(n_467), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_502), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_521), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_507), .A2(n_436), .B1(n_425), .B2(n_458), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_526), .B(n_418), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_484), .Y(n_545) );
OAI21xp33_ASAP7_75t_L g546 ( .A1(n_488), .A2(n_419), .B(n_449), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_476), .B(n_460), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_507), .A2(n_425), .B1(n_458), .B2(n_418), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_479), .B(n_427), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_476), .B(n_466), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_501), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_473), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_474), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_513), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_478), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_483), .B(n_470), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_501), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_491), .B(n_428), .Y(n_559) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_527), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_480), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_487), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_514), .B(n_458), .Y(n_564) );
OA21x2_ASAP7_75t_SL g565 ( .A1(n_471), .A2(n_419), .B(n_425), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_490), .Y(n_566) );
XNOR2x1_ASAP7_75t_L g567 ( .A(n_492), .B(n_466), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_483), .B(n_457), .Y(n_568) );
OAI21xp33_ASAP7_75t_SL g569 ( .A1(n_477), .A2(n_467), .B(n_457), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_481), .B(n_465), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_510), .Y(n_571) );
NAND2xp33_ASAP7_75t_L g572 ( .A(n_488), .B(n_453), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_517), .B(n_463), .Y(n_573) );
AOI321xp33_ASAP7_75t_L g574 ( .A1(n_516), .A2(n_465), .A3(n_454), .B1(n_463), .B2(n_456), .C(n_453), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_499), .Y(n_575) );
INVxp33_ASAP7_75t_L g576 ( .A(n_489), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_494), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_528), .B(n_456), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_482), .B(n_446), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_481), .B(n_446), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_571), .Y(n_581) );
NOR2xp33_ASAP7_75t_SL g582 ( .A(n_543), .B(n_508), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_531), .B(n_503), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_579), .B(n_528), .Y(n_584) );
AOI21xp33_ASAP7_75t_L g585 ( .A1(n_531), .A2(n_497), .B(n_500), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_553), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_542), .B(n_524), .Y(n_587) );
AOI21xp33_ASAP7_75t_SL g588 ( .A1(n_569), .A2(n_508), .B(n_485), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_541), .Y(n_589) );
INVxp33_ASAP7_75t_L g590 ( .A(n_548), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_542), .A2(n_363), .B(n_353), .C(n_529), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_554), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_568), .B(n_524), .Y(n_593) );
OAI21xp33_ASAP7_75t_L g594 ( .A1(n_551), .A2(n_495), .B(n_512), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_560), .A2(n_508), .B(n_522), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_568), .A2(n_496), .B1(n_520), .B2(n_515), .C(n_511), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_534), .B(n_467), .Y(n_597) );
OAI221xp5_ASAP7_75t_SL g598 ( .A1(n_574), .A2(n_519), .B1(n_467), .B2(n_506), .C(n_509), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_537), .B(n_498), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_547), .A2(n_505), .B1(n_503), .B2(n_518), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_575), .B(n_518), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_552), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_576), .A2(n_572), .B(n_546), .C(n_560), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_579), .B(n_505), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
OAI32xp33_ASAP7_75t_L g606 ( .A1(n_576), .A2(n_504), .A3(n_510), .B1(n_523), .B2(n_454), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_561), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_540), .B(n_523), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_563), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_566), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_577), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_547), .A2(n_467), .B1(n_362), .B2(n_452), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_575), .B(n_423), .Y(n_614) );
AOI21xp5_ASAP7_75t_SL g615 ( .A1(n_609), .A2(n_552), .B(n_544), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_582), .A2(n_557), .B1(n_555), .B2(n_567), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_590), .A2(n_538), .B(n_544), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_583), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_590), .A2(n_587), .B1(n_599), .B2(n_595), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_598), .A2(n_538), .B(n_558), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_588), .A2(n_565), .B1(n_558), .B2(n_533), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g622 ( .A1(n_603), .A2(n_559), .B1(n_564), .B2(n_545), .C(n_539), .Y(n_622) );
AOI21xp33_ASAP7_75t_L g623 ( .A1(n_591), .A2(n_530), .B(n_452), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_599), .A2(n_532), .B1(n_535), .B2(n_536), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_602), .A2(n_452), .B(n_571), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_600), .A2(n_549), .B1(n_573), .B2(n_578), .Y(n_626) );
AOI311xp33_ASAP7_75t_L g627 ( .A1(n_585), .A2(n_580), .A3(n_570), .B(n_541), .C(n_550), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_596), .B(n_550), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_594), .A2(n_452), .B1(n_362), .B2(n_462), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_581), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_601), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_602), .A2(n_452), .B1(n_462), .B2(n_426), .C(n_423), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_593), .B(n_608), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_613), .A2(n_452), .B(n_411), .Y(n_634) );
OAI321xp33_ASAP7_75t_L g635 ( .A1(n_621), .A2(n_609), .A3(n_614), .B1(n_611), .B2(n_610), .C(n_612), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_615), .A2(n_597), .B(n_606), .C(n_605), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_622), .A2(n_607), .B(n_592), .C(n_586), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_619), .A2(n_617), .B1(n_620), .B2(n_634), .C(n_628), .Y(n_638) );
AOI211x1_ASAP7_75t_L g639 ( .A1(n_623), .A2(n_584), .B(n_604), .C(n_364), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_625), .B(n_589), .C(n_411), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_618), .A2(n_589), .B1(n_426), .B2(n_432), .C(n_462), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_616), .B(n_423), .Y(n_642) );
AOI222xp33_ASAP7_75t_L g643 ( .A1(n_631), .A2(n_426), .B1(n_432), .B2(n_441), .C1(n_394), .C2(n_356), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_633), .Y(n_644) );
AOI221x1_ASAP7_75t_L g645 ( .A1(n_627), .A2(n_432), .B1(n_441), .B2(n_394), .C(n_364), .Y(n_645) );
AOI211x1_ASAP7_75t_L g646 ( .A1(n_626), .A2(n_394), .B(n_356), .C(n_441), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_644), .B(n_629), .Y(n_647) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_636), .B(n_630), .Y(n_648) );
AOI221x1_ASAP7_75t_L g649 ( .A1(n_640), .A2(n_632), .B1(n_624), .B2(n_394), .C(n_356), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_637), .Y(n_650) );
NOR3xp33_ASAP7_75t_SL g651 ( .A(n_635), .B(n_632), .C(n_356), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_638), .A2(n_356), .B(n_371), .C(n_642), .Y(n_652) );
OR5x1_ASAP7_75t_L g653 ( .A(n_651), .B(n_639), .C(n_645), .D(n_646), .E(n_643), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_650), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_648), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_652), .B(n_647), .C(n_641), .Y(n_656) );
OR3x1_ASAP7_75t_L g657 ( .A(n_656), .B(n_649), .C(n_371), .Y(n_657) );
INVx4_ASAP7_75t_L g658 ( .A(n_654), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_658), .Y(n_659) );
INVx2_ASAP7_75t_SL g660 ( .A(n_657), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_661), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_662), .B(n_655), .Y(n_663) );
OAI21x1_ASAP7_75t_SL g664 ( .A1(n_663), .A2(n_660), .B(n_653), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_371), .B1(n_661), .B2(n_663), .Y(n_665) );
endmodule