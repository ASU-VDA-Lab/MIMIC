module fake_jpeg_2781_n_550 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_550);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_52),
.B(n_67),
.Y(n_132)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_53),
.Y(n_122)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_33),
.Y(n_61)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_76),
.B(n_98),
.Y(n_117)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_71),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_0),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_18),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_80),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_34),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_18),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_88),
.Y(n_115)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_95),
.Y(n_130)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_25),
.B(n_2),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_63),
.A2(n_41),
.B1(n_39),
.B2(n_37),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_121),
.A2(n_126),
.B1(n_146),
.B2(n_165),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_41),
.B1(n_37),
.B2(n_46),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g213 ( 
.A1(n_124),
.A2(n_51),
.B1(n_100),
.B2(n_102),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_40),
.B1(n_48),
.B2(n_28),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_54),
.B(n_40),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_70),
.A2(n_44),
.B1(n_39),
.B2(n_41),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_144),
.B1(n_162),
.B2(n_20),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_55),
.B(n_48),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_145),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_74),
.A2(n_51),
.B1(n_22),
.B2(n_36),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_142),
.A2(n_64),
.B1(n_62),
.B2(n_66),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_41),
.B1(n_39),
.B2(n_46),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_75),
.B(n_43),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_67),
.A2(n_39),
.B1(n_46),
.B2(n_45),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_43),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_38),
.Y(n_155)
);

NAND2x1p5_ASAP7_75t_L g157 ( 
.A(n_53),
.B(n_44),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_94),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_61),
.B(n_38),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_160),
.B(n_163),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_68),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_73),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_85),
.A2(n_44),
.B1(n_45),
.B2(n_28),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_144),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_166),
.B(n_180),
.Y(n_264)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_170),
.A2(n_201),
.B1(n_217),
.B2(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_114),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_171),
.B(n_189),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_174),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_106),
.A2(n_47),
.B(n_22),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_190),
.Y(n_232)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_176),
.Y(n_271)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_181),
.Y(n_269)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_183),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_105),
.B(n_47),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_198),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_121),
.A2(n_91),
.B1(n_84),
.B2(n_97),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_185),
.A2(n_213),
.B(n_223),
.Y(n_247)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_105),
.A2(n_103),
.B1(n_20),
.B2(n_45),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_187),
.A2(n_92),
.B(n_118),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_36),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_108),
.C(n_133),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_112),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_191),
.B(n_212),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_58),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

BUFx4f_ASAP7_75t_SL g197 ( 
.A(n_131),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_117),
.B(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_57),
.B1(n_96),
.B2(n_90),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_109),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_204),
.Y(n_265)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_206),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_139),
.A2(n_56),
.B1(n_83),
.B2(n_82),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_164),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_81),
.B1(n_79),
.B2(n_77),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_124),
.A2(n_59),
.B1(n_22),
.B2(n_36),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_123),
.B(n_102),
.Y(n_212)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_123),
.B(n_100),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_219),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_157),
.B(n_51),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_218),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_124),
.A2(n_127),
.B1(n_134),
.B2(n_110),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_51),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_116),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_111),
.B(n_69),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_116),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_225),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_125),
.B(n_69),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_226),
.B(n_122),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_170),
.A2(n_124),
.B1(n_120),
.B2(n_154),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_227),
.A2(n_250),
.B1(n_262),
.B2(n_278),
.Y(n_286)
);

AO22x1_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_116),
.B1(n_134),
.B2(n_154),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_228),
.B(n_276),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_233),
.B(n_241),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_156),
.B(n_125),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_237),
.A2(n_218),
.B(n_223),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_150),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_253),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_167),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_166),
.A2(n_137),
.B1(n_147),
.B2(n_151),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_184),
.B(n_216),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_207),
.A2(n_137),
.B1(n_147),
.B2(n_151),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_189),
.B(n_193),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_272),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_172),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_197),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_192),
.A2(n_127),
.B1(n_136),
.B2(n_152),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_274),
.B1(n_187),
.B2(n_218),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_193),
.B(n_111),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_210),
.A2(n_156),
.B1(n_122),
.B2(n_118),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_275),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_173),
.B(n_164),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_197),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_209),
.A2(n_148),
.B1(n_119),
.B2(n_27),
.Y(n_280)
);

AO21x2_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_213),
.B(n_185),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_281),
.B(n_292),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_282),
.A2(n_306),
.B1(n_231),
.B2(n_280),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_188),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_283),
.B(n_297),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_284),
.B(n_290),
.Y(n_369)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_288),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_236),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_246),
.A2(n_185),
.B1(n_213),
.B2(n_226),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_291),
.A2(n_294),
.B1(n_295),
.B2(n_302),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_227),
.A2(n_185),
.B1(n_186),
.B2(n_183),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_252),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_296),
.B(n_310),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_237),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_239),
.A2(n_223),
.B1(n_179),
.B2(n_178),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_317),
.B1(n_318),
.B2(n_325),
.Y(n_332)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_247),
.A2(n_278),
.B1(n_267),
.B2(n_264),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_235),
.B(n_205),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_303),
.B(n_309),
.Y(n_356)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_264),
.A2(n_181),
.B1(n_195),
.B2(n_176),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_252),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_230),
.B(n_168),
.C(n_174),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_260),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_247),
.A2(n_204),
.B1(n_214),
.B2(n_211),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_312),
.A2(n_327),
.B1(n_260),
.B2(n_279),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_315),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_242),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_314),
.B(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_230),
.B(n_253),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_254),
.B(n_220),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_264),
.A2(n_244),
.B1(n_263),
.B2(n_247),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_244),
.A2(n_148),
.B1(n_202),
.B2(n_203),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_238),
.B(n_78),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_228),
.C(n_233),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_242),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_322),
.Y(n_349)
);

OAI21xp33_ASAP7_75t_SL g321 ( 
.A1(n_232),
.A2(n_177),
.B(n_169),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_3),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_261),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_261),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_328),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_274),
.A2(n_272),
.B1(n_276),
.B2(n_248),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_259),
.A2(n_78),
.B1(n_27),
.B2(n_26),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_326),
.A2(n_304),
.B(n_313),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_250),
.A2(n_119),
.B1(n_27),
.B2(n_26),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_238),
.B(n_258),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_228),
.B(n_2),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_330),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_235),
.B(n_2),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_L g394 ( 
.A1(n_331),
.A2(n_370),
.B1(n_310),
.B2(n_296),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_338),
.C(n_354),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_262),
.B1(n_268),
.B2(n_251),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_334),
.A2(n_337),
.B1(n_294),
.B2(n_327),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_335),
.Y(n_405)
);

AOI22x1_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_251),
.B1(n_240),
.B2(n_269),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_229),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_291),
.A2(n_266),
.B1(n_269),
.B2(n_273),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_348),
.B1(n_334),
.B2(n_344),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_286),
.A2(n_243),
.B1(n_273),
.B2(n_271),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_340),
.A2(n_360),
.B1(n_372),
.B2(n_295),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_288),
.A2(n_231),
.B(n_243),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_312),
.B(n_329),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_271),
.B1(n_265),
.B2(n_279),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_347),
.A2(n_350),
.B1(n_359),
.B2(n_365),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_286),
.A2(n_229),
.B1(n_265),
.B2(n_271),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_299),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_301),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_328),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_297),
.A2(n_304),
.B1(n_325),
.B2(n_282),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_289),
.B(n_326),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_234),
.B1(n_256),
.B2(n_270),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_304),
.A2(n_234),
.B1(n_256),
.B2(n_270),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_285),
.B(n_311),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_364),
.C(n_8),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_27),
.C(n_26),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_294),
.A2(n_27),
.B1(n_26),
.B2(n_5),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_318),
.A2(n_27),
.B1(n_26),
.B2(n_5),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_SL g408 ( 
.A(n_371),
.B(n_373),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_294),
.A2(n_26),
.B1(n_4),
.B2(n_5),
.Y(n_372)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_363),
.Y(n_375)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_380),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_377),
.A2(n_378),
.B(n_399),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_379),
.A2(n_397),
.B1(n_406),
.B2(n_407),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_373),
.Y(n_380)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_349),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_389),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_284),
.Y(n_383)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_372),
.A2(n_294),
.B1(n_289),
.B2(n_290),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_384),
.A2(n_390),
.B1(n_392),
.B2(n_387),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_311),
.Y(n_385)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_336),
.Y(n_386)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_332),
.A2(n_294),
.B1(n_300),
.B2(n_316),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_387),
.A2(n_340),
.B1(n_346),
.B2(n_342),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_330),
.Y(n_388)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_332),
.A2(n_287),
.B1(n_293),
.B2(n_298),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_398),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_357),
.A2(n_320),
.B1(n_314),
.B2(n_292),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_369),
.B(n_309),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_395),
.B(n_396),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_356),
.B(n_307),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_345),
.A2(n_305),
.B1(n_323),
.B2(n_322),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_345),
.B(n_3),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_SL g399 ( 
.A(n_353),
.B(n_3),
.C(n_4),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_402),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_358),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_368),
.B(n_3),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_403),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_343),
.B(n_4),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_409),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_355),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_355),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_361),
.B(n_6),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_364),
.C(n_333),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_358),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_411),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_335),
.C(n_362),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_425),
.C(n_431),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_382),
.A2(n_408),
.B(n_353),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_421),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_416),
.B(n_375),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_418),
.A2(n_401),
.B1(n_386),
.B2(n_400),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_371),
.B(n_343),
.Y(n_421)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_354),
.C(n_360),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_348),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_426),
.B(n_389),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_337),
.B1(n_361),
.B2(n_339),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_428),
.A2(n_436),
.B1(n_440),
.B2(n_441),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_337),
.B(n_367),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_391),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_385),
.C(n_383),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_381),
.A2(n_374),
.B1(n_367),
.B2(n_366),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_378),
.C(n_390),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_388),
.C(n_399),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_379),
.A2(n_341),
.B1(n_366),
.B2(n_351),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_376),
.A2(n_341),
.B1(n_374),
.B2(n_11),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_424),
.A2(n_377),
.B1(n_402),
.B2(n_411),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_445),
.A2(n_423),
.B1(n_430),
.B2(n_421),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_448),
.B(n_456),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_418),
.A2(n_380),
.B1(n_395),
.B2(n_396),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_449),
.A2(n_454),
.B1(n_466),
.B2(n_429),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_457),
.C(n_458),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_443),
.B(n_403),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_451),
.B(n_465),
.Y(n_483)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_452),
.A2(n_453),
.B1(n_455),
.B2(n_461),
.Y(n_487)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_398),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_426),
.B(n_409),
.C(n_404),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_407),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_464),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_425),
.B(n_406),
.C(n_10),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_462),
.C(n_468),
.Y(n_486)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_8),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_8),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_443),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_414),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_11),
.C(n_13),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_412),
.B(n_13),
.C(n_14),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_415),
.C(n_437),
.Y(n_488)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_471),
.A2(n_480),
.B1(n_485),
.B2(n_459),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_463),
.Y(n_474)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_444),
.A2(n_424),
.B1(n_422),
.B2(n_413),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_475),
.A2(n_482),
.B1(n_441),
.B2(n_448),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_445),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_477),
.B(n_491),
.Y(n_499)
);

AOI221xp5_ASAP7_75t_L g480 ( 
.A1(n_455),
.A2(n_438),
.B1(n_439),
.B2(n_419),
.C(n_413),
.Y(n_480)
);

BUFx12_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_481),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_444),
.A2(n_422),
.B1(n_440),
.B2(n_438),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_427),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_453),
.A2(n_428),
.B1(n_436),
.B2(n_420),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_469),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_447),
.B(n_454),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_489),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_461),
.A2(n_427),
.B(n_415),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_464),
.B(n_434),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_431),
.C(n_433),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_491),
.B(n_446),
.C(n_456),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_503),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_495),
.A2(n_496),
.B1(n_507),
.B2(n_489),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_497),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_446),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_473),
.C(n_490),
.Y(n_512)
);

FAx1_ASAP7_75t_SL g503 ( 
.A(n_473),
.B(n_458),
.CI(n_433),
.CON(n_503),
.SN(n_503)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_505),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_419),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_508),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_482),
.A2(n_475),
.B1(n_489),
.B2(n_471),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_479),
.B(n_462),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_460),
.C(n_468),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_509),
.B(n_486),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_434),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_510),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_512),
.B(n_517),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_513),
.A2(n_500),
.B1(n_493),
.B2(n_497),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_514),
.B(n_518),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_498),
.B(n_483),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_488),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_494),
.B(n_487),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_519),
.A2(n_522),
.B(n_503),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_492),
.C(n_486),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_523),
.C(n_509),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_502),
.A2(n_472),
.B(n_485),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_472),
.C(n_481),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_526),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_510),
.C(n_507),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_511),
.A2(n_500),
.B1(n_496),
.B2(n_481),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_528),
.B(n_529),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_442),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_533),
.Y(n_540)
);

OAI21x1_ASAP7_75t_SL g535 ( 
.A1(n_532),
.A2(n_516),
.B(n_522),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_503),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_481),
.C(n_437),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g537 ( 
.A1(n_534),
.A2(n_524),
.B(n_442),
.Y(n_537)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_535),
.A2(n_526),
.B(n_534),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_537),
.A2(n_531),
.B(n_533),
.Y(n_541)
);

A2O1A1Ixp33_ASAP7_75t_SL g538 ( 
.A1(n_527),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_538)
);

AOI31xp33_ASAP7_75t_L g544 ( 
.A1(n_538),
.A2(n_15),
.A3(n_16),
.B(n_17),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_541),
.B(n_542),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_528),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_544),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_545),
.B(n_539),
.C(n_540),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_547),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_548),
.A2(n_546),
.B(n_17),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_17),
.Y(n_550)
);


endmodule