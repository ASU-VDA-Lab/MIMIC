module fake_netlist_6_4258_n_1295 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1295);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1295;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_304;
wire n_694;
wire n_1294;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_177;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1287;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_172;
wire n_1272;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_50),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_26),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_102),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_71),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_38),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_40),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_72),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_116),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_31),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_74),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_63),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_17),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_32),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_134),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_68),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_110),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_93),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_38),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_81),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_100),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_162),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_105),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_130),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_50),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_46),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_85),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_62),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_112),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_151),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_139),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_65),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_41),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_45),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_33),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_107),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_159),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_7),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_113),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_106),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_16),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_164),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_26),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_21),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_97),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_78),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_161),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_66),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_148),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_31),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_114),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_101),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_43),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_165),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_20),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_146),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_152),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_109),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_18),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_7),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_33),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_158),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_86),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_163),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_64),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_28),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_4),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_133),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_154),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_96),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_10),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_45),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_55),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_145),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_79),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_88),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_147),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_22),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_140),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_27),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_60),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_10),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_25),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_19),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_36),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_0),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_43),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_149),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_99),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_42),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_187),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_178),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_181),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_181),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_197),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_216),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_231),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_190),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_180),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_190),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_189),
.B(n_0),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_195),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_204),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_211),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_185),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_272),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_172),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_191),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_179),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_204),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_227),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_227),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_195),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_211),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_251),
.B(n_1),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_189),
.B(n_1),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_215),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_215),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_193),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_171),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_218),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_251),
.B(n_2),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_174),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_200),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_177),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_173),
.B(n_4),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_218),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_230),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_212),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_214),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_223),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_173),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_230),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_233),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_233),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_173),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_182),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_226),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_203),
.B(n_5),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_183),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_184),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_243),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_232),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_243),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_250),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_241),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_242),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_186),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_175),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_188),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_228),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_253),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_250),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_192),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_260),
.B(n_5),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_257),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_252),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_252),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_258),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_266),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_196),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_236),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_254),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_260),
.B(n_6),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_236),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_203),
.B(n_6),
.Y(n_371)
);

INVxp33_ASAP7_75t_SL g372 ( 
.A(n_270),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_271),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_254),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_198),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_262),
.B(n_8),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_275),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_225),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_281),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_262),
.B(n_8),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_278),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_279),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_294),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_294),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_201),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_176),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_294),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_306),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_264),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g391 ( 
.A1(n_295),
.A2(n_248),
.B(n_239),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_292),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_379),
.A2(n_288),
.B1(n_285),
.B2(n_239),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_300),
.B(n_303),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_337),
.B(n_264),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_213),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

OA21x2_ASAP7_75t_L g405 ( 
.A1(n_305),
.A2(n_259),
.B(n_248),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_316),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_199),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_SL g408 ( 
.A(n_302),
.B(n_286),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_317),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_337),
.B(n_289),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_318),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_304),
.B(n_213),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_341),
.B(n_289),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_348),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_202),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_293),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

CKINVDCx6p67_ASAP7_75t_R g424 ( 
.A(n_311),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_293),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_340),
.B(n_290),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_347),
.Y(n_428)
);

CKINVDCx8_ASAP7_75t_R g429 ( 
.A(n_356),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_349),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_321),
.B(n_287),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_368),
.Y(n_436)
);

AND2x2_ASAP7_75t_SL g437 ( 
.A(n_376),
.B(n_244),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_364),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_307),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_353),
.B(n_290),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_301),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_309),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_327),
.Y(n_448)
);

INVx6_ASAP7_75t_L g449 ( 
.A(n_299),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_319),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_398),
.A2(n_314),
.B1(n_312),
.B2(n_308),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_388),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_444),
.B(n_372),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_244),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_386),
.B(n_372),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_261),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_383),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_386),
.B(n_373),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_437),
.A2(n_291),
.B1(n_285),
.B2(n_265),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_261),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_273),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_273),
.Y(n_469)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_444),
.B(n_373),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_396),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_274),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_274),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_427),
.B(n_282),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_388),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_444),
.B(n_301),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_444),
.B(n_310),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_402),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_396),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_390),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_383),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_383),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_415),
.B(n_282),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_435),
.B(n_359),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_328),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_407),
.B(n_330),
.Y(n_507)
);

AND2x6_ASAP7_75t_L g508 ( 
.A(n_389),
.B(n_201),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_405),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_444),
.B(n_310),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_409),
.Y(n_512)
);

OAI21xp33_ASAP7_75t_SL g513 ( 
.A1(n_414),
.A2(n_265),
.B(n_259),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_437),
.A2(n_291),
.B1(n_221),
.B2(n_201),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_393),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_409),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_383),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_415),
.B(n_201),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_437),
.A2(n_221),
.B1(n_201),
.B2(n_377),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_444),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_415),
.B(n_221),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_445),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_488),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_514),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_459),
.B(n_445),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_463),
.A2(n_414),
.B1(n_437),
.B2(n_445),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_470),
.B(n_444),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_445),
.Y(n_530)
);

A2O1A1Ixp33_ASAP7_75t_L g531 ( 
.A1(n_513),
.A2(n_414),
.B(n_407),
.C(n_389),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_464),
.B(n_451),
.C(n_444),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_414),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_457),
.B(n_445),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_488),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_514),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_470),
.B(n_502),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_499),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_470),
.B(n_451),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_488),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_493),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_470),
.B(n_389),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_502),
.B(n_451),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_499),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_502),
.B(n_443),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_496),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_502),
.B(n_451),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_494),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_451),
.C(n_324),
.Y(n_551)
);

NOR2xp67_ASAP7_75t_L g552 ( 
.A(n_504),
.B(n_313),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_496),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_466),
.B(n_443),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_455),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_471),
.B(n_451),
.Y(n_556)
);

OR2x2_ASAP7_75t_SL g557 ( 
.A(n_475),
.B(n_451),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_496),
.Y(n_558)
);

A2O1A1Ixp33_ASAP7_75t_L g559 ( 
.A1(n_513),
.A2(n_443),
.B(n_385),
.C(n_419),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_487),
.B(n_451),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_489),
.A2(n_426),
.B1(n_420),
.B2(n_345),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_511),
.B(n_420),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_475),
.Y(n_563)
);

AND2x6_ASAP7_75t_SL g564 ( 
.A(n_494),
.B(n_450),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_497),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_522),
.B(n_420),
.Y(n_566)
);

BUFx5_ASAP7_75t_L g567 ( 
.A(n_473),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_466),
.B(n_419),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_455),
.B(n_354),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_515),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_460),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_466),
.B(n_385),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_466),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_460),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_483),
.B(n_446),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_517),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_483),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_483),
.B(n_432),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_483),
.B(n_432),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_522),
.B(n_426),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_522),
.B(n_313),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_517),
.B(n_446),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_473),
.B(n_426),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_474),
.B(n_221),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_517),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_474),
.B(n_417),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_458),
.B(n_446),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_458),
.B(n_432),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_476),
.A2(n_346),
.B1(n_355),
.B2(n_342),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_461),
.B(n_432),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_476),
.B(n_417),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_481),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_481),
.B(n_438),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_461),
.Y(n_595)
);

NOR2x1_ASAP7_75t_L g596 ( 
.A(n_482),
.B(n_366),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_482),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_497),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_465),
.B(n_432),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_465),
.B(n_422),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_485),
.B(n_438),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_469),
.B(n_478),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_469),
.B(n_375),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_478),
.B(n_422),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_503),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_490),
.A2(n_297),
.B1(n_298),
.B2(n_408),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_479),
.B(n_422),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_479),
.B(n_422),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_490),
.B(n_422),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_508),
.B(n_205),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_491),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_491),
.B(n_425),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_492),
.B(n_324),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_492),
.B(n_425),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_495),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_495),
.B(n_425),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_503),
.B(n_398),
.C(n_408),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_509),
.B(n_425),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_509),
.B(n_221),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_L g621 ( 
.A(n_510),
.B(n_442),
.C(n_334),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_528),
.B(n_510),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_550),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_537),
.A2(n_501),
.B(n_401),
.Y(n_624)
);

O2A1O1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_531),
.A2(n_520),
.B(n_523),
.C(n_393),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_584),
.A2(n_520),
.B(n_523),
.C(n_393),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_527),
.B(n_329),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_527),
.B(n_453),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_530),
.B(n_453),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_555),
.B(n_329),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_530),
.B(n_453),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_606),
.B(n_453),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_574),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_603),
.A2(n_501),
.B(n_401),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_569),
.B(n_334),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_587),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_573),
.A2(n_501),
.B(n_401),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_462),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_567),
.B(n_462),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_543),
.A2(n_501),
.B(n_401),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_578),
.B(n_400),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_576),
.B(n_400),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_533),
.A2(n_401),
.B1(n_449),
.B2(n_429),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_585),
.A2(n_456),
.B(n_454),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_SL g647 ( 
.A1(n_559),
.A2(n_229),
.B(n_194),
.C(n_440),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_588),
.B(n_462),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_536),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_583),
.B(n_462),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_524),
.B(n_467),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_525),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_589),
.A2(n_401),
.B(n_454),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_585),
.A2(n_456),
.B(n_454),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_614),
.B(n_467),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_584),
.A2(n_428),
.B(n_430),
.C(n_421),
.Y(n_656)
);

O2A1O1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_587),
.A2(n_428),
.B(n_430),
.C(n_421),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_620),
.A2(n_468),
.B(n_456),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_620),
.A2(n_472),
.B(n_468),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_541),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_538),
.B(n_545),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_563),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_614),
.B(n_467),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_549),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_590),
.B(n_335),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_591),
.A2(n_401),
.B(n_468),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_607),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_554),
.B(n_568),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_600),
.A2(n_477),
.B(n_472),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_570),
.Y(n_670)
);

O2A1O1Ixp5_ASAP7_75t_L g671 ( 
.A1(n_539),
.A2(n_472),
.B(n_477),
.C(n_480),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_567),
.B(n_534),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_542),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_535),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_567),
.B(n_467),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_557),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_567),
.B(n_500),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_567),
.B(n_500),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_567),
.B(n_500),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_601),
.A2(n_480),
.B(n_477),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_542),
.B(n_500),
.Y(n_681)
);

A2O1A1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_592),
.A2(n_416),
.B(n_400),
.C(n_411),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_535),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_540),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_534),
.A2(n_508),
.B1(n_449),
.B2(n_399),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_556),
.B(n_519),
.Y(n_686)
);

BUFx8_ASAP7_75t_L g687 ( 
.A(n_564),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_540),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_547),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_605),
.A2(n_484),
.B(n_480),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_608),
.A2(n_486),
.B(n_484),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_609),
.A2(n_486),
.B(n_484),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_539),
.A2(n_486),
.B(n_519),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_593),
.B(n_425),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_556),
.A2(n_427),
.B(n_416),
.C(n_411),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_592),
.B(n_594),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_547),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_553),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_529),
.A2(n_519),
.B(n_506),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_594),
.B(n_335),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_544),
.A2(n_519),
.B(n_506),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_593),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_560),
.A2(n_416),
.B(n_411),
.C(n_450),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_542),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_546),
.B(n_602),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_561),
.B(n_424),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_553),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_548),
.A2(n_519),
.B(n_506),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_558),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_542),
.Y(n_710)
);

AO21x1_ASAP7_75t_L g711 ( 
.A1(n_560),
.A2(n_512),
.B(n_498),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_602),
.B(n_508),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_571),
.Y(n_713)
);

AOI21x1_ASAP7_75t_L g714 ( 
.A1(n_610),
.A2(n_512),
.B(n_498),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_604),
.B(n_336),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_562),
.Y(n_716)
);

AOI21x1_ASAP7_75t_L g717 ( 
.A1(n_613),
.A2(n_512),
.B(n_498),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_579),
.A2(n_519),
.B(n_518),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_558),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_532),
.A2(n_449),
.B1(n_429),
.B2(n_392),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_552),
.B(n_452),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_551),
.B(n_452),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_704),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_627),
.A2(n_618),
.B(n_596),
.C(n_621),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_639),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_644),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_702),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_627),
.A2(n_581),
.B1(n_580),
.B2(n_566),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_668),
.A2(n_575),
.B(n_571),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_705),
.A2(n_599),
.B1(n_597),
.B2(n_616),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_649),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_700),
.A2(n_581),
.B1(n_577),
.B2(n_586),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_700),
.B(n_582),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_634),
.A2(n_575),
.B(n_612),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_643),
.A2(n_508),
.B1(n_611),
.B2(n_399),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_648),
.A2(n_617),
.B(n_615),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_664),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_670),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_L g739 ( 
.A(n_710),
.B(n_565),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_630),
.B(n_392),
.Y(n_740)
);

OAI21xp33_ASAP7_75t_L g741 ( 
.A1(n_635),
.A2(n_343),
.B(n_336),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_702),
.A2(n_619),
.B1(n_429),
.B2(n_572),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_623),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_630),
.B(n_440),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_636),
.A2(n_598),
.B1(n_572),
.B2(n_565),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_704),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_637),
.A2(n_598),
.B(n_387),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_674),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_696),
.B(n_399),
.Y(n_749)
);

AO32x1_ASAP7_75t_L g750 ( 
.A1(n_645),
.A2(n_418),
.A3(n_447),
.B1(n_448),
.B2(n_518),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_623),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_636),
.B(n_399),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_622),
.A2(n_518),
.B(n_508),
.Y(n_753)
);

INVx6_ASAP7_75t_L g754 ( 
.A(n_687),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_704),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_643),
.B(n_399),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_672),
.A2(n_387),
.B(n_383),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_721),
.B(n_343),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_635),
.B(n_424),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_672),
.A2(n_387),
.B(n_383),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_704),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_660),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_710),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_676),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_716),
.B(n_351),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_667),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_665),
.B(n_424),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_642),
.B(n_351),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_707),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_650),
.A2(n_624),
.B(n_686),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_661),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_686),
.A2(n_387),
.B(n_384),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_652),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_622),
.A2(n_449),
.B1(n_352),
.B2(n_361),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_662),
.Y(n_775)
);

OR2x6_ASAP7_75t_L g776 ( 
.A(n_642),
.B(n_449),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_665),
.B(n_352),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_675),
.A2(n_387),
.B(n_384),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_722),
.B(n_361),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_715),
.B(n_365),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_712),
.A2(n_449),
.B1(n_365),
.B2(n_377),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_678),
.A2(n_387),
.B(n_384),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_638),
.B(n_381),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_SL g784 ( 
.A(n_706),
.B(n_447),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_715),
.B(n_381),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_720),
.A2(n_508),
.B1(n_382),
.B2(n_418),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_683),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_673),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_628),
.B(n_382),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_633),
.B(n_448),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_684),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_625),
.A2(n_423),
.B(n_439),
.C(n_436),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_632),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_713),
.A2(n_267),
.B1(n_207),
.B2(n_208),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_688),
.Y(n_795)
);

OAI21xp33_ASAP7_75t_L g796 ( 
.A1(n_682),
.A2(n_397),
.B(n_394),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_734),
.A2(n_717),
.B(n_714),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_726),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_763),
.B(n_682),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_747),
.A2(n_693),
.B(n_659),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_770),
.A2(n_631),
.B(n_629),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_777),
.A2(n_713),
.B1(n_673),
.B2(n_695),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_775),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_757),
.A2(n_671),
.B(n_718),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_760),
.A2(n_671),
.B(n_680),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_SL g806 ( 
.A1(n_724),
.A2(n_703),
.B(n_694),
.C(n_655),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_763),
.B(n_640),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_789),
.B(n_657),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_729),
.A2(n_736),
.B(n_733),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_759),
.A2(n_647),
.B(n_656),
.C(n_663),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_730),
.A2(n_641),
.B(n_651),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_783),
.B(n_689),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_776),
.B(n_697),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_728),
.A2(n_666),
.B(n_653),
.Y(n_814)
);

BUFx12f_ASAP7_75t_L g815 ( 
.A(n_754),
.Y(n_815)
);

AOI21x1_ASAP7_75t_SL g816 ( 
.A1(n_779),
.A2(n_647),
.B(n_711),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_728),
.A2(n_626),
.B(n_690),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_749),
.A2(n_677),
.B(n_640),
.Y(n_818)
);

OA21x2_ASAP7_75t_L g819 ( 
.A1(n_792),
.A2(n_669),
.B(n_691),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_772),
.A2(n_692),
.B(n_699),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_731),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_732),
.A2(n_685),
.B(n_701),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_764),
.Y(n_823)
);

AO21x2_ASAP7_75t_L g824 ( 
.A1(n_796),
.A2(n_654),
.B(n_646),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_763),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_751),
.Y(n_826)
);

BUFx4_ASAP7_75t_SL g827 ( 
.A(n_762),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_778),
.A2(n_708),
.B(n_658),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_793),
.B(n_698),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_753),
.A2(n_679),
.B(n_677),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_784),
.A2(n_679),
.B(n_681),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_758),
.B(n_709),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_776),
.B(n_719),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_723),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_740),
.A2(n_687),
.B1(n_276),
.B2(n_269),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_764),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_737),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_782),
.A2(n_681),
.B(n_423),
.Y(n_838)
);

AO21x1_ASAP7_75t_L g839 ( 
.A1(n_732),
.A2(n_397),
.B(n_394),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_752),
.A2(n_742),
.B(n_786),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_776),
.B(n_412),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_786),
.A2(n_508),
.B(n_423),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_738),
.Y(n_843)
);

AOI221xp5_ASAP7_75t_L g844 ( 
.A1(n_767),
.A2(n_410),
.B1(n_403),
.B2(n_404),
.C(n_406),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_744),
.B(n_412),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_748),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_735),
.A2(n_756),
.B(n_745),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_769),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_743),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_766),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_750),
.A2(n_387),
.B(n_413),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_739),
.A2(n_395),
.B(n_412),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_L g853 ( 
.A(n_741),
.B(n_404),
.C(n_403),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_781),
.A2(n_508),
.B(n_434),
.Y(n_854)
);

AO21x2_ASAP7_75t_L g855 ( 
.A1(n_796),
.A2(n_410),
.B(n_406),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_771),
.B(n_433),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_790),
.A2(n_439),
.B(n_436),
.C(n_434),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_727),
.B(n_433),
.Y(n_858)
);

AO21x2_ASAP7_75t_L g859 ( 
.A1(n_750),
.A2(n_434),
.B(n_433),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_827),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_849),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_850),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_834),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_L g864 ( 
.A1(n_835),
.A2(n_780),
.B1(n_785),
.B2(n_768),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_840),
.A2(n_774),
.B1(n_791),
.B2(n_765),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_825),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_850),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_808),
.A2(n_764),
.B1(n_794),
.B2(n_788),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_799),
.A2(n_754),
.B1(n_788),
.B2(n_755),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_798),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_821),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_815),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_853),
.A2(n_795),
.B1(n_787),
.B2(n_773),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_837),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_843),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_815),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_814),
.A2(n_725),
.B1(n_436),
.B2(n_439),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_826),
.B(n_755),
.Y(n_878)
);

INVx8_ASAP7_75t_L g879 ( 
.A(n_813),
.Y(n_879)
);

OAI22xp33_ASAP7_75t_SL g880 ( 
.A1(n_812),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_832),
.A2(n_761),
.B1(n_723),
.B2(n_746),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_799),
.A2(n_395),
.B1(n_431),
.B2(n_413),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_817),
.A2(n_395),
.B1(n_431),
.B2(n_413),
.Y(n_883)
);

CKINVDCx11_ASAP7_75t_R g884 ( 
.A(n_803),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_825),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_839),
.A2(n_413),
.B1(n_431),
.B2(n_746),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_826),
.A2(n_761),
.B1(n_723),
.B2(n_746),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_846),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_803),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_848),
.Y(n_890)
);

CKINVDCx11_ASAP7_75t_R g891 ( 
.A(n_836),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_841),
.A2(n_247),
.B1(n_219),
.B2(n_220),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_SL g893 ( 
.A1(n_802),
.A2(n_761),
.B1(n_246),
.B2(n_280),
.Y(n_893)
);

INVx6_ASAP7_75t_L g894 ( 
.A(n_836),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_829),
.A2(n_249),
.B1(n_222),
.B2(n_224),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_855),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_823),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_858),
.Y(n_898)
);

BUFx8_ASAP7_75t_SL g899 ( 
.A(n_841),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_856),
.Y(n_900)
);

BUFx6f_ASAP7_75t_SL g901 ( 
.A(n_841),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_822),
.A2(n_413),
.B1(n_431),
.B2(n_256),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_807),
.A2(n_255),
.B1(n_234),
.B2(n_235),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_855),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_834),
.Y(n_905)
);

BUFx10_ASAP7_75t_L g906 ( 
.A(n_813),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_834),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_845),
.A2(n_413),
.B1(n_431),
.B2(n_268),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_807),
.Y(n_909)
);

OAI21xp33_ASAP7_75t_L g910 ( 
.A1(n_845),
.A2(n_263),
.B(n_237),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_859),
.Y(n_911)
);

INVx6_ASAP7_75t_L g912 ( 
.A(n_813),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_833),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_831),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_833),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_833),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_859),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_857),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_857),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_818),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_852),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_838),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_SL g923 ( 
.A1(n_842),
.A2(n_277),
.B1(n_245),
.B2(n_240),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_SL g924 ( 
.A1(n_847),
.A2(n_238),
.B1(n_217),
.B2(n_750),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_810),
.A2(n_431),
.B1(n_413),
.B2(n_409),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_819),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_911),
.B(n_824),
.Y(n_927)
);

AO21x2_ASAP7_75t_L g928 ( 
.A1(n_904),
.A2(n_809),
.B(n_801),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_896),
.A2(n_797),
.B(n_811),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_922),
.B(n_838),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_896),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_865),
.A2(n_806),
.B(n_830),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_864),
.B(n_806),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_914),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_911),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_917),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_917),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_SL g938 ( 
.A1(n_920),
.A2(n_819),
.B1(n_854),
.B2(n_851),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_925),
.A2(n_797),
.B(n_800),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_922),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_926),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_870),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_926),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_921),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_870),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_874),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_874),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_875),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_875),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_916),
.B(n_804),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_888),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_888),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_871),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_865),
.A2(n_844),
.B1(n_824),
.B2(n_819),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_890),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_909),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_918),
.B(n_805),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_919),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_898),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_886),
.A2(n_820),
.B(n_805),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_900),
.Y(n_961)
);

NOR2x1_ASAP7_75t_SL g962 ( 
.A(n_868),
.B(n_816),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_913),
.B(n_804),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_915),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_877),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_877),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_916),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_861),
.B(n_9),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_873),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_878),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_879),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_912),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_912),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_970),
.B(n_897),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_952),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_933),
.A2(n_902),
.B(n_893),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_952),
.Y(n_977)
);

CKINVDCx11_ASAP7_75t_R g978 ( 
.A(n_934),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_933),
.A2(n_902),
.B(n_924),
.C(n_923),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_938),
.A2(n_882),
.B(n_869),
.C(n_886),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_938),
.A2(n_882),
.B(n_910),
.C(n_908),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_932),
.A2(n_883),
.B(n_880),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_970),
.B(n_912),
.Y(n_983)
);

NOR2x1_ASAP7_75t_SL g984 ( 
.A(n_934),
.B(n_887),
.Y(n_984)
);

BUFx2_ASAP7_75t_R g985 ( 
.A(n_934),
.Y(n_985)
);

NOR2x1_ASAP7_75t_SL g986 ( 
.A(n_934),
.B(n_940),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_954),
.A2(n_905),
.B1(n_889),
.B2(n_867),
.Y(n_987)
);

AO21x2_ASAP7_75t_L g988 ( 
.A1(n_962),
.A2(n_820),
.B(n_828),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_959),
.B(n_881),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_968),
.A2(n_895),
.B1(n_903),
.B2(n_908),
.C(n_892),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_961),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_967),
.B(n_906),
.Y(n_992)
);

NOR2x1_ASAP7_75t_SL g993 ( 
.A(n_940),
.B(n_907),
.Y(n_993)
);

AOI221xp5_ASAP7_75t_L g994 ( 
.A1(n_968),
.A2(n_901),
.B1(n_879),
.B2(n_872),
.C(n_876),
.Y(n_994)
);

AND2x6_ASAP7_75t_L g995 ( 
.A(n_958),
.B(n_863),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_932),
.A2(n_862),
.B(n_828),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_959),
.B(n_879),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_951),
.B(n_885),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_951),
.B(n_885),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_951),
.B(n_885),
.Y(n_1000)
);

AO21x2_ASAP7_75t_L g1001 ( 
.A1(n_962),
.A2(n_883),
.B(n_906),
.Y(n_1001)
);

AOI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_954),
.A2(n_901),
.B1(n_885),
.B2(n_866),
.C(n_413),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_969),
.A2(n_863),
.B(n_866),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_973),
.A2(n_972),
.B1(n_884),
.B2(n_969),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_951),
.B(n_907),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_L g1006 ( 
.A(n_961),
.B(n_884),
.C(n_891),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_967),
.B(n_972),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_949),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_967),
.B(n_894),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_L g1010 ( 
.A(n_971),
.B(n_965),
.Y(n_1010)
);

AOI211xp5_ASAP7_75t_L g1011 ( 
.A1(n_972),
.A2(n_860),
.B(n_409),
.C(n_13),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_942),
.B(n_894),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_953),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_942),
.B(n_894),
.Y(n_1014)
);

NOR2x1_ASAP7_75t_SL g1015 ( 
.A(n_940),
.B(n_958),
.Y(n_1015)
);

BUFx12f_ASAP7_75t_L g1016 ( 
.A(n_971),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_929),
.A2(n_899),
.B(n_891),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_967),
.B(n_11),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_929),
.A2(n_899),
.B(n_409),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_1013),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1007),
.B(n_927),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_SL g1022 ( 
.A1(n_987),
.A2(n_965),
.B1(n_966),
.B2(n_971),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1008),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_991),
.B(n_950),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1019),
.B(n_927),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_1015),
.B(n_950),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_975),
.B(n_977),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_998),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_991),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1019),
.B(n_927),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_995),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1019),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_976),
.A2(n_973),
.B1(n_972),
.B2(n_950),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_995),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_999),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_995),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_988),
.B(n_941),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_995),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_1017),
.B(n_950),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_995),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_1006),
.B(n_941),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1005),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_1000),
.B(n_931),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_988),
.B(n_941),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1012),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1014),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_979),
.A2(n_966),
.B(n_963),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_996),
.B(n_953),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1025),
.B(n_941),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1029),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1021),
.B(n_1035),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1029),
.B(n_989),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1025),
.B(n_943),
.Y(n_1053)
);

INVx5_ASAP7_75t_SL g1054 ( 
.A(n_1026),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1029),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1025),
.B(n_1030),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1022),
.A2(n_1011),
.B1(n_980),
.B2(n_981),
.Y(n_1057)
);

OAI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_1047),
.A2(n_990),
.B1(n_979),
.B2(n_981),
.C(n_982),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1030),
.B(n_943),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1020),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1020),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1020),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_1032),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1021),
.B(n_1035),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1023),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_1026),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_1026),
.Y(n_1067)
);

OAI211xp5_ASAP7_75t_L g1068 ( 
.A1(n_1047),
.A2(n_980),
.B(n_1002),
.C(n_978),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1030),
.B(n_1021),
.Y(n_1069)
);

AO22x1_ASAP7_75t_L g1070 ( 
.A1(n_1046),
.A2(n_1003),
.B1(n_985),
.B2(n_989),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1028),
.B(n_986),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1024),
.B(n_943),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_1027),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_1057),
.B(n_1041),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1058),
.B(n_978),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1052),
.B(n_1046),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1060),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1058),
.B(n_1041),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1052),
.B(n_1028),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1071),
.B(n_1045),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1071),
.B(n_1045),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1060),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1051),
.B(n_1042),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1073),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1051),
.B(n_1042),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1064),
.B(n_1039),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1064),
.B(n_1039),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1086),
.B(n_1054),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1087),
.B(n_1067),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1074),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_1074),
.B(n_1057),
.C(n_1068),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_1084),
.Y(n_1092)
);

OAI21xp33_ASAP7_75t_L g1093 ( 
.A1(n_1078),
.A2(n_1068),
.B(n_1033),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1083),
.B(n_1054),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1079),
.B(n_1073),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1090),
.B(n_1078),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1088),
.B(n_1067),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1092),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1092),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1093),
.B(n_1075),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1094),
.B(n_1054),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1098),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1098),
.Y(n_1103)
);

AOI222xp33_ASAP7_75t_L g1104 ( 
.A1(n_1100),
.A2(n_1091),
.B1(n_1096),
.B2(n_1075),
.C1(n_1099),
.C2(n_1070),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1097),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1097),
.A2(n_1095),
.B(n_994),
.C(n_1076),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1101),
.A2(n_1054),
.B1(n_1022),
.B2(n_1089),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1100),
.A2(n_1010),
.B(n_1004),
.C(n_1048),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1100),
.B(n_1080),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1098),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1098),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1101),
.B(n_1089),
.Y(n_1112)
);

AOI211xp5_ASAP7_75t_SL g1113 ( 
.A1(n_1100),
.A2(n_1010),
.B(n_1048),
.C(n_1018),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1111),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1111),
.B(n_1077),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1112),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1105),
.B(n_1081),
.Y(n_1117)
);

OAI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1104),
.A2(n_1066),
.B1(n_1082),
.B2(n_1077),
.C(n_1045),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1109),
.B(n_1102),
.Y(n_1119)
);

OAI211xp5_ASAP7_75t_L g1120 ( 
.A1(n_1108),
.A2(n_1063),
.B(n_1066),
.C(n_974),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1108),
.A2(n_1063),
.B1(n_1054),
.B2(n_1066),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1109),
.B(n_1085),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1103),
.B(n_1082),
.Y(n_1123)
);

AO21x1_ASAP7_75t_L g1124 ( 
.A1(n_1110),
.A2(n_1062),
.B(n_1056),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1106),
.Y(n_1125)
);

OAI211xp5_ASAP7_75t_L g1126 ( 
.A1(n_1113),
.A2(n_1063),
.B(n_997),
.C(n_1034),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1107),
.B(n_1056),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_1111),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1111),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1111),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1128),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1125),
.A2(n_1070),
.B1(n_1062),
.B2(n_1050),
.C(n_1055),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1116),
.B(n_1056),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_1119),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1114),
.B(n_1069),
.Y(n_1135)
);

XNOR2x1_ASAP7_75t_L g1136 ( 
.A(n_1129),
.B(n_11),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1130),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1122),
.B(n_1069),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1117),
.B(n_1069),
.Y(n_1139)
);

AOI221xp5_ASAP7_75t_L g1140 ( 
.A1(n_1118),
.A2(n_1055),
.B1(n_1050),
.B2(n_1061),
.C(n_1060),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1115),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1115),
.Y(n_1142)
);

OAI21xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1127),
.A2(n_1061),
.B(n_1053),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1123),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1121),
.Y(n_1145)
);

NAND4xp25_ASAP7_75t_SL g1146 ( 
.A(n_1120),
.B(n_1126),
.C(n_1124),
.D(n_1121),
.Y(n_1146)
);

AOI32xp33_ASAP7_75t_L g1147 ( 
.A1(n_1125),
.A2(n_1059),
.A3(n_1053),
.B1(n_1049),
.B2(n_1061),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1125),
.A2(n_1063),
.B(n_1039),
.C(n_997),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1128),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1128),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1131),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1149),
.B(n_1063),
.C(n_955),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1134),
.B(n_983),
.C(n_973),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1150),
.B(n_1049),
.Y(n_1154)
);

NAND4xp25_ASAP7_75t_L g1155 ( 
.A(n_1145),
.B(n_1039),
.C(n_1026),
.D(n_1009),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1136),
.B(n_1065),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1144),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1132),
.A2(n_1039),
.B(n_1063),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1137),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1141),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1142),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1133),
.B(n_1049),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_L g1163 ( 
.A(n_1146),
.B(n_12),
.C(n_13),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1140),
.B(n_1063),
.C(n_955),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1138),
.B(n_1053),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1139),
.Y(n_1166)
);

NAND4xp25_ASAP7_75t_L g1167 ( 
.A(n_1135),
.B(n_1026),
.C(n_973),
.D(n_1038),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1143),
.B(n_1065),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1163),
.A2(n_1143),
.B1(n_1148),
.B2(n_1147),
.C(n_1065),
.Y(n_1169)
);

NOR3xp33_ASAP7_75t_L g1170 ( 
.A(n_1163),
.B(n_1034),
.C(n_1031),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1157),
.B(n_1059),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1166),
.A2(n_1036),
.B1(n_1040),
.B2(n_1038),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_SL g1173 ( 
.A(n_1161),
.B(n_1036),
.C(n_1031),
.Y(n_1173)
);

AOI211xp5_ASAP7_75t_L g1174 ( 
.A1(n_1151),
.A2(n_1156),
.B(n_1159),
.C(n_1160),
.Y(n_1174)
);

OAI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_1158),
.A2(n_1040),
.B1(n_1027),
.B2(n_971),
.C(n_1059),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1153),
.B(n_1072),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1154),
.B(n_12),
.Y(n_1177)
);

AOI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_1155),
.A2(n_1044),
.B1(n_1037),
.B2(n_1001),
.C(n_1032),
.Y(n_1178)
);

AOI21xp33_ASAP7_75t_L g1179 ( 
.A1(n_1152),
.A2(n_14),
.B(n_15),
.Y(n_1179)
);

OAI211xp5_ASAP7_75t_L g1180 ( 
.A1(n_1167),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1164),
.B(n_1044),
.C(n_1037),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_R g1182 ( 
.A(n_1165),
.B(n_17),
.Y(n_1182)
);

NAND4xp25_ASAP7_75t_L g1183 ( 
.A(n_1162),
.B(n_1024),
.C(n_992),
.D(n_1037),
.Y(n_1183)
);

AOI21xp33_ASAP7_75t_L g1184 ( 
.A1(n_1168),
.A2(n_18),
.B(n_20),
.Y(n_1184)
);

NOR4xp25_ASAP7_75t_L g1185 ( 
.A(n_1161),
.B(n_21),
.C(n_22),
.D(n_23),
.Y(n_1185)
);

OAI31xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1161),
.A2(n_984),
.A3(n_1072),
.B(n_1044),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1157),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1157),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1163),
.A2(n_1016),
.B1(n_1072),
.B2(n_1001),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1163),
.A2(n_1032),
.B1(n_956),
.B2(n_1023),
.C(n_27),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_R g1191 ( 
.A(n_1157),
.B(n_23),
.Y(n_1191)
);

OAI211xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1163),
.A2(n_24),
.B(n_25),
.C(n_28),
.Y(n_1192)
);

AOI311xp33_ASAP7_75t_L g1193 ( 
.A1(n_1163),
.A2(n_24),
.A3(n_29),
.B(n_30),
.C(n_32),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1192),
.A2(n_29),
.B(n_30),
.C(n_34),
.Y(n_1194)
);

OAI211xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1174),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1187),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.C(n_40),
.Y(n_1196)
);

OAI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1190),
.A2(n_971),
.B1(n_1043),
.B2(n_964),
.C(n_963),
.Y(n_1197)
);

AOI211xp5_ASAP7_75t_L g1198 ( 
.A1(n_1185),
.A2(n_37),
.B(n_39),
.C(n_41),
.Y(n_1198)
);

XNOR2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1188),
.B(n_42),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1177),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_1184),
.A2(n_44),
.B(n_47),
.C(n_48),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1170),
.B(n_44),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1191),
.Y(n_1203)
);

XOR2x2_ASAP7_75t_L g1204 ( 
.A(n_1189),
.B(n_48),
.Y(n_1204)
);

OAI221xp5_ASAP7_75t_L g1205 ( 
.A1(n_1193),
.A2(n_971),
.B1(n_1043),
.B2(n_964),
.C(n_1023),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1180),
.A2(n_971),
.B1(n_956),
.B2(n_940),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_SL g1207 ( 
.A(n_1182),
.B(n_49),
.C(n_993),
.Y(n_1207)
);

AOI221xp5_ASAP7_75t_L g1208 ( 
.A1(n_1179),
.A2(n_1169),
.B1(n_1171),
.B2(n_1175),
.C(n_1173),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1172),
.B(n_49),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1178),
.A2(n_945),
.B(n_946),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1183),
.A2(n_940),
.B1(n_947),
.B2(n_945),
.C(n_946),
.Y(n_1211)
);

AOI211xp5_ASAP7_75t_L g1212 ( 
.A1(n_1186),
.A2(n_971),
.B(n_947),
.C(n_948),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1176),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1181),
.A2(n_956),
.B1(n_948),
.B2(n_950),
.C(n_940),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1188),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1187),
.B(n_956),
.Y(n_1216)
);

AOI211xp5_ASAP7_75t_L g1217 ( 
.A1(n_1185),
.A2(n_51),
.B(n_52),
.C(n_56),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1203),
.Y(n_1218)
);

NAND4xp75_ASAP7_75t_L g1219 ( 
.A(n_1215),
.B(n_58),
.C(n_59),
.D(n_61),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1200),
.B(n_956),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1204),
.Y(n_1221)
);

NAND4xp75_ASAP7_75t_L g1222 ( 
.A(n_1209),
.B(n_69),
.C(n_70),
.D(n_73),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1216),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1202),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1213),
.B(n_940),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1195),
.A2(n_1217),
.B1(n_1198),
.B2(n_1207),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1199),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1194),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1208),
.B(n_940),
.Y(n_1229)
);

NAND4xp75_ASAP7_75t_L g1230 ( 
.A(n_1196),
.B(n_75),
.C(n_76),
.D(n_77),
.Y(n_1230)
);

XOR2xp5_ASAP7_75t_L g1231 ( 
.A(n_1206),
.B(n_80),
.Y(n_1231)
);

CKINVDCx6p67_ASAP7_75t_R g1232 ( 
.A(n_1201),
.Y(n_1232)
);

NAND4xp75_ASAP7_75t_L g1233 ( 
.A(n_1211),
.B(n_82),
.C(n_83),
.D(n_84),
.Y(n_1233)
);

XNOR2xp5_ASAP7_75t_L g1234 ( 
.A(n_1217),
.B(n_89),
.Y(n_1234)
);

NAND4xp75_ASAP7_75t_L g1235 ( 
.A(n_1210),
.B(n_90),
.C(n_91),
.D(n_94),
.Y(n_1235)
);

NOR2x1_ASAP7_75t_L g1236 ( 
.A(n_1197),
.B(n_431),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1205),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1212),
.B(n_949),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1214),
.Y(n_1239)
);

AOI221xp5_ASAP7_75t_L g1240 ( 
.A1(n_1227),
.A2(n_409),
.B1(n_943),
.B2(n_949),
.C(n_958),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1232),
.A2(n_958),
.B1(n_957),
.B2(n_944),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1218),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1226),
.B(n_431),
.Y(n_1243)
);

OAI211xp5_ASAP7_75t_L g1244 ( 
.A1(n_1226),
.A2(n_95),
.B(n_98),
.C(n_103),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1218),
.B(n_387),
.C(n_957),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1221),
.B(n_928),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1229),
.Y(n_1247)
);

NAND4xp75_ASAP7_75t_L g1248 ( 
.A(n_1228),
.B(n_1237),
.C(n_1236),
.D(n_1223),
.Y(n_1248)
);

OAI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1231),
.A2(n_957),
.B1(n_944),
.B2(n_931),
.C(n_935),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1239),
.A2(n_1224),
.B1(n_1238),
.B2(n_1225),
.Y(n_1250)
);

NOR4xp75_ASAP7_75t_L g1251 ( 
.A(n_1233),
.B(n_104),
.C(n_108),
.D(n_111),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1224),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1220),
.A2(n_944),
.B1(n_930),
.B2(n_928),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1236),
.A2(n_928),
.B1(n_930),
.B2(n_944),
.Y(n_1254)
);

CKINVDCx14_ASAP7_75t_R g1255 ( 
.A(n_1252),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1242),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1251),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1247),
.A2(n_1234),
.B1(n_1230),
.B2(n_1222),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1248),
.Y(n_1259)
);

AND2x2_ASAP7_75t_SL g1260 ( 
.A(n_1246),
.B(n_1240),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1250),
.B(n_1235),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1243),
.Y(n_1262)
);

AOI22x1_ASAP7_75t_L g1263 ( 
.A1(n_1244),
.A2(n_1219),
.B1(n_117),
.B2(n_118),
.Y(n_1263)
);

AOI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1245),
.A2(n_115),
.B(n_119),
.Y(n_1264)
);

XNOR2xp5_ASAP7_75t_L g1265 ( 
.A(n_1241),
.B(n_120),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1254),
.B(n_928),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1249),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1253),
.B(n_121),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1242),
.A2(n_928),
.B1(n_930),
.B2(n_944),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1255),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1256),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1259),
.A2(n_930),
.B1(n_935),
.B2(n_936),
.Y(n_1272)
);

OAI22x1_ASAP7_75t_L g1273 ( 
.A1(n_1263),
.A2(n_1257),
.B1(n_1256),
.B2(n_1261),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1258),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1262),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1267),
.A2(n_930),
.B1(n_937),
.B2(n_936),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1265),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1260),
.A2(n_937),
.B1(n_936),
.B2(n_929),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1268),
.A2(n_937),
.B1(n_936),
.B2(n_939),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1270),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1271),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1275),
.B(n_1264),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1274),
.A2(n_1262),
.B(n_1266),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1277),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1276),
.B(n_1269),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1280),
.A2(n_1273),
.B1(n_1279),
.B2(n_1272),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1281),
.A2(n_1278),
.B1(n_937),
.B2(n_960),
.Y(n_1287)
);

XNOR2xp5_ASAP7_75t_L g1288 ( 
.A(n_1284),
.B(n_1282),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1283),
.B(n_122),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_1289),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1290),
.B(n_1288),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1291),
.A2(n_1285),
.B(n_1287),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1292),
.A2(n_1286),
.B1(n_124),
.B2(n_126),
.Y(n_1293)
);

OAI221xp5_ASAP7_75t_R g1294 ( 
.A1(n_1293),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.C(n_129),
.Y(n_1294)
);

AOI211xp5_ASAP7_75t_L g1295 ( 
.A1(n_1294),
.A2(n_131),
.B(n_135),
.C(n_136),
.Y(n_1295)
);


endmodule