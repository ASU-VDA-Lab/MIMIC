module fake_ariane_1307_n_1268 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1268);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1268;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_209;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_212;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_179;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1257;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_211;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_363;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_63),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_4),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_70),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_97),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_26),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_29),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_34),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_33),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_67),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_93),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_23),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_33),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_94),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_132),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_61),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_69),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_78),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_39),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_44),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_122),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_124),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_11),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_40),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_106),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_119),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_92),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_130),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_80),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_143),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_24),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_26),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_50),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_200),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_222),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_226),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_206),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_179),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_180),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_182),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_184),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_198),
.Y(n_262)
);

BUFx8_ASAP7_75t_SL g263 ( 
.A(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_241),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_263),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_265),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_248),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_251),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_239),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_253),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_252),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_220),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_255),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_241),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_239),
.Y(n_314)
);

BUFx8_ASAP7_75t_SL g315 ( 
.A(n_263),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_249),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_241),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_277),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_303),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_280),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_269),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_288),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_296),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_269),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_284),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_303),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_270),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_272),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_296),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_292),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_267),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_294),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_275),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_312),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_281),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_282),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_291),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_283),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_305),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_285),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_287),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_289),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_295),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_291),
.Y(n_379)
);

BUFx12f_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_291),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_271),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_350),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

CKINVDCx6p67_ASAP7_75t_R g389 ( 
.A(n_366),
.Y(n_389)
);

BUFx12f_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_346),
.B(n_275),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

BUFx12f_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_276),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_276),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_320),
.B(n_278),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_358),
.B(n_278),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_323),
.B(n_302),
.Y(n_404)
);

BUFx8_ASAP7_75t_SL g405 ( 
.A(n_362),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_330),
.B(n_290),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_361),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_319),
.B(n_225),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_325),
.B(n_293),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_360),
.B(n_318),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_360),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_412),
.A2(n_347),
.B1(n_335),
.B2(n_298),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_329),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_372),
.B(n_392),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_371),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_353),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_403),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_411),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_372),
.A2(n_318),
.B1(n_366),
.B2(n_365),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_391),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_370),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_385),
.B(n_364),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_409),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_388),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_385),
.B(n_364),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_393),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

CKINVDCx6p67_ASAP7_75t_R g451 ( 
.A(n_390),
.Y(n_451)
);

BUFx8_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_398),
.B(n_365),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_374),
.A2(n_322),
.B(n_321),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_398),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_373),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_374),
.B(n_337),
.Y(n_462)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_413),
.B(n_337),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_374),
.B(n_338),
.Y(n_467)
);

BUFx8_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_392),
.B(n_321),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_374),
.B(n_338),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_404),
.A2(n_341),
.B1(n_340),
.B2(n_342),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_375),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_394),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_397),
.A2(n_341),
.B1(n_340),
.B2(n_342),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_413),
.A2(n_293),
.B1(n_326),
.B2(n_332),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_376),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_376),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_405),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

NOR2x1_ASAP7_75t_L g484 ( 
.A(n_379),
.B(n_314),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

CKINVDCx6p67_ASAP7_75t_R g487 ( 
.A(n_389),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_370),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_377),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_407),
.B(n_322),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_377),
.Y(n_492)
);

OAI22x1_ASAP7_75t_SL g493 ( 
.A1(n_403),
.A2(n_273),
.B1(n_315),
.B2(n_188),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_379),
.B(n_343),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_370),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_395),
.A2(n_331),
.B1(n_332),
.B2(n_326),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_396),
.B(n_343),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_396),
.B(n_377),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_384),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_400),
.A2(n_273),
.B1(n_315),
.B2(n_187),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_441),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_452),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_499),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_482),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_452),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_454),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_457),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_468),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_432),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_457),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_420),
.B(n_383),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_468),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_476),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_451),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_440),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_458),
.B(n_407),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_487),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_444),
.B(n_407),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_427),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_418),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_418),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_445),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_454),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_433),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_422),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_416),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_435),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_439),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_420),
.B(n_401),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_446),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_419),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_442),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_445),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_455),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_503),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_423),
.B(n_357),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_428),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_455),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_428),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_499),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_493),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_477),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_477),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_430),
.B(n_494),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_463),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_470),
.B(n_202),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_470),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_521),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_516),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_568),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_568),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_570),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_519),
.B(n_424),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_538),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_538),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_528),
.B(n_494),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_535),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_540),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_567),
.B(n_478),
.C(n_479),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_555),
.B(n_465),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_531),
.B(n_483),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_550),
.B(n_465),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_541),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_528),
.B(n_429),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_528),
.B(n_469),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_526),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_542),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_561),
.Y(n_596)
);

INVxp33_ASAP7_75t_SL g597 ( 
.A(n_505),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_547),
.B(n_429),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_542),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_553),
.B(n_469),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_514),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_545),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_526),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_518),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_518),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_545),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_522),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_561),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_581),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_571),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_572),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_576),
.B(n_516),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_572),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_603),
.B(n_449),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_597),
.B(n_505),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_573),
.B(n_523),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_582),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_601),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_581),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_573),
.B(n_508),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_586),
.A2(n_569),
.B1(n_489),
.B2(n_543),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_596),
.B(n_559),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_587),
.B(n_504),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_600),
.B(n_516),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_591),
.A2(n_472),
.B1(n_478),
.B2(n_415),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_598),
.B(n_536),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_L g628 ( 
.A(n_593),
.B(n_472),
.C(n_486),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_571),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_591),
.B(n_525),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_603),
.B(n_463),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_598),
.B(n_509),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_601),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_591),
.A2(n_543),
.B1(n_484),
.B2(n_554),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_571),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_604),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_604),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_577),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_574),
.B(n_508),
.Y(n_639)
);

AND2x2_ASAP7_75t_SL g640 ( 
.A(n_603),
.B(n_449),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_605),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_577),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_577),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_574),
.B(n_516),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_583),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_578),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_583),
.B(n_529),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_605),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_572),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_606),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_598),
.B(n_511),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_603),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_591),
.A2(n_554),
.B1(n_486),
.B2(n_533),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_591),
.B(n_534),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_572),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_580),
.B(n_534),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_589),
.B(n_513),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_578),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_588),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_606),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_572),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_598),
.B(n_517),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_594),
.B(n_529),
.Y(n_664)
);

AO22x1_ASAP7_75t_L g665 ( 
.A1(n_575),
.A2(n_562),
.B1(n_520),
.B2(n_510),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_578),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_579),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_596),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_598),
.B(n_537),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_579),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_596),
.B(n_453),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_607),
.B(n_189),
.C(n_185),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_596),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_608),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_584),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_584),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_584),
.B(n_544),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_608),
.B(n_453),
.C(n_524),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_594),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_585),
.B(n_548),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_608),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_608),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_585),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_585),
.B(n_549),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_590),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_590),
.B(n_534),
.Y(n_687)
);

AO22x2_ASAP7_75t_L g688 ( 
.A1(n_590),
.A2(n_564),
.B1(n_551),
.B2(n_546),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_592),
.B(n_539),
.Y(n_689)
);

INVx8_ASAP7_75t_L g690 ( 
.A(n_592),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_592),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_595),
.A2(n_460),
.B1(n_490),
.B2(n_464),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_595),
.B(n_563),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_617),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_645),
.B(n_595),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_618),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_620),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_619),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_628),
.B(n_463),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_633),
.Y(n_700)
);

XOR2xp5_ASAP7_75t_L g701 ( 
.A(n_665),
.B(n_506),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_609),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_693),
.B(n_659),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_613),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_625),
.A2(n_599),
.B(n_602),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_615),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_636),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_637),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_653),
.B(n_530),
.Y(n_709)
);

XNOR2x2_ASAP7_75t_L g710 ( 
.A(n_628),
.B(n_193),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_641),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_669),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_648),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_650),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_661),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_621),
.B(n_563),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_626),
.B(n_680),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_632),
.B(n_599),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_653),
.B(n_530),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_651),
.B(n_663),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_684),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_626),
.A2(n_501),
.B(n_496),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_681),
.Y(n_724)
);

XOR2x2_ASAP7_75t_L g725 ( 
.A(n_622),
.B(n_506),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_669),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_681),
.Y(n_727)
);

AND2x2_ASAP7_75t_SL g728 ( 
.A(n_640),
.B(n_561),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_651),
.B(n_566),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_639),
.B(n_566),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_685),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_685),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_616),
.Y(n_733)
);

XOR2x2_ASAP7_75t_L g734 ( 
.A(n_634),
.B(n_515),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_663),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_666),
.Y(n_736)
);

XNOR2xp5_ASAP7_75t_L g737 ( 
.A(n_662),
.B(n_515),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_654),
.B(n_532),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_654),
.B(n_599),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_610),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_629),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_635),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_630),
.B(n_602),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_627),
.B(n_532),
.Y(n_744)
);

AND2x2_ASAP7_75t_SL g745 ( 
.A(n_614),
.B(n_602),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_670),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_676),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_638),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_677),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_678),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_627),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_642),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_643),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_646),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_658),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_667),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_673),
.Y(n_757)
);

XOR2xp5_ASAP7_75t_L g758 ( 
.A(n_657),
.B(n_510),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_691),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_688),
.Y(n_760)
);

AOI21x1_ASAP7_75t_L g761 ( 
.A1(n_644),
.A2(n_612),
.B(n_647),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_688),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_686),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_683),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_614),
.B(n_526),
.Y(n_765)
);

INVx4_ASAP7_75t_SL g766 ( 
.A(n_623),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_686),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_613),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_624),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_630),
.B(n_552),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_690),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_613),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_656),
.B(n_552),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_660),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_672),
.B(n_680),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_690),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_656),
.B(n_539),
.Y(n_777)
);

XOR2x2_ASAP7_75t_L g778 ( 
.A(n_672),
.B(n_520),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_671),
.B(n_539),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_664),
.B(n_556),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_721),
.B(n_623),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_775),
.B(n_679),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_696),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_712),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_721),
.B(n_623),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_751),
.B(n_623),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_775),
.B(n_682),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_715),
.B(n_668),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_735),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_715),
.B(n_668),
.Y(n_790)
);

AO221x1_ASAP7_75t_L g791 ( 
.A1(n_704),
.A2(n_652),
.B1(n_660),
.B2(n_682),
.C(n_675),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_764),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_702),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_694),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_769),
.B(n_675),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_698),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_718),
.B(n_196),
.C(n_194),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_706),
.B(n_524),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_729),
.B(n_674),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_699),
.A2(n_631),
.B1(n_689),
.B2(n_687),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_717),
.B(n_682),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_703),
.B(n_660),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_729),
.B(n_649),
.Y(n_803)
);

OAI21xp33_ASAP7_75t_L g804 ( 
.A1(n_718),
.A2(n_186),
.B(n_183),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_744),
.B(n_687),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_712),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_710),
.A2(n_461),
.B1(n_466),
.B2(n_459),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_765),
.A2(n_631),
.B1(n_652),
.B2(n_415),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_730),
.B(n_611),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_733),
.B(n_527),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_697),
.B(n_527),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_700),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_707),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_766),
.B(n_611),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_766),
.B(n_611),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_744),
.B(n_687),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_726),
.B(n_687),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_704),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_699),
.A2(n_631),
.B1(n_689),
.B2(n_526),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_737),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_726),
.B(n_689),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_734),
.A2(n_474),
.B1(n_475),
.B2(n_473),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_708),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_765),
.A2(n_689),
.B1(n_526),
.B2(n_692),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_763),
.B(n_216),
.C(n_197),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_724),
.B(n_649),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_727),
.B(n_655),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_711),
.Y(n_828)
);

NOR2x1p5_ASAP7_75t_L g829 ( 
.A(n_709),
.B(n_655),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_720),
.A2(n_526),
.B1(n_481),
.B2(n_485),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_745),
.B(n_529),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_695),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_738),
.B(n_529),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_758),
.B(n_0),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_731),
.B(n_690),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_713),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_704),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_714),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_701),
.B(n_0),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_768),
.B(n_565),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_768),
.B(n_565),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_723),
.A2(n_557),
.B1(n_558),
.B2(n_556),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_770),
.B(n_565),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_766),
.B(n_565),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_728),
.B(n_556),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_732),
.B(n_1),
.Y(n_846)
);

O2A1O1Ixp5_ASAP7_75t_L g847 ( 
.A1(n_723),
.A2(n_558),
.B(n_560),
.C(n_557),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_750),
.B(n_1),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_740),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_L g850 ( 
.A(n_767),
.B(n_719),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_728),
.B(n_557),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_741),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_716),
.Y(n_853)
);

AO221x1_ASAP7_75t_L g854 ( 
.A1(n_768),
.A2(n_560),
.B1(n_558),
.B2(n_233),
.C(n_225),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_773),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_725),
.A2(n_492),
.B1(n_498),
.B2(n_480),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_792),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_784),
.B(n_736),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_829),
.B(n_722),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_797),
.B(n_782),
.C(n_806),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_784),
.B(n_746),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_781),
.B(n_772),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_818),
.Y(n_863)
);

O2A1O1Ixp5_ASAP7_75t_L g864 ( 
.A1(n_787),
.A2(n_761),
.B(n_780),
.C(n_776),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_SL g865 ( 
.A(n_808),
.B(n_739),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_806),
.B(n_747),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_789),
.B(n_749),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_832),
.B(n_739),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_792),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_797),
.A2(n_778),
.B1(n_777),
.B2(n_780),
.Y(n_870)
);

O2A1O1Ixp5_ASAP7_75t_L g871 ( 
.A1(n_839),
.A2(n_771),
.B(n_779),
.C(n_762),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_802),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_832),
.B(n_795),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_783),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_794),
.Y(n_875)
);

AND2x6_ASAP7_75t_L g876 ( 
.A(n_819),
.B(n_743),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_820),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_785),
.B(n_772),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_804),
.A2(n_760),
.B1(n_743),
.B2(n_754),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_796),
.B(n_772),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_793),
.B(n_779),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_813),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_849),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_812),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_823),
.B(n_774),
.Y(n_885)
);

AND3x1_ASAP7_75t_L g886 ( 
.A(n_834),
.B(n_218),
.C(n_217),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_850),
.B(n_753),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_828),
.B(n_774),
.Y(n_888)
);

O2A1O1Ixp5_ASAP7_75t_L g889 ( 
.A1(n_801),
.A2(n_705),
.B(n_223),
.C(n_228),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_808),
.A2(n_774),
.B(n_507),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_852),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_836),
.B(n_755),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_838),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_853),
.B(n_756),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_788),
.B(n_757),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_790),
.B(n_759),
.Y(n_896)
);

O2A1O1Ixp5_ASAP7_75t_L g897 ( 
.A1(n_809),
.A2(n_224),
.B(n_560),
.C(n_742),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_826),
.B(n_752),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_856),
.A2(n_748),
.B1(n_551),
.B2(n_546),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_827),
.B(n_803),
.Y(n_900)
);

AND2x2_ASAP7_75t_SL g901 ( 
.A(n_805),
.B(n_225),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_855),
.B(n_2),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_817),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_798),
.B(n_810),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_799),
.B(n_2),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_821),
.B(n_3),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_786),
.B(n_3),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_846),
.B(n_4),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_811),
.B(n_5),
.Y(n_909)
);

AND2x2_ASAP7_75t_SL g910 ( 
.A(n_816),
.B(n_230),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_837),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_835),
.B(n_5),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_848),
.B(n_6),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_831),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_831),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_837),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_825),
.B(n_507),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_791),
.B(n_6),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_843),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_800),
.B(n_499),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_856),
.A2(n_448),
.B1(n_450),
.B2(n_186),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_847),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_847),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_830),
.B(n_499),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_833),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_842),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_845),
.B(n_7),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_818),
.Y(n_928)
);

INVx8_ASAP7_75t_L g929 ( 
.A(n_840),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_824),
.B(n_438),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_851),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_814),
.B(n_7),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_815),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_844),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_L g935 ( 
.A(n_807),
.B(n_491),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_822),
.B(n_8),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_935),
.A2(n_822),
.B1(n_807),
.B2(n_854),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_877),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_903),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_886),
.A2(n_841),
.B1(n_195),
.B2(n_215),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_858),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_872),
.B(n_8),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_858),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_863),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_904),
.B(n_9),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_857),
.B(n_9),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_869),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_881),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_861),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_863),
.B(n_10),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_909),
.B(n_10),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_861),
.B(n_11),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_860),
.A2(n_208),
.B(n_195),
.C(n_190),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_859),
.B(n_933),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_866),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_866),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_871),
.A2(n_190),
.B(n_233),
.C(n_230),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_872),
.B(n_12),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_867),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_859),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_873),
.B(n_12),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_893),
.B(n_13),
.Y(n_962)
);

CKINVDCx8_ASAP7_75t_R g963 ( 
.A(n_934),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_895),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_928),
.Y(n_965)
);

CKINVDCx11_ASAP7_75t_R g966 ( 
.A(n_929),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_887),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_887),
.Y(n_968)
);

BUFx2_ASAP7_75t_SL g969 ( 
.A(n_902),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_875),
.Y(n_970)
);

BUFx4f_ASAP7_75t_L g971 ( 
.A(n_901),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_867),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_929),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_925),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_911),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_884),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_936),
.A2(n_865),
.B1(n_930),
.B2(n_926),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_918),
.Y(n_978)
);

CKINVDCx8_ASAP7_75t_R g979 ( 
.A(n_929),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_910),
.B(n_438),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_905),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_892),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_865),
.A2(n_437),
.B1(n_500),
.B2(n_204),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_894),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_876),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_874),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_931),
.B(n_13),
.Y(n_987)
);

AOI211xp5_ASAP7_75t_L g988 ( 
.A1(n_918),
.A2(n_233),
.B(n_230),
.C(n_16),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_913),
.B(n_14),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_922),
.B(n_14),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_906),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_896),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_907),
.Y(n_993)
);

INVxp33_ASAP7_75t_SL g994 ( 
.A(n_938),
.Y(n_994)
);

AO21x1_ASAP7_75t_L g995 ( 
.A1(n_945),
.A2(n_913),
.B(n_908),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_978),
.B(n_898),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_977),
.A2(n_870),
.B1(n_900),
.B2(n_878),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_970),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_988),
.A2(n_908),
.B(n_917),
.C(n_889),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_990),
.A2(n_912),
.B(n_923),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_971),
.A2(n_991),
.B1(n_993),
.B2(n_985),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_966),
.B(n_912),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_944),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_985),
.B(n_914),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_939),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_971),
.A2(n_862),
.B(n_924),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_956),
.B(n_919),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_L g1008 ( 
.A(n_985),
.B(n_916),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_959),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_948),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_953),
.A2(n_951),
.B(n_989),
.C(n_993),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_957),
.A2(n_953),
.B(n_990),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_963),
.B(n_932),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_985),
.B(n_868),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_991),
.A2(n_920),
.B1(n_915),
.B2(n_927),
.Y(n_1015)
);

INVx3_ASAP7_75t_SL g1016 ( 
.A(n_944),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_944),
.B(n_864),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_952),
.A2(n_890),
.B(n_885),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_979),
.B(n_876),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_981),
.B(n_880),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_952),
.A2(n_888),
.B(n_897),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_969),
.A2(n_879),
.B1(n_899),
.B2(n_921),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_968),
.A2(n_882),
.B(n_883),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_968),
.A2(n_891),
.B(n_876),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_954),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_955),
.B(n_876),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_962),
.A2(n_233),
.B1(n_230),
.B2(n_209),
.C(n_210),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_954),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_987),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_967),
.A2(n_204),
.B1(n_434),
.B2(n_426),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_937),
.A2(n_204),
.B1(n_437),
.B2(n_500),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_980),
.A2(n_467),
.B(n_462),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_972),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_986),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_962),
.A2(n_306),
.B(n_297),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_950),
.A2(n_201),
.B(n_207),
.C(n_211),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_L g1037 ( 
.A1(n_992),
.A2(n_497),
.B(n_471),
.C(n_467),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_941),
.A2(n_949),
.B(n_943),
.Y(n_1038)
);

OR2x6_ASAP7_75t_L g1039 ( 
.A(n_973),
.B(n_438),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_982),
.B(n_204),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_961),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_964),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_975),
.B(n_15),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_984),
.A2(n_471),
.B(n_462),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_965),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_947),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_946),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_976),
.B(n_204),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_942),
.B(n_204),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_987),
.A2(n_960),
.B(n_983),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_960),
.A2(n_497),
.B(n_501),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_958),
.A2(n_974),
.B(n_940),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_978),
.B(n_204),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_979),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_985),
.B(n_18),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_971),
.A2(n_488),
.B(n_443),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_938),
.B(n_19),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_978),
.B(n_20),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_938),
.B(n_20),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_995),
.B(n_21),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1025),
.B(n_21),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1000),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1025),
.B(n_22),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1048),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1028),
.B(n_22),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_1028),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1042),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_996),
.B(n_23),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_1010),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_998),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1005),
.B(n_24),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_1009),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_1011),
.A2(n_212),
.B(n_214),
.C(n_219),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1038),
.B(n_25),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1040),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1003),
.B(n_25),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_994),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_1054),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_999),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1054),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_1041),
.A2(n_221),
.B(n_227),
.C(n_231),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1066),
.A2(n_1023),
.B(n_1001),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1072),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1060),
.B(n_1053),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1066),
.A2(n_1024),
.B(n_1052),
.Y(n_1085)
);

NAND3xp33_ASAP7_75t_SL g1086 ( 
.A(n_1079),
.B(n_1017),
.C(n_1047),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1074),
.A2(n_1012),
.B(n_1058),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1066),
.A2(n_1018),
.B(n_1026),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1080),
.A2(n_1045),
.B1(n_1029),
.B2(n_1046),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1078),
.B(n_1016),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1078),
.B(n_1033),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1062),
.A2(n_1050),
.B(n_1034),
.Y(n_1092)
);

OAI211xp5_ASAP7_75t_SL g1093 ( 
.A1(n_1071),
.A2(n_1059),
.B(n_1057),
.C(n_1036),
.Y(n_1093)
);

OAI21xp33_ASAP7_75t_L g1094 ( 
.A1(n_1073),
.A2(n_1043),
.B(n_1031),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1073),
.A2(n_1049),
.B(n_1019),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1069),
.B(n_1002),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1062),
.A2(n_1013),
.B(n_1021),
.C(n_1027),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_1075),
.A2(n_1015),
.B(n_1055),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1068),
.A2(n_997),
.B(n_1006),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1063),
.B(n_1029),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_1077),
.B(n_1029),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_SL g1102 ( 
.A1(n_1061),
.A2(n_1055),
.B(n_1008),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1063),
.B(n_1007),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1081),
.A2(n_1037),
.B(n_1022),
.Y(n_1104)
);

INVx6_ASAP7_75t_L g1105 ( 
.A(n_1061),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1061),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1065),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1107),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_1107),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1083),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1086),
.A2(n_1014),
.B1(n_1064),
.B2(n_1067),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1087),
.B(n_1070),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_1096),
.B(n_1065),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1104),
.B(n_1065),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_1113),
.B(n_1101),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1109),
.Y(n_1116)
);

INVx5_ASAP7_75t_L g1117 ( 
.A(n_1116),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1115),
.B(n_1105),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1117),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_1118),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_SL g1121 ( 
.A1(n_1120),
.A2(n_1114),
.B1(n_1112),
.B2(n_1109),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1120),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1122),
.A2(n_1119),
.B(n_1108),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1121),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1124),
.A2(n_1084),
.B1(n_1111),
.B2(n_1092),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1124),
.A2(n_1094),
.B1(n_1107),
.B2(n_1110),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1123),
.B(n_1106),
.Y(n_1127)
);

INVx11_ASAP7_75t_L g1128 ( 
.A(n_1127),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1126),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1125),
.A2(n_1090),
.B(n_1097),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1129),
.A2(n_1099),
.B(n_1088),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1128),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1131),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_1134),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1133),
.B(n_1130),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1135),
.B(n_1105),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1136),
.B(n_1094),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_1137),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1138),
.B(n_1100),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_1139),
.B(n_1089),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_1140),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1142),
.B(n_1091),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_1141),
.B(n_27),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1142),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1145),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_1143),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_1082),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1147),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1146),
.Y(n_1150)
);

XOR2x1_ASAP7_75t_L g1151 ( 
.A(n_1150),
.B(n_1148),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1149),
.B(n_1085),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_1076),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1153),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1154),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1155),
.B(n_28),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1156),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1158),
.B(n_30),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1157),
.B(n_30),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1160),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1159),
.A2(n_1093),
.B1(n_1103),
.B2(n_1076),
.Y(n_1162)
);

AOI221xp5_ASAP7_75t_L g1163 ( 
.A1(n_1160),
.A2(n_236),
.B1(n_1098),
.B2(n_1102),
.C(n_286),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1161),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1162),
.B(n_1020),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1163),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1164),
.B(n_31),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1166),
.A2(n_1095),
.B1(n_1081),
.B2(n_31),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1167),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1168),
.B(n_1165),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1169),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1170),
.Y(n_1172)
);

AOI211xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1172),
.A2(n_297),
.B(n_306),
.C(n_32),
.Y(n_1173)
);

OAI211xp5_ASAP7_75t_L g1174 ( 
.A1(n_1171),
.A2(n_286),
.B(n_32),
.C(n_339),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1173),
.A2(n_286),
.B(n_324),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1174),
.B(n_359),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1176),
.Y(n_1177)
);

O2A1O1Ixp5_ASAP7_75t_SL g1178 ( 
.A1(n_1175),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1178)
);

NAND4xp75_ASAP7_75t_L g1179 ( 
.A(n_1177),
.B(n_1178),
.C(n_363),
.D(n_359),
.Y(n_1179)
);

XOR2x2_ASAP7_75t_L g1180 ( 
.A(n_1177),
.B(n_38),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_L g1181 ( 
.A(n_1177),
.B(n_363),
.C(n_1056),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1180),
.B(n_1179),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1181),
.A2(n_363),
.B(n_1039),
.Y(n_1183)
);

NOR3x1_ASAP7_75t_L g1184 ( 
.A(n_1179),
.B(n_41),
.C(n_42),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1182),
.B(n_1184),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_L g1186 ( 
.A(n_1183),
.B(n_1039),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1185),
.Y(n_1187)
);

NAND2xp33_ASAP7_75t_L g1188 ( 
.A(n_1186),
.B(n_410),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1187),
.B(n_43),
.Y(n_1189)
);

NOR2x1_ASAP7_75t_L g1190 ( 
.A(n_1188),
.B(n_1004),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1189),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1190),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1192),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_L g1194 ( 
.A(n_1191),
.B(n_45),
.C(n_46),
.Y(n_1194)
);

NOR3xp33_ASAP7_75t_L g1195 ( 
.A(n_1193),
.B(n_1004),
.C(n_48),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1194),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1196),
.B(n_47),
.Y(n_1197)
);

NOR4xp25_ASAP7_75t_L g1198 ( 
.A(n_1195),
.B(n_49),
.C(n_51),
.D(n_52),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_L g1199 ( 
.A(n_1196),
.B(n_53),
.C(n_54),
.Y(n_1199)
);

NAND4xp25_ASAP7_75t_L g1200 ( 
.A(n_1198),
.B(n_55),
.C(n_56),
.D(n_57),
.Y(n_1200)
);

AND3x1_ASAP7_75t_L g1201 ( 
.A(n_1197),
.B(n_1199),
.C(n_59),
.Y(n_1201)
);

OR4x2_ASAP7_75t_L g1202 ( 
.A(n_1198),
.B(n_58),
.C(n_60),
.D(n_62),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1201),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1202),
.Y(n_1204)
);

OAI22x1_ASAP7_75t_L g1205 ( 
.A1(n_1203),
.A2(n_1200),
.B1(n_65),
.B2(n_66),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1204),
.B(n_64),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1205),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1206),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1208),
.A2(n_79),
.B(n_81),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1207),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1210),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_SL g1212 ( 
.A(n_1209),
.B(n_82),
.C(n_84),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_L g1213 ( 
.A(n_1211),
.B(n_85),
.Y(n_1213)
);

XNOR2xp5_ASAP7_75t_L g1214 ( 
.A(n_1212),
.B(n_86),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1213),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1214),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1213),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_1217)
);

XNOR2x1_ASAP7_75t_L g1218 ( 
.A(n_1216),
.B(n_90),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1215),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1217),
.Y(n_1220)
);

AOI21xp33_ASAP7_75t_L g1221 ( 
.A1(n_1219),
.A2(n_91),
.B(n_96),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1218),
.Y(n_1222)
);

AOI222xp33_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_1220),
.B1(n_99),
.B2(n_100),
.C1(n_101),
.C2(n_103),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1221),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1222),
.A2(n_98),
.B1(n_104),
.B2(n_105),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1224),
.A2(n_1223),
.B(n_1225),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1224),
.B(n_107),
.Y(n_1227)
);

XNOR2xp5_ASAP7_75t_L g1228 ( 
.A(n_1224),
.B(n_108),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1226),
.B(n_109),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1227),
.A2(n_110),
.B(n_112),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1228),
.A2(n_113),
.B(n_115),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1229),
.A2(n_1230),
.B1(n_1231),
.B2(n_118),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1229),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_1233)
);

AO22x2_ASAP7_75t_L g1234 ( 
.A1(n_1229),
.A2(n_123),
.B1(n_126),
.B2(n_129),
.Y(n_1234)
);

AO22x2_ASAP7_75t_L g1235 ( 
.A1(n_1229),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1229),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1229),
.A2(n_139),
.B1(n_140),
.B2(n_145),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1229),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1229),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1229),
.A2(n_156),
.B(n_157),
.Y(n_1240)
);

AO22x2_ASAP7_75t_L g1241 ( 
.A1(n_1229),
.A2(n_158),
.B1(n_160),
.B2(n_162),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1229),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1229),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_1243)
);

AO22x2_ASAP7_75t_L g1244 ( 
.A1(n_1229),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_1244)
);

AOI222xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1240),
.A2(n_176),
.B1(n_177),
.B2(n_1035),
.C1(n_1030),
.C2(n_410),
.Y(n_1245)
);

AOI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_1233),
.A2(n_1051),
.B(n_1032),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1236),
.A2(n_1044),
.B1(n_443),
.B2(n_502),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1237),
.A2(n_502),
.B1(n_443),
.B2(n_488),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1238),
.A2(n_410),
.B(n_491),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1243),
.A2(n_502),
.B(n_488),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1239),
.A2(n_410),
.B(n_491),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1234),
.A2(n_502),
.B1(n_443),
.B2(n_488),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1244),
.A2(n_410),
.B(n_491),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1246),
.B(n_1235),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1249),
.A2(n_1241),
.B(n_1232),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1253),
.A2(n_1242),
.B(n_495),
.Y(n_1256)
);

XNOR2xp5_ASAP7_75t_L g1257 ( 
.A(n_1251),
.B(n_410),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1247),
.B(n_495),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1250),
.Y(n_1259)
);

OAI221xp5_ASAP7_75t_R g1260 ( 
.A1(n_1259),
.A2(n_1245),
.B1(n_1248),
.B2(n_1252),
.C(n_410),
.Y(n_1260)
);

AOI322xp5_ASAP7_75t_L g1261 ( 
.A1(n_1255),
.A2(n_495),
.A3(n_410),
.B1(n_381),
.B2(n_382),
.C1(n_378),
.C2(n_386),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1254),
.A2(n_491),
.B1(n_495),
.B2(n_381),
.Y(n_1262)
);

OAI32xp33_ASAP7_75t_L g1263 ( 
.A1(n_1260),
.A2(n_1257),
.A3(n_1258),
.B1(n_1256),
.B2(n_382),
.Y(n_1263)
);

AOI221xp5_ASAP7_75t_L g1264 ( 
.A1(n_1263),
.A2(n_1262),
.B1(n_1261),
.B2(n_381),
.C(n_382),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1264),
.A2(n_378),
.B(n_381),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1265),
.A2(n_378),
.B1(n_381),
.B2(n_382),
.Y(n_1266)
);

AOI211xp5_ASAP7_75t_L g1267 ( 
.A1(n_1266),
.A2(n_384),
.B(n_456),
.C(n_381),
.Y(n_1267)
);

AOI211xp5_ASAP7_75t_L g1268 ( 
.A1(n_1267),
.A2(n_384),
.B(n_378),
.C(n_381),
.Y(n_1268)
);


endmodule