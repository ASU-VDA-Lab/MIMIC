module fake_jpeg_21332_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_17),
.B1(n_32),
.B2(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_40),
.B1(n_36),
.B2(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_17),
.B1(n_32),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_55),
.B1(n_42),
.B2(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_17),
.B1(n_19),
.B2(n_30),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_35),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_69),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_36),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_61),
.A2(n_62),
.B1(n_85),
.B2(n_92),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_18),
.B1(n_22),
.B2(n_30),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_60),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_70),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_18),
.B1(n_30),
.B2(n_19),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_75),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_77),
.Y(n_122)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_78),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_91),
.B1(n_21),
.B2(n_31),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_56),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_88),
.C(n_37),
.Y(n_119)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_18),
.B1(n_36),
.B2(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_94),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_43),
.B1(n_42),
.B2(n_38),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_36),
.B1(n_20),
.B2(n_31),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_42),
.B(n_43),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_61),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_46),
.B(n_38),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_117),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_42),
.B(n_43),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_111),
.B(n_119),
.C(n_75),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_59),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_94),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_37),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_34),
.C(n_35),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_80),
.B1(n_82),
.B2(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_37),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_89),
.B1(n_74),
.B2(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_73),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_93),
.B1(n_65),
.B2(n_95),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_131),
.B1(n_133),
.B2(n_136),
.Y(n_173)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_135),
.Y(n_154)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_79),
.B1(n_87),
.B2(n_64),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_83),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_88),
.B1(n_84),
.B2(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_148),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_111),
.B(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_144),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_117),
.C(n_125),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_146),
.C(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_33),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_152),
.B1(n_153),
.B2(n_140),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_73),
.C(n_34),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_33),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_33),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_77),
.B1(n_35),
.B2(n_37),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_119),
.B1(n_101),
.B2(n_104),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_90),
.B1(n_67),
.B2(n_70),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_35),
.B1(n_71),
.B2(n_73),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_163),
.B1(n_165),
.B2(n_179),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_175),
.C(n_183),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_123),
.B(n_105),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_160),
.A2(n_164),
.B(n_184),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_108),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_121),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_105),
.B1(n_109),
.B2(n_113),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_108),
.B1(n_98),
.B2(n_122),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_96),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_169),
.B(n_171),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_112),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_122),
.B(n_106),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_178),
.B(n_26),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_114),
.C(n_98),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_176),
.B(n_132),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_178),
.B1(n_173),
.B2(n_174),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_101),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_111),
.B1(n_124),
.B2(n_110),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_111),
.B1(n_97),
.B2(n_110),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_182),
.B1(n_185),
.B2(n_1),
.Y(n_216)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_133),
.A2(n_97),
.B1(n_21),
.B2(n_25),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_151),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_33),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_118),
.B(n_97),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_121),
.B1(n_102),
.B2(n_21),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_191),
.B1(n_195),
.B2(n_185),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_173),
.A2(n_145),
.B1(n_136),
.B2(n_129),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_127),
.B1(n_102),
.B2(n_25),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_167),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_197),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_206),
.C(n_210),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_28),
.B(n_33),
.Y(n_202)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_186),
.B(n_28),
.Y(n_234)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_163),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_23),
.C(n_29),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_25),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_211),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_23),
.C(n_29),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_27),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_154),
.B(n_16),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_33),
.Y(n_214)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_29),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_29),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_23),
.C(n_27),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_156),
.C(n_179),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_239),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_168),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_222),
.B(n_195),
.C(n_199),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_188),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_241),
.C(n_218),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_216),
.B1(n_199),
.B2(n_215),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_172),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_238),
.Y(n_251)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_196),
.B(n_200),
.Y(n_254)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_176),
.B1(n_168),
.B2(n_162),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_200),
.B(n_203),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_155),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_155),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_157),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_247),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_206),
.C(n_210),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_249),
.C(n_261),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_238),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_226),
.C(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_192),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_23),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_189),
.B1(n_191),
.B2(n_211),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_227),
.B1(n_230),
.B2(n_225),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_231),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_254),
.B(n_256),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_237),
.B1(n_232),
.B2(n_220),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_217),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_260),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_242),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_201),
.C(n_157),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_262),
.A2(n_240),
.B(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_272),
.B1(n_2),
.B2(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_193),
.C(n_196),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_279),
.C(n_14),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_272)
);

A2O1A1O1Ixp25_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_28),
.B(n_23),
.C(n_10),
.D(n_11),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_10),
.C(n_15),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_258),
.B1(n_254),
.B2(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_12),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_2),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_246),
.B(n_247),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_14),
.C(n_13),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_251),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_281),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_244),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_291),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_251),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_14),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_273),
.B1(n_264),
.B2(n_266),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_263),
.C(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_269),
.C(n_268),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_267),
.Y(n_300)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_275),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_13),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_283),
.B1(n_272),
.B2(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_310),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_289),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_295),
.C(n_298),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_264),
.B(n_278),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_282),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_13),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_302),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_301),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_312),
.B(n_309),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_320),
.B(n_321),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_307),
.B(n_305),
.C(n_296),
.Y(n_320)
);

AOI221xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_316),
.B1(n_318),
.B2(n_5),
.C(n_6),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_3),
.B(n_4),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_3),
.C(n_4),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_326)
);


endmodule