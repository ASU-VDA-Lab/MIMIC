module fake_jpeg_13695_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_9),
.B(n_12),
.Y(n_27)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_13),
.B(n_16),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_31),
.C(n_17),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_22),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_36),
.B1(n_23),
.B2(n_25),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_31),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B(n_13),
.Y(n_45)
);

FAx1_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_6),
.CI(n_7),
.CON(n_43),
.SN(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_42),
.C(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_37),
.B1(n_33),
.B2(n_16),
.Y(n_46)
);

XNOR2x1_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_43),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_50),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

AOI322xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_52),
.A3(n_44),
.B1(n_6),
.B2(n_35),
.C1(n_41),
.C2(n_17),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_44),
.Y(n_55)
);


endmodule