module real_aes_7910_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g500 ( .A(n_1), .Y(n_500) );
INVx1_ASAP7_75t_L g206 ( .A(n_2), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_3), .A2(n_38), .B1(n_167), .B2(n_530), .Y(n_545) );
AOI21xp33_ASAP7_75t_L g174 ( .A1(n_4), .A2(n_148), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_5), .B(n_141), .Y(n_513) );
AND2x6_ASAP7_75t_L g153 ( .A(n_6), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_7), .A2(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_8), .B(n_39), .Y(n_465) );
INVx1_ASAP7_75t_L g181 ( .A(n_9), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_10), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g146 ( .A(n_11), .Y(n_146) );
INVx1_ASAP7_75t_L g494 ( .A(n_12), .Y(n_494) );
INVx1_ASAP7_75t_L g262 ( .A(n_13), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_14), .B(n_189), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_15), .A2(n_105), .B1(n_116), .B2(n_779), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_16), .B(n_142), .Y(n_571) );
AO32x2_ASAP7_75t_L g543 ( .A1(n_17), .A2(n_141), .A3(n_186), .B1(n_522), .B2(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_18), .A2(n_63), .B1(n_130), .B2(n_131), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_18), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_19), .B(n_167), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_20), .B(n_162), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_21), .B(n_142), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_22), .A2(n_51), .B1(n_167), .B2(n_530), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_23), .B(n_148), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_24), .A2(n_80), .B1(n_167), .B2(n_189), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_25), .B(n_167), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_26), .B(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_27), .A2(n_260), .B(n_261), .C(n_263), .Y(n_259) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_29), .B(n_183), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_30), .B(n_179), .Y(n_208) );
INVx1_ASAP7_75t_L g195 ( .A(n_31), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_32), .A2(n_33), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_32), .Y(n_125) );
INVxp67_ASAP7_75t_L g124 ( .A(n_33), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_33), .B(n_183), .Y(n_560) );
INVx2_ASAP7_75t_L g151 ( .A(n_34), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_35), .B(n_167), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_36), .B(n_183), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_37), .A2(n_153), .B(n_157), .C(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g193 ( .A(n_40), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_41), .A2(n_473), .B1(n_476), .B2(n_477), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_41), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_42), .B(n_179), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_43), .B(n_167), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_44), .A2(n_90), .B1(n_225), .B2(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_45), .B(n_167), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_46), .B(n_167), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_47), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_48), .A2(n_70), .B1(n_474), .B2(n_475), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_48), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_49), .B(n_499), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_50), .B(n_148), .Y(n_250) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_52), .A2(n_61), .B1(n_167), .B2(n_189), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_53), .A2(n_157), .B1(n_189), .B2(n_191), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_54), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_55), .B(n_167), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_56), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_57), .B(n_167), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_58), .A2(n_166), .B(n_178), .C(n_180), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_59), .Y(n_238) );
INVx1_ASAP7_75t_L g176 ( .A(n_60), .Y(n_176) );
INVx1_ASAP7_75t_L g154 ( .A(n_62), .Y(n_154) );
INVx1_ASAP7_75t_L g130 ( .A(n_63), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_64), .B(n_167), .Y(n_501) );
INVx1_ASAP7_75t_L g145 ( .A(n_65), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
AO32x2_ASAP7_75t_L g527 ( .A1(n_67), .A2(n_141), .A3(n_242), .B1(n_522), .B2(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g520 ( .A(n_68), .Y(n_520) );
INVx1_ASAP7_75t_L g555 ( .A(n_69), .Y(n_555) );
INVx1_ASAP7_75t_L g474 ( .A(n_70), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_SL g161 ( .A1(n_71), .A2(n_162), .B(n_163), .C(n_166), .Y(n_161) );
INVxp67_ASAP7_75t_L g164 ( .A(n_72), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_73), .B(n_189), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_74), .A2(n_471), .B1(n_472), .B2(n_478), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_74), .Y(n_471) );
INVx1_ASAP7_75t_L g115 ( .A(n_75), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_76), .B(n_461), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_77), .A2(n_463), .B1(n_469), .B2(n_774), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_78), .Y(n_199) );
INVx1_ASAP7_75t_L g231 ( .A(n_79), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_81), .A2(n_153), .B(n_157), .C(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_82), .B(n_530), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_83), .B(n_189), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_84), .B(n_207), .Y(n_221) );
INVx2_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_86), .B(n_162), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_87), .B(n_189), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_88), .A2(n_153), .B(n_157), .C(n_205), .Y(n_204) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_89), .B(n_112), .C(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g462 ( .A(n_89), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g480 ( .A(n_89), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_91), .A2(n_103), .B1(n_189), .B2(n_190), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_92), .B(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_93), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_94), .A2(n_153), .B(n_157), .C(n_245), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_95), .Y(n_252) );
INVx1_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_97), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_98), .B(n_207), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_99), .B(n_189), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_100), .B(n_141), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_101), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_102), .A2(n_148), .B(n_155), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx5_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_108), .Y(n_780) );
OR2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g464 ( .A(n_112), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_467), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g778 ( .A(n_120), .Y(n_778) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_459), .B(n_466), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B1(n_127), .B2(n_458), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_123), .Y(n_458) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_132), .B2(n_457), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g457 ( .A(n_132), .Y(n_457) );
AOI22xp5_ASAP7_75t_SL g479 ( .A1(n_132), .A2(n_480), .B1(n_481), .B2(n_773), .Y(n_479) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND4x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_375), .C(n_422), .D(n_442), .Y(n_133) );
NOR3xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_305), .C(n_330), .Y(n_134) );
OAI211xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_213), .B(n_265), .C(n_295), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_184), .Y(n_137) );
INVx3_ASAP7_75t_SL g347 ( .A(n_138), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_138), .B(n_278), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_138), .B(n_200), .Y(n_428) );
AND2x2_ASAP7_75t_L g451 ( .A(n_138), .B(n_317), .Y(n_451) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_172), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g269 ( .A(n_140), .B(n_173), .Y(n_269) );
INVx3_ASAP7_75t_L g282 ( .A(n_140), .Y(n_282) );
AND2x2_ASAP7_75t_L g287 ( .A(n_140), .B(n_172), .Y(n_287) );
OR2x2_ASAP7_75t_L g338 ( .A(n_140), .B(n_279), .Y(n_338) );
BUFx2_ASAP7_75t_L g358 ( .A(n_140), .Y(n_358) );
AND2x2_ASAP7_75t_L g368 ( .A(n_140), .B(n_279), .Y(n_368) );
AND2x2_ASAP7_75t_L g374 ( .A(n_140), .B(n_185), .Y(n_374) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_147), .B(n_169), .Y(n_140) );
INVx4_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_141), .A2(n_506), .B(n_513), .Y(n_505) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_143), .B(n_144), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx2_ASAP7_75t_L g256 ( .A(n_148), .Y(n_256) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_149), .B(n_153), .Y(n_197) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g499 ( .A(n_150), .Y(n_499) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
INVx1_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
INVx1_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
INVx1_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
INVx3_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx4_ASAP7_75t_SL g168 ( .A(n_153), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_153), .A2(n_493), .B(n_497), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_153), .A2(n_507), .B(n_510), .Y(n_506) );
BUFx3_ASAP7_75t_L g522 ( .A(n_153), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_153), .A2(n_535), .B(n_539), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_153), .A2(n_554), .B(n_557), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_160), .B(n_161), .C(n_168), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_156), .A2(n_168), .B(n_176), .C(n_177), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_156), .A2(n_168), .B(n_258), .C(n_259), .Y(n_257) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
BUFx3_ASAP7_75t_L g225 ( .A(n_158), .Y(n_225) );
INVx1_ASAP7_75t_L g530 ( .A(n_158), .Y(n_530) );
INVx1_ASAP7_75t_L g538 ( .A(n_162), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_165), .B(n_181), .Y(n_180) );
INVx5_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
OAI22xp5_ASAP7_75t_SL g528 ( .A1(n_165), .A2(n_179), .B1(n_529), .B2(n_531), .Y(n_528) );
O2A1O1Ixp5_ASAP7_75t_SL g554 ( .A1(n_166), .A2(n_207), .B(n_555), .C(n_556), .Y(n_554) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_167), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_168), .A2(n_188), .B1(n_196), .B2(n_197), .Y(n_187) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_170), .A2(n_174), .B(n_182), .Y(n_173) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g227 ( .A(n_171), .B(n_228), .Y(n_227) );
AO21x1_ASAP7_75t_L g566 ( .A1(n_171), .A2(n_567), .B(n_570), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_171), .B(n_522), .C(n_567), .Y(n_585) );
INVx1_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_173), .B(n_279), .Y(n_293) );
INVx2_ASAP7_75t_L g303 ( .A(n_173), .Y(n_303) );
AND2x2_ASAP7_75t_L g316 ( .A(n_173), .B(n_282), .Y(n_316) );
OR2x2_ASAP7_75t_L g327 ( .A(n_173), .B(n_279), .Y(n_327) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_173), .B(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g385 ( .A(n_173), .Y(n_385) );
AND2x2_ASAP7_75t_L g431 ( .A(n_173), .B(n_185), .Y(n_431) );
O2A1O1Ixp5_ASAP7_75t_L g519 ( .A1(n_178), .A2(n_498), .B(n_520), .C(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_178), .A2(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g248 ( .A(n_179), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_179), .A2(n_502), .B1(n_545), .B2(n_546), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_179), .A2(n_502), .B1(n_568), .B2(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g212 ( .A(n_183), .Y(n_212) );
INVx2_ASAP7_75t_L g242 ( .A(n_183), .Y(n_242) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_183), .A2(n_255), .B(n_264), .Y(n_254) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_183), .A2(n_534), .B(n_542), .Y(n_533) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_183), .A2(n_553), .B(n_560), .Y(n_552) );
INVx3_ASAP7_75t_SL g304 ( .A(n_184), .Y(n_304) );
OR2x2_ASAP7_75t_L g357 ( .A(n_184), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
INVx3_ASAP7_75t_L g279 ( .A(n_185), .Y(n_279) );
AND2x2_ASAP7_75t_L g346 ( .A(n_185), .B(n_201), .Y(n_346) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_185), .Y(n_414) );
AOI33xp33_ASAP7_75t_L g418 ( .A1(n_185), .A2(n_347), .A3(n_354), .B1(n_363), .B2(n_419), .B3(n_420), .Y(n_418) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_198), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_186), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_186), .A2(n_202), .B(n_210), .Y(n_201) );
INVx2_ASAP7_75t_L g226 ( .A(n_186), .Y(n_226) );
INVx2_ASAP7_75t_L g209 ( .A(n_189), .Y(n_209) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g191 ( .A1(n_192), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_191) );
INVx2_ASAP7_75t_L g194 ( .A(n_192), .Y(n_194) );
INVx4_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_197), .A2(n_203), .B(n_204), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_197), .A2(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g267 ( .A(n_200), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_200), .B(n_282), .Y(n_281) );
NOR3xp33_ASAP7_75t_L g341 ( .A(n_200), .B(n_342), .C(n_344), .Y(n_341) );
AND2x2_ASAP7_75t_L g367 ( .A(n_200), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_200), .B(n_374), .Y(n_377) );
AND2x2_ASAP7_75t_L g430 ( .A(n_200), .B(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g286 ( .A(n_201), .Y(n_286) );
OR2x2_ASAP7_75t_L g380 ( .A(n_201), .B(n_279), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .C(n_209), .Y(n_205) );
INVx2_ASAP7_75t_L g502 ( .A(n_207), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_207), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_207), .A2(n_517), .B(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_209), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_212), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_212), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_239), .Y(n_213) );
AOI32xp33_ASAP7_75t_L g331 ( .A1(n_214), .A2(n_332), .A3(n_334), .B1(n_336), .B2(n_339), .Y(n_331) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_214), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g434 ( .A(n_214), .Y(n_434) );
INVx4_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g366 ( .A(n_215), .B(n_350), .Y(n_366) );
AND2x2_ASAP7_75t_L g386 ( .A(n_215), .B(n_312), .Y(n_386) );
AND2x2_ASAP7_75t_L g454 ( .A(n_215), .B(n_372), .Y(n_454) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_229), .Y(n_215) );
INVx3_ASAP7_75t_L g275 ( .A(n_216), .Y(n_275) );
AND2x2_ASAP7_75t_L g289 ( .A(n_216), .B(n_273), .Y(n_289) );
OR2x2_ASAP7_75t_L g294 ( .A(n_216), .B(n_272), .Y(n_294) );
INVx1_ASAP7_75t_L g301 ( .A(n_216), .Y(n_301) );
AND2x2_ASAP7_75t_L g309 ( .A(n_216), .B(n_283), .Y(n_309) );
AND2x2_ASAP7_75t_L g311 ( .A(n_216), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_216), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g364 ( .A(n_216), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_216), .B(n_449), .Y(n_448) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
AOI21xp5_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_219), .B(n_226), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_223), .A2(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g263 ( .A(n_225), .Y(n_263) );
INVx1_ASAP7_75t_L g236 ( .A(n_226), .Y(n_236) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_226), .A2(n_492), .B(n_503), .Y(n_491) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_226), .A2(n_515), .B(n_523), .Y(n_514) );
INVx2_ASAP7_75t_L g273 ( .A(n_229), .Y(n_273) );
AND2x2_ASAP7_75t_L g319 ( .A(n_229), .B(n_240), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_229), .B(n_254), .Y(n_329) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_236), .B(n_237), .Y(n_229) );
INVx2_ASAP7_75t_L g449 ( .A(n_239), .Y(n_449) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_253), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_240), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g290 ( .A(n_240), .Y(n_290) );
AND2x2_ASAP7_75t_L g334 ( .A(n_240), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g350 ( .A(n_240), .B(n_313), .Y(n_350) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g298 ( .A(n_241), .Y(n_298) );
AND2x2_ASAP7_75t_L g312 ( .A(n_241), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g363 ( .A(n_241), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_241), .B(n_273), .Y(n_395) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_251), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_250), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_249), .Y(n_245) );
AND2x2_ASAP7_75t_L g274 ( .A(n_253), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g335 ( .A(n_253), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_253), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g372 ( .A(n_253), .Y(n_372) );
INVx1_ASAP7_75t_L g405 ( .A(n_253), .Y(n_405) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g283 ( .A(n_254), .B(n_273), .Y(n_283) );
INVx1_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_260), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g496 ( .A(n_260), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_260), .A2(n_558), .B(n_559), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_270), .B1(n_276), .B2(n_283), .C(n_284), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_267), .B(n_287), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_267), .B(n_350), .Y(n_427) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_269), .B(n_317), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_269), .B(n_278), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_269), .B(n_292), .Y(n_421) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g343 ( .A(n_273), .Y(n_343) );
AND2x2_ASAP7_75t_L g318 ( .A(n_274), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g396 ( .A(n_274), .Y(n_396) );
AND2x2_ASAP7_75t_L g328 ( .A(n_275), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_275), .B(n_298), .Y(n_344) );
AND2x2_ASAP7_75t_L g408 ( .A(n_275), .B(n_334), .Y(n_408) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g317 ( .A(n_279), .B(n_286), .Y(n_317) );
AND2x2_ASAP7_75t_L g413 ( .A(n_280), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_282), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_283), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_283), .B(n_290), .Y(n_378) );
AND2x2_ASAP7_75t_L g398 ( .A(n_283), .B(n_298), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_283), .B(n_363), .Y(n_419) );
OAI32xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .A3(n_290), .B1(n_291), .B2(n_294), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_SL g292 ( .A(n_286), .Y(n_292) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_286), .B(n_316), .Y(n_333) );
OR2x2_ASAP7_75t_L g337 ( .A(n_286), .B(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_286), .B(n_385), .Y(n_438) );
INVx1_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
OAI221xp5_ASAP7_75t_SL g424 ( .A1(n_288), .A2(n_379), .B1(n_425), .B2(n_428), .C(n_429), .Y(n_424) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_289), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g339 ( .A(n_289), .B(n_312), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_289), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g417 ( .A(n_289), .B(n_350), .Y(n_417) );
INVxp67_ASAP7_75t_L g353 ( .A(n_290), .Y(n_353) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g423 ( .A(n_292), .B(n_410), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_292), .B(n_373), .Y(n_446) );
INVx1_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_294), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g439 ( .A(n_294), .B(n_440), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_299), .B(n_302), .Y(n_295) );
AND2x2_ASAP7_75t_L g308 ( .A(n_297), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g392 ( .A(n_301), .B(n_312), .Y(n_392) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g410 ( .A(n_303), .B(n_368), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_303), .B(n_367), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_304), .B(n_316), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_310), .C(n_320), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_306), .A2(n_341), .B1(n_345), .B2(n_348), .C(n_351), .Y(n_340) );
AOI31xp33_ASAP7_75t_L g435 ( .A1(n_306), .A2(n_436), .A3(n_437), .B(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B1(n_316), .B2(n_318), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g436 ( .A(n_316), .Y(n_436) );
INVx1_ASAP7_75t_L g399 ( .A(n_317), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_319), .A2(n_443), .B(n_445), .C(n_447), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_324), .B2(n_328), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_325), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_327), .A2(n_361), .B1(n_380), .B2(n_416), .C(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g411 ( .A(n_328), .Y(n_411) );
INVx1_ASAP7_75t_L g365 ( .A(n_329), .Y(n_365) );
NAND3xp33_ASAP7_75t_SL g330 ( .A(n_331), .B(n_340), .C(n_355), .Y(n_330) );
OAI21xp33_ASAP7_75t_L g381 ( .A1(n_332), .A2(n_382), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_334), .B(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g441 ( .A(n_335), .Y(n_441) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g379 ( .A(n_342), .B(n_362), .Y(n_379) );
INVx1_ASAP7_75t_L g354 ( .A(n_343), .Y(n_354) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g352 ( .A(n_346), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_346), .B(n_384), .Y(n_383) );
NOR4xp25_ASAP7_75t_L g351 ( .A(n_347), .B(n_352), .C(n_353), .D(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI222xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_360), .B1(n_366), .B2(n_367), .C1(n_369), .C2(n_373), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g453 ( .A(n_357), .Y(n_453) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_369), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g429 ( .A1(n_374), .A2(n_430), .B(n_432), .Y(n_429) );
NOR4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_387), .C(n_400), .D(n_415), .Y(n_375) );
OAI221xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_378), .B1(n_379), .B2(n_380), .C(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g456 ( .A(n_377), .Y(n_456) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_384), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OAI222xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_391), .B1(n_393), .B2(n_394), .C1(n_397), .C2(n_399), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_423), .B(n_424), .C(n_435), .Y(n_422) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
OAI222xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_406), .B1(n_407), .B2(n_409), .C1(n_411), .C2(n_412), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_417), .A2(n_420), .B1(n_453), .B2(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_450), .B(n_452), .C(n_455), .Y(n_447) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NOR2x2_ASAP7_75t_L g776 ( .A(n_463), .B(n_480), .Y(n_776) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_466), .A2(n_468), .B(n_777), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
INVx1_ASAP7_75t_L g478 ( .A(n_472), .Y(n_478) );
INVx1_ASAP7_75t_L g476 ( .A(n_473), .Y(n_476) );
INVx2_ASAP7_75t_L g773 ( .A(n_480), .Y(n_773) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_SL g482 ( .A(n_483), .B(n_739), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_643), .C(n_727), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_485), .B(n_586), .C(n_608), .D(n_624), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_524), .B1(n_547), .B2(n_565), .C(n_572), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_504), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_488), .B(n_565), .Y(n_598) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_488), .B(n_626), .C(n_639), .D(n_641), .Y(n_638) );
INVxp67_ASAP7_75t_L g755 ( .A(n_488), .Y(n_755) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g637 ( .A(n_489), .B(n_575), .Y(n_637) );
AND2x2_ASAP7_75t_L g661 ( .A(n_489), .B(n_504), .Y(n_661) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g628 ( .A(n_490), .B(n_564), .Y(n_628) );
AND2x2_ASAP7_75t_L g668 ( .A(n_490), .B(n_649), .Y(n_668) );
AND2x2_ASAP7_75t_L g685 ( .A(n_490), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_490), .B(n_505), .Y(n_709) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g563 ( .A(n_491), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g592 ( .A(n_491), .B(n_505), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_491), .B(n_514), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_500), .B(n_501), .C(n_502), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_502), .A2(n_511), .B(n_512), .Y(n_510) );
AND2x2_ASAP7_75t_L g595 ( .A(n_504), .B(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_504), .A2(n_645), .B1(n_648), .B2(n_650), .C(n_654), .Y(n_644) );
AND2x2_ASAP7_75t_L g703 ( .A(n_504), .B(n_668), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_504), .B(n_685), .Y(n_737) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
INVx3_ASAP7_75t_L g564 ( .A(n_505), .Y(n_564) );
AND2x2_ASAP7_75t_L g612 ( .A(n_505), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g666 ( .A(n_505), .B(n_581), .Y(n_666) );
AND2x2_ASAP7_75t_L g724 ( .A(n_505), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g565 ( .A(n_514), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g581 ( .A(n_514), .Y(n_581) );
INVx1_ASAP7_75t_L g636 ( .A(n_514), .Y(n_636) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_514), .Y(n_642) );
AND2x2_ASAP7_75t_L g687 ( .A(n_514), .B(n_564), .Y(n_687) );
OR2x2_ASAP7_75t_L g726 ( .A(n_514), .B(n_566), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_519), .B(n_522), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_524), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_532), .Y(n_524) );
AND2x2_ASAP7_75t_L g722 ( .A(n_525), .B(n_719), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_525), .B(n_704), .Y(n_754) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g653 ( .A(n_526), .B(n_577), .Y(n_653) );
AND2x2_ASAP7_75t_L g702 ( .A(n_526), .B(n_550), .Y(n_702) );
INVx1_ASAP7_75t_L g748 ( .A(n_526), .Y(n_748) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_527), .Y(n_562) );
AND2x2_ASAP7_75t_L g603 ( .A(n_527), .B(n_577), .Y(n_603) );
INVx1_ASAP7_75t_L g620 ( .A(n_527), .Y(n_620) );
AND2x2_ASAP7_75t_L g626 ( .A(n_527), .B(n_543), .Y(n_626) );
AND2x2_ASAP7_75t_L g694 ( .A(n_532), .B(n_602), .Y(n_694) );
INVx2_ASAP7_75t_L g759 ( .A(n_532), .Y(n_759) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_543), .Y(n_532) );
AND2x2_ASAP7_75t_L g576 ( .A(n_533), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g589 ( .A(n_533), .B(n_551), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_533), .B(n_550), .Y(n_617) );
INVx1_ASAP7_75t_L g623 ( .A(n_533), .Y(n_623) );
INVx1_ASAP7_75t_L g640 ( .A(n_533), .Y(n_640) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_533), .Y(n_652) );
INVx2_ASAP7_75t_L g720 ( .A(n_533), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B(n_538), .Y(n_535) );
INVx2_ASAP7_75t_L g577 ( .A(n_543), .Y(n_577) );
BUFx2_ASAP7_75t_L g674 ( .A(n_543), .Y(n_674) );
AND2x2_ASAP7_75t_L g719 ( .A(n_543), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_561), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_549), .B(n_656), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_549), .A2(n_718), .B(n_732), .Y(n_742) );
AND2x2_ASAP7_75t_L g767 ( .A(n_549), .B(n_653), .Y(n_767) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g689 ( .A(n_551), .Y(n_689) );
AND2x2_ASAP7_75t_L g718 ( .A(n_551), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_552), .Y(n_602) );
INVx2_ASAP7_75t_L g621 ( .A(n_552), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_552), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g575 ( .A(n_562), .Y(n_575) );
OR2x2_ASAP7_75t_L g588 ( .A(n_562), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g656 ( .A(n_562), .B(n_652), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_562), .B(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g757 ( .A(n_562), .B(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_562), .B(n_694), .Y(n_769) );
AND2x2_ASAP7_75t_L g648 ( .A(n_563), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g671 ( .A(n_563), .B(n_565), .Y(n_671) );
INVx2_ASAP7_75t_L g583 ( .A(n_564), .Y(n_583) );
AND2x2_ASAP7_75t_L g611 ( .A(n_564), .B(n_584), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_564), .B(n_636), .Y(n_692) );
AND2x2_ASAP7_75t_L g606 ( .A(n_565), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g753 ( .A(n_565), .Y(n_753) );
AND2x2_ASAP7_75t_L g765 ( .A(n_565), .B(n_628), .Y(n_765) );
AND2x2_ASAP7_75t_L g591 ( .A(n_566), .B(n_581), .Y(n_591) );
INVx1_ASAP7_75t_L g686 ( .A(n_566), .Y(n_686) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g584 ( .A(n_571), .B(n_585), .Y(n_584) );
INVxp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_575), .B(n_622), .Y(n_631) );
OR2x2_ASAP7_75t_L g763 ( .A(n_575), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g680 ( .A(n_576), .B(n_621), .Y(n_680) );
AND2x2_ASAP7_75t_L g688 ( .A(n_576), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g747 ( .A(n_576), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g771 ( .A(n_576), .B(n_618), .Y(n_771) );
NOR2xp67_ASAP7_75t_L g729 ( .A(n_577), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g758 ( .A(n_577), .B(n_621), .Y(n_758) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2x1p5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AND2x2_ASAP7_75t_L g610 ( .A(n_580), .B(n_611), .Y(n_610) );
INVxp67_ASAP7_75t_L g772 ( .A(n_580), .Y(n_772) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g607 ( .A(n_583), .Y(n_607) );
AND2x2_ASAP7_75t_L g658 ( .A(n_583), .B(n_591), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_583), .B(n_726), .Y(n_752) );
INVx2_ASAP7_75t_L g597 ( .A(n_584), .Y(n_597) );
INVx3_ASAP7_75t_L g649 ( .A(n_584), .Y(n_649) );
OR2x2_ASAP7_75t_L g677 ( .A(n_584), .B(n_678), .Y(n_677) );
AOI311xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_590), .A3(n_592), .B(n_593), .C(n_604), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_587), .A2(n_625), .B(n_627), .C(n_629), .Y(n_624) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_SL g609 ( .A(n_589), .Y(n_609) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g627 ( .A(n_591), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_591), .B(n_607), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_591), .B(n_592), .Y(n_760) );
AND2x2_ASAP7_75t_L g682 ( .A(n_592), .B(n_596), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B(n_599), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g740 ( .A(n_596), .B(n_628), .Y(n_740) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_597), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g634 ( .A(n_597), .Y(n_634) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g625 ( .A(n_601), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g670 ( .A(n_603), .Y(n_670) );
AND2x4_ASAP7_75t_L g732 ( .A(n_603), .B(n_701), .Y(n_732) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_606), .A2(n_672), .B1(n_684), .B2(n_688), .C1(n_690), .C2(n_694), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_612), .C(n_615), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_609), .B(n_653), .Y(n_676) );
INVx1_ASAP7_75t_L g698 ( .A(n_611), .Y(n_698) );
INVx1_ASAP7_75t_L g632 ( .A(n_613), .Y(n_632) );
OR2x2_ASAP7_75t_L g697 ( .A(n_614), .B(n_698), .Y(n_697) );
OAI21xp33_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_618), .B(n_622), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_616), .B(n_634), .C(n_635), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_616), .A2(n_653), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_620), .Y(n_673) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_621), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g730 ( .A(n_621), .Y(n_730) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_621), .Y(n_746) );
INVx2_ASAP7_75t_L g704 ( .A(n_622), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_626), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g678 ( .A(n_628), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B1(n_633), .B2(n_637), .C(n_638), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_632), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g766 ( .A(n_632), .Y(n_766) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g647 ( .A(n_639), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_639), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g705 ( .A(n_639), .B(n_653), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_639), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g738 ( .A(n_639), .B(n_673), .Y(n_738) );
BUFx3_ASAP7_75t_L g701 ( .A(n_640), .Y(n_701) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND5xp2_ASAP7_75t_L g643 ( .A(n_644), .B(n_662), .C(n_683), .D(n_695), .E(n_710), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI32xp33_ASAP7_75t_L g735 ( .A1(n_647), .A2(n_674), .A3(n_690), .B1(n_736), .B2(n_738), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_649), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g659 ( .A(n_653), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_669), .B1(n_671), .B2(n_672), .C(n_675), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g734 ( .A(n_666), .B(n_685), .Y(n_734) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_671), .A2(n_732), .B1(n_750), .B2(n_755), .C(n_756), .Y(n_749) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx2_ASAP7_75t_L g715 ( .A(n_674), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_679), .B2(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g693 ( .A(n_685), .Y(n_693) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_699), .B1(n_703), .B2(n_704), .C1(n_705), .C2(n_706), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_704), .A2(n_751), .B1(n_753), .B2(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .B(n_716), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_721), .B(n_723), .Y(n_716) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g764 ( .A(n_719), .Y(n_764) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_731), .B(n_733), .C(n_735), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AOI211xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_743), .C(n_768), .Y(n_739) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_740), .Y(n_744) );
INVxp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_749), .C(n_761), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B(n_760), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AOI21xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B(n_772), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
endmodule