module real_jpeg_377_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_0),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_1),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_147),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_147),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_66),
.B1(n_67),
.B2(n_147),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_2),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_125),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_125),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_125),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_47),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_47),
.B1(n_66),
.B2(n_67),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_6),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_7),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_87),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_87),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_87),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_55),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_8),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_56),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_9),
.B(n_29),
.C(n_31),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_9),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_28),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_9),
.B(n_63),
.C(n_66),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_214),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_9),
.B(n_115),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_9),
.B(n_69),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_214),
.Y(n_279)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B(n_345),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_13),
.B(n_346),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_14),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_79),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_79),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_14),
.A2(n_66),
.B1(n_67),
.B2(n_79),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_16),
.A2(n_44),
.B1(n_45),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_179),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_16),
.A2(n_66),
.B1(n_67),
.B2(n_179),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_17),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_40),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_17),
.A2(n_40),
.B1(n_66),
.B2(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_17),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_340),
.B(n_343),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_332),
.B(n_336),
.Y(n_21)
);

AOI21x1_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_92),
.B(n_331),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_80),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_24),
.B(n_80),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_59),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_27),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_28),
.B(n_176),
.Y(n_280)
);

AO22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_30),
.A2(n_31),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_31),
.B(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_35),
.B(n_204),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g228 ( 
.A(n_35),
.B(n_51),
.Y(n_228)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g226 ( 
.A1(n_36),
.A2(n_45),
.A3(n_50),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_41),
.B(n_57),
.C(n_59),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_54),
.B2(n_56),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_49),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_45),
.A2(n_77),
.B(n_214),
.C(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_45),
.B(n_214),
.Y(n_215)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_48),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_48),
.A2(n_56),
.B1(n_146),
.B2(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_48),
.A2(n_54),
.B1(n_56),
.B2(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_48),
.A2(n_56),
.B(n_334),
.Y(n_342)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_77),
.B1(n_78),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_49),
.A2(n_86),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_49),
.B(n_124),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_49),
.A2(n_122),
.B(n_300),
.Y(n_299)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_72),
.C(n_76),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_72),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_85),
.C(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_61),
.A2(n_69),
.B1(n_120),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_61),
.A2(n_69),
.B1(n_141),
.B2(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_61),
.A2(n_196),
.B(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_61),
.B(n_200),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_71),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_101),
.B1(n_102),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_65),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_65),
.A2(n_221),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_65),
.A2(n_101),
.B1(n_197),
.B2(n_247),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_66),
.B(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_69),
.B(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_75),
.B1(n_91),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_73),
.A2(n_75),
.B1(n_99),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_73),
.A2(n_75),
.B1(n_187),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_73),
.A2(n_279),
.B(n_280),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_73),
.A2(n_218),
.B(n_280),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_75),
.A2(n_143),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_75),
.A2(n_175),
.B(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_77),
.A2(n_145),
.B(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_88),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_81),
.A2(n_85),
.B1(n_105),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_155),
.B(n_328),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_150),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_126),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_95),
.B(n_126),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_103),
.C(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_101),
.A2(n_199),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_121),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_109),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_111),
.B1(n_121),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_111),
.B1(n_118),
.B2(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_115),
.B(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_112),
.A2(n_115),
.B1(n_138),
.B2(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_112),
.A2(n_214),
.B(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_113),
.A2(n_114),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_113),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_113),
.A2(n_114),
.B1(n_194),
.B2(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_113),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_113),
.A2(n_114),
.B1(n_239),
.B2(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_114),
.A2(n_193),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_114),
.B(n_208),
.Y(n_241)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_115),
.A2(n_207),
.B(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_133),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_142),
.C(n_144),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_135),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_136),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_144),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_149),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_150),
.A2(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_151),
.B(n_154),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_180),
.B(n_327),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_157),
.B(n_160),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_161),
.B(n_164),
.Y(n_325)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_166),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.C(n_177),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_167),
.A2(n_168),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_169),
.B(n_171),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_177),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_178),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_322),
.B(n_326),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_291),
.B(n_319),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_233),
.B(n_290),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_209),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_184),
.B(n_209),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.C(n_201),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_185),
.B(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_189),
.C(n_192),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_201),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_223),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_210),
.B(n_224),
.C(n_232),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_222),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_211),
.B(n_217),
.C(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_232),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_225),
.B(n_230),
.Y(n_295)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_285),
.B(n_289),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_274),
.B(n_284),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_256),
.B(n_273),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_250),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_250),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_242),
.B1(n_248),
.B2(n_249),
.Y(n_237)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_245),
.C(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_267),
.B(n_272),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_262),
.B(n_266),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_265),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_264),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_270),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_276),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_306),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_305),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_305),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_302),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_303),
.C(n_304),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_297),
.C(n_301),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_301),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_318),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_318),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_312),
.C(n_314),
.Y(n_323)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_324),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_333),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_333),
.B(n_341),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_335),
.Y(n_339)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_338),
.B(n_342),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);


endmodule