module fake_jpeg_31806_n_497 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_497);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_497;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_461;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_13),
.B(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_8),
.C(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_52),
.B(n_64),
.Y(n_154)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_8),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_54),
.B(n_67),
.Y(n_143)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_18),
.B(n_8),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_75),
.B(n_83),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx12f_ASAP7_75t_SL g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_7),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_7),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_95),
.B(n_24),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_34),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_9),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

CKINVDCx9p33_ASAP7_75t_R g98 ( 
.A(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_22),
.B1(n_25),
.B2(n_46),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_102),
.A2(n_114),
.B1(n_130),
.B2(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_105),
.B(n_10),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_109),
.B1(n_116),
.B2(n_121),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_44),
.B1(n_49),
.B2(n_37),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_78),
.B1(n_72),
.B2(n_68),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_35),
.B1(n_47),
.B2(n_45),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_63),
.A2(n_87),
.B1(n_82),
.B2(n_84),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_51),
.A2(n_37),
.B1(n_44),
.B2(n_49),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_129),
.A2(n_20),
.B1(n_17),
.B2(n_50),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_61),
.A2(n_38),
.B1(n_32),
.B2(n_29),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_69),
.A2(n_38),
.B1(n_32),
.B2(n_29),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_60),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_142),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_65),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_76),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_152),
.B1(n_86),
.B2(n_81),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_90),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_155),
.B(n_188),
.Y(n_209)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_104),
.A2(n_94),
.B1(n_53),
.B2(n_96),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_183),
.B1(n_193),
.B2(n_203),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_74),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_189),
.Y(n_221)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_58),
.C(n_70),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_176),
.Y(n_217)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_79),
.B1(n_62),
.B2(n_89),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_126),
.B(n_80),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_179),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_17),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_131),
.B1(n_117),
.B2(n_113),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_182),
.A2(n_187),
.B1(n_190),
.B2(n_192),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_109),
.A2(n_77),
.B1(n_89),
.B2(n_97),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_185),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_50),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_122),
.A2(n_17),
.B1(n_20),
.B2(n_2),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_191),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_122),
.A2(n_133),
.B1(n_127),
.B2(n_103),
.Y(n_192)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_202),
.B1(n_205),
.B2(n_135),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_140),
.A2(n_50),
.B1(n_39),
.B2(n_2),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_195),
.A2(n_108),
.B1(n_110),
.B2(n_124),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_199),
.Y(n_231)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_198),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_108),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_50),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_39),
.B1(n_9),
.B2(n_3),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_206),
.Y(n_227)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_107),
.B(n_39),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_133),
.B1(n_127),
.B2(n_103),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_208),
.A2(n_234),
.B1(n_184),
.B2(n_1),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_155),
.A2(n_107),
.B1(n_134),
.B2(n_136),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_153),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_236),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_177),
.A2(n_115),
.B1(n_141),
.B2(n_123),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_153),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_164),
.A2(n_141),
.B1(n_140),
.B2(n_115),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_243),
.B1(n_187),
.B2(n_213),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_161),
.B1(n_183),
.B2(n_179),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_124),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_246),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_177),
.A2(n_110),
.B1(n_112),
.B2(n_5),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_171),
.B(n_180),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_161),
.A2(n_12),
.B(n_5),
.C(n_6),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_176),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_180),
.B(n_0),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_249),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_163),
.B(n_0),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g251 ( 
.A1(n_161),
.A2(n_112),
.A3(n_39),
.B1(n_6),
.B2(n_11),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_183),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_252),
.A2(n_266),
.B(n_235),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_160),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_253),
.B(n_255),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_250),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_254),
.B(n_257),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_200),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_256),
.A2(n_265),
.B1(n_268),
.B2(n_271),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_189),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_211),
.B(n_175),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_261),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_207),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_241),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_262),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_209),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_263),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_211),
.B(n_159),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_282),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_243),
.A2(n_183),
.B1(n_204),
.B2(n_167),
.Y(n_265)
);

BUFx8_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_176),
.B1(n_170),
.B2(n_158),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_236),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_279),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_205),
.B1(n_202),
.B2(n_198),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_212),
.A2(n_232),
.B1(n_213),
.B2(n_234),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_272),
.A2(n_274),
.B1(n_283),
.B2(n_245),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_273),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_239),
.A2(n_191),
.B1(n_194),
.B2(n_156),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_277),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_220),
.B(n_222),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_278),
.B(n_288),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_216),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_157),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_221),
.B(n_173),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_221),
.A2(n_165),
.B1(n_181),
.B2(n_172),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_196),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_284),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_285),
.A2(n_286),
.B1(n_215),
.B2(n_235),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_208),
.A2(n_12),
.B1(n_15),
.B2(n_6),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_228),
.B(n_0),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_227),
.B(n_184),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_290),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_184),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_291),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_266),
.A2(n_212),
.B(n_247),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_292),
.A2(n_294),
.B(n_310),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_293),
.A2(n_295),
.B1(n_314),
.B2(n_268),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_238),
.B(n_248),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_252),
.A2(n_238),
.B1(n_222),
.B2(n_251),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_298),
.B(n_309),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_270),
.B(n_229),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_328),
.Y(n_329)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_312),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_233),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_258),
.C(n_290),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_280),
.A2(n_242),
.B1(n_245),
.B2(n_229),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_315),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_317),
.A2(n_257),
.B1(n_285),
.B2(n_282),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_318),
.B(n_261),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_262),
.A2(n_233),
.B(n_225),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_291),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_330),
.B(n_331),
.C(n_352),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_291),
.C(n_275),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_263),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_339),
.Y(n_378)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_310),
.A2(n_260),
.A3(n_287),
.B1(n_279),
.B2(n_255),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_353),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_289),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_338),
.B(n_292),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_319),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_340),
.A2(n_360),
.B1(n_311),
.B2(n_301),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_320),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_346),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_309),
.A2(n_272),
.B1(n_256),
.B2(n_278),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_343),
.A2(n_347),
.B1(n_355),
.B2(n_307),
.Y(n_365)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_296),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_348),
.Y(n_383)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_303),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_357),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_275),
.C(n_289),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_299),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_253),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_354),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_311),
.A2(n_317),
.B1(n_326),
.B2(n_319),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_328),
.C(n_294),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_226),
.C(n_237),
.Y(n_387)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_296),
.B(n_284),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_316),
.C(n_300),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_288),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_267),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_307),
.A2(n_293),
.B1(n_301),
.B2(n_295),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_307),
.B(n_319),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_361),
.A2(n_369),
.B(n_332),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_375),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_363),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_365),
.A2(n_367),
.B1(n_372),
.B2(n_374),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_342),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_347),
.A2(n_314),
.B1(n_316),
.B2(n_324),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_310),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_344),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_344),
.A2(n_322),
.B(n_323),
.Y(n_369)
);

AOI22x1_ASAP7_75t_L g370 ( 
.A1(n_351),
.A2(n_325),
.B1(n_265),
.B2(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_341),
.A2(n_325),
.B1(n_274),
.B2(n_305),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_355),
.A2(n_300),
.B1(n_305),
.B2(n_315),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_340),
.A2(n_321),
.B1(n_304),
.B2(n_308),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_336),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_376),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_335),
.A2(n_321),
.B(n_306),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_377),
.B(n_388),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_306),
.B1(n_327),
.B2(n_254),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_379),
.A2(n_382),
.B1(n_372),
.B2(n_367),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_327),
.Y(n_381)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_381),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_254),
.B1(n_273),
.B2(n_286),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_329),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_386),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_356),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_329),
.Y(n_388)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_389),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_381),
.B(n_379),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_371),
.A2(n_360),
.B1(n_349),
.B2(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_391),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_368),
.C(n_387),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_393),
.C(n_395),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_330),
.C(n_338),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_399),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_352),
.C(n_332),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_377),
.C(n_374),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_401),
.C(n_403),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_344),
.C(n_357),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_388),
.C(n_386),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_407),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_342),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_408),
.A2(n_364),
.B1(n_383),
.B2(n_382),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_337),
.C(n_333),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_371),
.C(n_376),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_361),
.A2(n_337),
.B(n_333),
.Y(n_411)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_411),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_410),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_416),
.Y(n_446)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_399),
.B(n_375),
.CI(n_362),
.CON(n_416),
.SN(n_416)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_396),
.A2(n_380),
.B1(n_378),
.B2(n_370),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_421),
.A2(n_230),
.B1(n_237),
.B2(n_226),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_403),
.A2(n_385),
.B(n_370),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_427),
.B(n_390),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_385),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_424),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_389),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_425),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_433),
.C(n_406),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_364),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_429),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_383),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_397),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_405),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_267),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_432),
.A2(n_396),
.B1(n_402),
.B2(n_404),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_395),
.B(n_401),
.C(n_400),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_440),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_449),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_407),
.C(n_408),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_438),
.C(n_443),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_397),
.C(n_413),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_448),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_409),
.C(n_402),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_409),
.C(n_412),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_428),
.C(n_430),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_445),
.A2(n_432),
.B1(n_417),
.B2(n_419),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_422),
.A2(n_230),
.B(n_210),
.Y(n_447)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_447),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_418),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_452),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_446),
.A2(n_418),
.B(n_433),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_439),
.A2(n_445),
.B1(n_441),
.B2(n_421),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_458),
.Y(n_468)
);

XNOR2x1_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_223),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_442),
.A2(n_427),
.B1(n_426),
.B2(n_416),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_426),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_460),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_416),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_420),
.C(n_225),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_440),
.C(n_210),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_437),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_214),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_460),
.A2(n_443),
.B(n_436),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_469),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_470),
.Y(n_483)
);

AOI21xp33_ASAP7_75t_L g467 ( 
.A1(n_455),
.A2(n_267),
.B(n_223),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_467),
.A2(n_11),
.B(n_14),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_267),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_451),
.B(n_214),
.Y(n_472)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_472),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_475),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_0),
.C(n_1),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_474),
.B(n_1),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_6),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_479),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_471),
.A2(n_461),
.B(n_454),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_462),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_462),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_464),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_484),
.B(n_485),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_481),
.Y(n_485)
);

NOR2x1_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_472),
.Y(n_486)
);

NAND4xp25_ASAP7_75t_SL g489 ( 
.A(n_486),
.B(n_476),
.C(n_468),
.D(n_465),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_457),
.C(n_470),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_489),
.A2(n_490),
.B(n_486),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_492),
.A2(n_493),
.B(n_483),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_491),
.A2(n_466),
.B(n_478),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_494),
.A2(n_483),
.B(n_457),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_487),
.B(n_15),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_496),
.A2(n_15),
.B(n_1),
.Y(n_497)
);


endmodule