module fake_aes_4105_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
HB1xp67_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_10), .B(n_4), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_0), .B(n_3), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_1), .B(n_9), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_13), .B(n_15), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_11), .B(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_14), .B(n_2), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_17), .B1(n_18), .B2(n_3), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_17), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_21), .B(n_19), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_18), .B1(n_26), .B2(n_23), .Y(n_28) );
NAND4xp25_ASAP7_75t_L g29 ( .A(n_25), .B(n_1), .C(n_2), .D(n_4), .Y(n_29) );
OAI221xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_19), .B1(n_20), .B2(n_7), .C(n_8), .Y(n_30) );
OAI211xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_20), .B(n_19), .C(n_7), .Y(n_31) );
OAI222xp33_ASAP7_75t_L g32 ( .A1(n_27), .A2(n_5), .B1(n_6), .B2(n_8), .C1(n_9), .C2(n_20), .Y(n_32) );
INVx2_ASAP7_75t_SL g33 ( .A(n_30), .Y(n_33) );
CKINVDCx16_ASAP7_75t_R g34 ( .A(n_32), .Y(n_34) );
AOI221xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_30), .B1(n_31), .B2(n_19), .C(n_5), .Y(n_35) );
AO221x1_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_19), .B1(n_33), .B2(n_32), .C(n_34), .Y(n_36) );
endmodule