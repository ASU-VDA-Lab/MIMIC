module fake_ibex_1202_n_837 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_837);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_837;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_682;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_798;
wire n_832;
wire n_732;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_787;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_772;
wire n_810;
wire n_768;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_640;
wire n_477;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_801;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_71),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_60),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_10),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_86),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_21),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_18),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_39),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_147),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_127),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_36),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_32),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx4_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_62),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_49),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_4),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_73),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_120),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_67),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_23),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_80),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_87),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_46),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_157),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_15),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_74),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_119),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_17),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_124),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_109),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_72),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_133),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_55),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_130),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_152),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_117),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_160),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_9),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_114),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_51),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_10),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_138),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_128),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_92),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_18),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_171),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_L g258 ( 
.A(n_70),
.B(n_163),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_26),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_143),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_15),
.B(n_8),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_123),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_153),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_85),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_76),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_27),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_26),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_155),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_174),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_167),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_33),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_90),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_58),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_112),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_129),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_6),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_135),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_47),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_27),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_35),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_33),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_156),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_3),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_108),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_144),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_162),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_173),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_131),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_259),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_180),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_185),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_2),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_182),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_182),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_196),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

BUFx8_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_211),
.B(n_3),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_196),
.B(n_4),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_259),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_187),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_176),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_223),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_288),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_243),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_223),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_177),
.B(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_187),
.B(n_12),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_192),
.B(n_193),
.Y(n_316)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_190),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_186),
.A2(n_81),
.B(n_170),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_265),
.B(n_13),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_180),
.B(n_13),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_206),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_186),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_234),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_238),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_275),
.B(n_16),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_195),
.A2(n_78),
.B(n_168),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_195),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_181),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_178),
.B(n_16),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_200),
.B(n_17),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_217),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_217),
.B(n_19),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_275),
.B(n_19),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_202),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_218),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_219),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_247),
.B(n_20),
.Y(n_342)
);

BUFx8_ASAP7_75t_L g343 ( 
.A(n_219),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_250),
.B(n_252),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_224),
.B(n_20),
.Y(n_345)
);

CKINVDCx11_ASAP7_75t_R g346 ( 
.A(n_234),
.Y(n_346)
);

OAI21x1_ASAP7_75t_L g347 ( 
.A1(n_224),
.A2(n_84),
.B(n_165),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_267),
.B(n_292),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_236),
.B(n_21),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g351 ( 
.A(n_292),
.B(n_42),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_179),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_183),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_184),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_191),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_188),
.B(n_22),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_194),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_197),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_260),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_356),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_322),
.B(n_199),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_189),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_304),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_317),
.B(n_208),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_326),
.Y(n_367)
);

OR2x6_ASAP7_75t_L g368 ( 
.A(n_294),
.B(n_261),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_347),
.A2(n_216),
.B(n_213),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_306),
.B(n_236),
.Y(n_372)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_317),
.B(n_221),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

OR2x6_ASAP7_75t_L g379 ( 
.A(n_305),
.B(n_269),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_322),
.B(n_222),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_304),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_304),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_356),
.A2(n_293),
.B1(n_282),
.B2(n_257),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_348),
.B(n_225),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_317),
.B(n_228),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_317),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_297),
.B(n_324),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_300),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_310),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_301),
.B(n_230),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_310),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_348),
.B(n_231),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_303),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_316),
.A2(n_293),
.B1(n_282),
.B2(n_257),
.Y(n_401)
);

AOI21x1_ASAP7_75t_L g402 ( 
.A1(n_347),
.A2(n_233),
.B(n_232),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_310),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_349),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_324),
.B(n_237),
.Y(n_405)
);

NAND3xp33_ASAP7_75t_L g406 ( 
.A(n_296),
.B(n_227),
.C(n_212),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_298),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_326),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_302),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_311),
.B(n_268),
.C(n_229),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_299),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_325),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_295),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_324),
.Y(n_416)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_332),
.B(n_239),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_352),
.B(n_240),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_332),
.B(n_242),
.Y(n_421)
);

OAI22x1_ASAP7_75t_L g422 ( 
.A1(n_357),
.A2(n_281),
.B1(n_280),
.B2(n_286),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g423 ( 
.A1(n_319),
.A2(n_245),
.B(n_244),
.Y(n_423)
);

AO21x2_ASAP7_75t_L g424 ( 
.A1(n_357),
.A2(n_249),
.B(n_246),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_308),
.Y(n_425)
);

AO21x2_ASAP7_75t_L g426 ( 
.A1(n_342),
.A2(n_253),
.B(n_251),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_308),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_302),
.B(n_255),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_L g429 ( 
.A(n_351),
.B(n_198),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_309),
.B(n_263),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_411),
.B(n_343),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_343),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_343),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_415),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_360),
.B(n_355),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_363),
.B(n_318),
.Y(n_438)
);

OAI22xp33_ASAP7_75t_L g439 ( 
.A1(n_379),
.A2(n_315),
.B1(n_320),
.B2(n_329),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_404),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_337),
.Y(n_441)
);

NOR3xp33_ASAP7_75t_L g442 ( 
.A(n_412),
.B(n_333),
.C(n_314),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_398),
.B(n_323),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_339),
.Y(n_444)
);

BUFx6f_ASAP7_75t_SL g445 ( 
.A(n_379),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_388),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_372),
.B(n_359),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_387),
.B(n_344),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_365),
.A2(n_358),
.B1(n_353),
.B2(n_341),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

OAI22x1_ASAP7_75t_L g451 ( 
.A1(n_401),
.A2(n_346),
.B1(n_285),
.B2(n_272),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_340),
.Y(n_452)
);

BUFx12f_ASAP7_75t_SL g453 ( 
.A(n_379),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_382),
.B(n_264),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_393),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_384),
.B(n_264),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_346),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_361),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_381),
.B(n_354),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_279),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_366),
.B(n_279),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_364),
.A2(n_289),
.B1(n_290),
.B2(n_214),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_374),
.B(n_289),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_391),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_375),
.A2(n_350),
.B1(n_341),
.B2(n_335),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_417),
.B(n_351),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_390),
.B(n_201),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_362),
.B(n_266),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_413),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_389),
.B(n_203),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_362),
.B(n_270),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_364),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_369),
.B(n_204),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_370),
.A2(n_271),
.B1(n_273),
.B2(n_277),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_368),
.B(n_22),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_380),
.B(n_278),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_379),
.B(n_330),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_389),
.B(n_205),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_399),
.B(n_210),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_406),
.B(n_226),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_376),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_396),
.B(n_330),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_391),
.B(n_215),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_378),
.B(n_258),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_431),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_416),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_380),
.A2(n_207),
.B1(n_287),
.B2(n_291),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_399),
.B(n_220),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_368),
.B(n_330),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_417),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_426),
.A2(n_283),
.B1(n_276),
.B2(n_254),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_368),
.A2(n_209),
.B1(n_24),
.B2(n_25),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_426),
.B(n_23),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_373),
.B(n_44),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_422),
.B(n_24),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_420),
.B(n_28),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_424),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_405),
.B(n_45),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_429),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_368),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_468),
.B(n_487),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_459),
.B(n_367),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_459),
.B(n_367),
.Y(n_512)
);

AO21x1_ASAP7_75t_L g513 ( 
.A1(n_498),
.A2(n_371),
.B(n_402),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_460),
.B(n_423),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_458),
.B(n_409),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_457),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_480),
.A2(n_437),
.B(n_494),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_444),
.B(n_427),
.Y(n_519)
);

A2O1A1Ixp33_ASAP7_75t_L g520 ( 
.A1(n_438),
.A2(n_377),
.B(n_383),
.C(n_385),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_452),
.A2(n_427),
.B(n_386),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_444),
.B(n_31),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_458),
.B(n_448),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_475),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_32),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_34),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_451),
.B(n_409),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_497),
.B(n_478),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_470),
.B(n_37),
.Y(n_532)
);

AO21x1_ASAP7_75t_L g533 ( 
.A1(n_502),
.A2(n_410),
.B(n_394),
.Y(n_533)
);

BUFx8_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

CKINVDCx10_ASAP7_75t_R g535 ( 
.A(n_445),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_482),
.A2(n_425),
.B1(n_408),
.B2(n_397),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_474),
.B(n_37),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_479),
.B(n_38),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_464),
.B(n_40),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_L g540 ( 
.A1(n_462),
.A2(n_479),
.B(n_443),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_453),
.B(n_40),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_433),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_454),
.A2(n_403),
.B(n_48),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_443),
.B(n_41),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_456),
.B(n_50),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_432),
.Y(n_546)
);

OAI321xp33_ASAP7_75t_L g547 ( 
.A1(n_506),
.A2(n_403),
.A3(n_53),
.B1(n_54),
.B2(n_56),
.C(n_57),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_435),
.Y(n_548)
);

CKINVDCx10_ASAP7_75t_R g549 ( 
.A(n_500),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_496),
.A2(n_52),
.B1(n_59),
.B2(n_61),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_476),
.B(n_63),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_461),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_491),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_489),
.B(n_66),
.Y(n_554)
);

AO21x1_ASAP7_75t_L g555 ( 
.A1(n_499),
.A2(n_68),
.B(n_69),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_446),
.A2(n_436),
.B(n_450),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_449),
.B(n_75),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_466),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_504),
.A2(n_77),
.B(n_82),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_473),
.A2(n_493),
.B(n_483),
.Y(n_560)
);

BUFx4f_ASAP7_75t_L g561 ( 
.A(n_485),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_481),
.A2(n_88),
.B(n_89),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_484),
.A2(n_95),
.B(n_96),
.C(n_98),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_455),
.A2(n_99),
.B(n_101),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_501),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_467),
.B(n_102),
.Y(n_566)
);

OAI321xp33_ASAP7_75t_L g567 ( 
.A1(n_506),
.A2(n_103),
.A3(n_105),
.B1(n_106),
.B2(n_110),
.C(n_111),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_463),
.A2(n_113),
.B1(n_121),
.B2(n_126),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_492),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_465),
.B(n_164),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_469),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_486),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_488),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_523),
.B(n_505),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_511),
.Y(n_575)
);

BUFx12f_ASAP7_75t_L g576 ( 
.A(n_534),
.Y(n_576)
);

NAND2x1p5_ASAP7_75t_L g577 ( 
.A(n_507),
.B(n_527),
.Y(n_577)
);

AO31x2_ASAP7_75t_L g578 ( 
.A1(n_509),
.A2(n_141),
.A3(n_142),
.B(n_146),
.Y(n_578)
);

AO31x2_ASAP7_75t_L g579 ( 
.A1(n_520),
.A2(n_555),
.A3(n_518),
.B(n_550),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_569),
.B(n_526),
.Y(n_580)
);

AO31x2_ASAP7_75t_L g581 ( 
.A1(n_563),
.A2(n_529),
.A3(n_544),
.B(n_562),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_512),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_508),
.B(n_517),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

OR2x6_ASAP7_75t_L g585 ( 
.A(n_541),
.B(n_524),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_552),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_561),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_531),
.B(n_516),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_528),
.A2(n_522),
.B1(n_519),
.B2(n_571),
.Y(n_589)
);

AO31x2_ASAP7_75t_L g590 ( 
.A1(n_559),
.A2(n_565),
.A3(n_557),
.B(n_566),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_535),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_539),
.B(n_573),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_546),
.B(n_548),
.Y(n_593)
);

AO31x2_ASAP7_75t_L g594 ( 
.A1(n_532),
.A2(n_537),
.A3(n_538),
.B(n_564),
.Y(n_594)
);

AO31x2_ASAP7_75t_L g595 ( 
.A1(n_570),
.A2(n_525),
.A3(n_556),
.B(n_543),
.Y(n_595)
);

INVx6_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_542),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_515),
.Y(n_598)
);

AO31x2_ASAP7_75t_L g599 ( 
.A1(n_521),
.A2(n_545),
.A3(n_536),
.B(n_554),
.Y(n_599)
);

OAI21xp33_ASAP7_75t_SL g600 ( 
.A1(n_551),
.A2(n_568),
.B(n_553),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_572),
.A2(n_547),
.B(n_567),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_530),
.B(n_558),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_510),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_510),
.B(n_490),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_527),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_L g607 ( 
.A1(n_540),
.A2(n_444),
.B(n_460),
.Y(n_607)
);

A2O1A1Ixp33_ASAP7_75t_L g608 ( 
.A1(n_540),
.A2(n_444),
.B(n_560),
.C(n_438),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_527),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_511),
.B(n_459),
.Y(n_610)
);

NAND2x1p5_ASAP7_75t_L g611 ( 
.A(n_507),
.B(n_527),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_510),
.B(n_490),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_510),
.B(n_490),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_523),
.A2(n_531),
.B1(n_528),
.B2(n_526),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_510),
.B(n_490),
.Y(n_615)
);

AO31x2_ASAP7_75t_L g616 ( 
.A1(n_533),
.A2(n_513),
.A3(n_509),
.B(n_514),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_540),
.A2(n_444),
.B(n_560),
.C(n_438),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_510),
.B(n_448),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_527),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_527),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_510),
.B(n_448),
.Y(n_621)
);

AOI21xp33_ASAP7_75t_L g622 ( 
.A1(n_523),
.A2(n_434),
.B(n_419),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_523),
.B(n_472),
.Y(n_623)
);

AOI21x1_ASAP7_75t_L g624 ( 
.A1(n_513),
.A2(n_509),
.B(n_518),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_SL g625 ( 
.A(n_529),
.B(n_326),
.C(n_367),
.Y(n_625)
);

AOI21xp33_ASAP7_75t_L g626 ( 
.A1(n_523),
.A2(n_434),
.B(n_419),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_515),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_541),
.B(n_387),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_510),
.B(n_490),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_510),
.B(n_490),
.Y(n_630)
);

AND3x4_ASAP7_75t_L g631 ( 
.A(n_531),
.B(n_412),
.C(n_441),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_510),
.B(n_490),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_510),
.B(n_490),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_SL g634 ( 
.A1(n_523),
.A2(n_439),
.B(n_434),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_511),
.B(n_459),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_510),
.B(n_490),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_510),
.B(n_490),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_490),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_510),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_510),
.B(n_490),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_510),
.B(n_490),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_510),
.B(n_490),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_510),
.B(n_448),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_514),
.A2(n_560),
.B(n_509),
.Y(n_644)
);

BUFx2_ASAP7_75t_R g645 ( 
.A(n_517),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_510),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_527),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_510),
.B(n_490),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_608),
.A2(n_617),
.B(n_607),
.C(n_634),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_607),
.A2(n_628),
.B1(n_618),
.B2(n_643),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_632),
.B1(n_648),
.B2(n_629),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_639),
.B(n_646),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_612),
.B(n_613),
.Y(n_653)
);

AO21x2_ASAP7_75t_L g654 ( 
.A1(n_601),
.A2(n_644),
.B(n_624),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_610),
.B(n_635),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_620),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_645),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_576),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_606),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_L g660 ( 
.A1(n_634),
.A2(n_592),
.B1(n_638),
.B2(n_615),
.C(n_642),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_577),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_584),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_611),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_586),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_598),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_646),
.B(n_582),
.Y(n_666)
);

A2O1A1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_630),
.A2(n_633),
.B(n_636),
.C(n_637),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_640),
.A2(n_641),
.B(n_574),
.C(n_600),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_591),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_596),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_596),
.Y(n_671)
);

AOI221xp5_ASAP7_75t_L g672 ( 
.A1(n_622),
.A2(n_626),
.B1(n_575),
.B2(n_625),
.C(n_623),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_621),
.B(n_614),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_628),
.A2(n_631),
.B1(n_614),
.B2(n_583),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_580),
.B(n_588),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_603),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_588),
.B(n_589),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_603),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_597),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_581),
.B(n_600),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_593),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_581),
.B(n_616),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_627),
.A2(n_581),
.B(n_616),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_609),
.Y(n_684)
);

AO31x2_ASAP7_75t_L g685 ( 
.A1(n_616),
.A2(n_579),
.A3(n_578),
.B(n_594),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_603),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_595),
.A2(n_579),
.B(n_590),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_587),
.B(n_585),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_SL g689 ( 
.A1(n_578),
.A2(n_579),
.B(n_590),
.C(n_594),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_619),
.B(n_647),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_595),
.A2(n_590),
.B(n_599),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_585),
.A2(n_602),
.B1(n_599),
.B2(n_594),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_599),
.A2(n_617),
.B(n_608),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_576),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_576),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_605),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_592),
.B(n_622),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_576),
.B(n_387),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_607),
.A2(n_628),
.B1(n_618),
.B2(n_621),
.Y(n_699)
);

AO32x2_ASAP7_75t_L g700 ( 
.A1(n_589),
.A2(n_550),
.A3(n_497),
.B1(n_477),
.B2(n_616),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

OAI222xp33_ASAP7_75t_L g702 ( 
.A1(n_628),
.A2(n_588),
.B1(n_614),
.B2(n_585),
.C1(n_387),
.C2(n_448),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_SL g703 ( 
.A1(n_628),
.A2(n_326),
.B1(n_409),
.B2(n_367),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_605),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_584),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_604),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_679),
.B(n_652),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_653),
.A2(n_667),
.B(n_660),
.C(n_677),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_666),
.Y(n_709)
);

BUFx12f_ASAP7_75t_L g710 ( 
.A(n_695),
.Y(n_710)
);

INVxp33_ASAP7_75t_SL g711 ( 
.A(n_658),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_661),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_663),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_660),
.A2(n_703),
.B1(n_699),
.B2(n_650),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_655),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_SL g716 ( 
.A(n_702),
.B(n_669),
.C(n_676),
.Y(n_716)
);

AO21x2_ASAP7_75t_L g717 ( 
.A1(n_693),
.A2(n_683),
.B(n_689),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_656),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_706),
.B(n_668),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_662),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_664),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_702),
.A2(n_667),
.B(n_651),
.C(n_696),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_674),
.B(n_675),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_705),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_690),
.Y(n_725)
);

INVxp33_ASAP7_75t_L g726 ( 
.A(n_690),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_673),
.B(n_704),
.Y(n_727)
);

OA21x2_ASAP7_75t_L g728 ( 
.A1(n_691),
.A2(n_687),
.B(n_649),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_665),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_684),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_682),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_688),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_697),
.B(n_704),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_673),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_680),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_735),
.B(n_685),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_731),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_714),
.A2(n_699),
.B1(n_650),
.B2(n_677),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_707),
.B(n_692),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_727),
.B(n_685),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_727),
.B(n_685),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_649),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_707),
.B(n_654),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_720),
.B(n_685),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_710),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_725),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_711),
.B(n_701),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_729),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_729),
.Y(n_749)
);

NOR2x1_ASAP7_75t_L g750 ( 
.A(n_729),
.B(n_686),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_721),
.B(n_659),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_719),
.B(n_700),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_721),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_737),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_743),
.B(n_728),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_739),
.B(n_728),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_739),
.B(n_728),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_750),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_740),
.B(n_709),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_747),
.B(n_686),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_736),
.B(n_717),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_742),
.B(n_724),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_749),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_740),
.B(n_741),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_756),
.B(n_752),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_754),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_754),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_760),
.B(n_657),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_764),
.B(n_741),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_756),
.B(n_752),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_759),
.B(n_753),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_763),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_759),
.B(n_753),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_762),
.B(n_751),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_764),
.B(n_744),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_766),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_765),
.B(n_755),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_765),
.B(n_755),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_766),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_767),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_767),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_774),
.B(n_757),
.Y(n_782)
);

AOI222xp33_ASAP7_75t_L g783 ( 
.A1(n_771),
.A2(n_733),
.B1(n_715),
.B2(n_723),
.C1(n_672),
.C2(n_757),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_775),
.B(n_761),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_775),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_785),
.Y(n_786)
);

NOR2x1_ASAP7_75t_L g787 ( 
.A(n_784),
.B(n_763),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_784),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_779),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_779),
.B(n_772),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_776),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_782),
.B(n_770),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_783),
.A2(n_716),
.B1(n_773),
.B2(n_768),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_777),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_777),
.A2(n_769),
.B1(n_763),
.B2(n_738),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_780),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_781),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_795),
.B(n_778),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_787),
.B(n_748),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_788),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_795),
.B(n_778),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_789),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_800),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_798),
.B(n_786),
.Y(n_804)
);

AOI221x1_ASAP7_75t_L g805 ( 
.A1(n_801),
.A2(n_802),
.B1(n_797),
.B2(n_791),
.C(n_790),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_803),
.B(n_793),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_804),
.Y(n_807)
);

NOR2x1_ASAP7_75t_SL g808 ( 
.A(n_806),
.B(n_710),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_807),
.B(n_794),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_809),
.B(n_805),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_808),
.B(n_701),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_SL g812 ( 
.A(n_811),
.B(n_678),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_810),
.Y(n_813)
);

NAND2x1_ASAP7_75t_SL g814 ( 
.A(n_813),
.B(n_809),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_812),
.A2(n_694),
.B1(n_745),
.B2(n_671),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_813),
.B(n_698),
.C(n_670),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_814),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_815),
.B(n_718),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_816),
.A2(n_799),
.B1(n_792),
.B2(n_730),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_815),
.B(n_712),
.Y(n_820)
);

NOR2x1_ASAP7_75t_L g821 ( 
.A(n_816),
.B(n_688),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_817),
.A2(n_672),
.B(n_799),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_818),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_820),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_821),
.A2(n_792),
.B1(n_746),
.B2(n_790),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_819),
.B(n_796),
.Y(n_826)
);

AOI21xp33_ASAP7_75t_L g827 ( 
.A1(n_817),
.A2(n_726),
.B(n_681),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_820),
.A2(n_713),
.B1(n_712),
.B2(n_750),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_824),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_823),
.B(n_713),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_827),
.A2(n_751),
.B(n_722),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_822),
.A2(n_708),
.B(n_758),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_829),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_832),
.B(n_826),
.Y(n_834)
);

OAI211xp5_ASAP7_75t_L g835 ( 
.A1(n_833),
.A2(n_828),
.B(n_831),
.C(n_830),
.Y(n_835)
);

NAND2xp67_ASAP7_75t_L g836 ( 
.A(n_835),
.B(n_834),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_836),
.A2(n_825),
.B1(n_732),
.B2(n_746),
.Y(n_837)
);


endmodule