module fake_jpeg_10672_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_71),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_50),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_0),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_78),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_0),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_66),
.C(n_49),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_95),
.C(n_11),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_86),
.Y(n_111)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_42),
.B1(n_43),
.B2(n_61),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_97),
.B1(n_100),
.B2(n_58),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_65),
.B1(n_56),
.B2(n_60),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_3),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_63),
.B(n_62),
.C(n_58),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_62),
.B1(n_51),
.B2(n_53),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_51),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_105),
.B1(n_106),
.B2(n_115),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_98),
.B(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_114),
.C(n_117),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_47),
.B1(n_5),
.B2(n_7),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_10),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_112),
.B1(n_116),
.B2(n_118),
.Y(n_124)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_103),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_125),
.A2(n_126),
.B(n_120),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_121),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_115),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_120),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_113),
.B(n_119),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_122),
.C(n_110),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_111),
.B(n_108),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_18),
.B(n_19),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_111),
.B(n_22),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_21),
.C(n_23),
.Y(n_140)
);

OAI221xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_124),
.B1(n_27),
.B2(n_30),
.C(n_31),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_25),
.Y(n_142)
);


endmodule