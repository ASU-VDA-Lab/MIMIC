module fake_jpeg_17574_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_43),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_3),
.Y(n_87)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_40),
.B1(n_45),
.B2(n_44),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_39),
.Y(n_80)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_51),
.B1(n_46),
.B2(n_48),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_75),
.B1(n_85),
.B2(n_67),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_46),
.B1(n_25),
.B2(n_26),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_4),
.B(n_5),
.Y(n_92)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_85),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_73),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_94),
.B1(n_68),
.B2(n_63),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_7),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_6),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_9),
.Y(n_102)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_78),
.C(n_64),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_91),
.C(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_102),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_105),
.B(n_12),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_88),
.B(n_98),
.C(n_97),
.D(n_89),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_109),
.B(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

OAI21x1_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_14),
.B(n_16),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_108),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_116),
.A2(n_117),
.B(n_19),
.Y(n_118)
);

NAND2x1p5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_18),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.C(n_21),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_112),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_22),
.B(n_27),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_28),
.C(n_29),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_30),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_31),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_33),
.Y(n_127)
);


endmodule