module fake_netlist_1_6769_n_907 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_907);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_907;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_522;
wire n_264;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_91), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_78), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_84), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_44), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_51), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_89), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_55), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_90), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_66), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_34), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_22), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_57), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_81), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_10), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_86), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_105), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_85), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_31), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_56), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_21), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_14), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_82), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_80), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_34), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_45), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_21), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_1), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_35), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_52), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_22), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_20), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_20), .Y(n_138) );
INVx1_ASAP7_75t_SL g139 ( .A(n_92), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_7), .Y(n_140) );
INVx2_ASAP7_75t_SL g141 ( .A(n_31), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_49), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_75), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_38), .Y(n_144) );
BUFx10_ASAP7_75t_L g145 ( .A(n_62), .Y(n_145) );
BUFx10_ASAP7_75t_L g146 ( .A(n_50), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_71), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_39), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_101), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_6), .Y(n_150) );
INVx5_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_141), .B(n_0), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
BUFx12f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_144), .B(n_40), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_116), .B(n_0), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_116), .B(n_1), .Y(n_160) );
BUFx8_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_141), .B(n_2), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_145), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_127), .B(n_2), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_145), .B(n_3), .Y(n_170) );
INVx5_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_140), .B(n_3), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_127), .B(n_4), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_141), .B(n_4), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_153), .A2(n_174), .B1(n_164), .B2(n_156), .Y(n_175) );
OR2x6_ASAP7_75t_L g176 ( .A(n_159), .B(n_115), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_153), .A2(n_115), .B1(n_117), .B2(n_120), .Y(n_177) );
AO22x2_ASAP7_75t_L g178 ( .A1(n_172), .A2(n_159), .B1(n_160), .B2(n_170), .Y(n_178) );
AO22x2_ASAP7_75t_L g179 ( .A1(n_172), .A2(n_123), .B1(n_111), .B2(n_112), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_172), .Y(n_180) );
OR2x6_ASAP7_75t_L g181 ( .A(n_159), .B(n_160), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_165), .B(n_145), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
OAI22xp33_ASAP7_75t_SL g184 ( .A1(n_170), .A2(n_126), .B1(n_134), .B2(n_133), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_156), .B(n_118), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_165), .B(n_146), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_165), .B(n_146), .Y(n_188) );
AO22x2_ASAP7_75t_L g189 ( .A1(n_172), .A2(n_123), .B1(n_111), .B2(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_165), .B(n_146), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_159), .A2(n_121), .B1(n_129), .B2(n_124), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_154), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_156), .A2(n_121), .B1(n_129), .B2(n_136), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_137), .B1(n_132), .B2(n_138), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_160), .B(n_146), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_153), .A2(n_117), .B1(n_120), .B2(n_150), .Y(n_198) );
AO22x2_ASAP7_75t_L g199 ( .A1(n_172), .A2(n_174), .B1(n_164), .B2(n_155), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_156), .A2(n_140), .B1(n_150), .B2(n_130), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_166), .B(n_108), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_166), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_169), .A2(n_150), .B1(n_130), .B2(n_125), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_166), .A2(n_130), .B1(n_108), .B2(n_112), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_154), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_166), .B(n_146), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_169), .A2(n_122), .B1(n_113), .B2(n_142), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_152), .B(n_139), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_173), .A2(n_122), .B1(n_113), .B2(n_125), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_155), .B(n_131), .Y(n_212) );
AO22x2_ASAP7_75t_L g213 ( .A1(n_172), .A2(n_131), .B1(n_139), .B2(n_7), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_152), .B(n_106), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_152), .B(n_107), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_161), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_172), .B(n_109), .Y(n_218) );
NAND3x1_ASAP7_75t_L g219 ( .A(n_173), .B(n_5), .C(n_6), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_149), .B1(n_147), .B2(n_135), .Y(n_221) );
XNOR2xp5_ASAP7_75t_L g222 ( .A(n_192), .B(n_174), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_202), .B(n_180), .Y(n_223) );
INVxp67_ASAP7_75t_SL g224 ( .A(n_196), .Y(n_224) );
XOR2xp5_ASAP7_75t_L g225 ( .A(n_192), .B(n_194), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_197), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_197), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_180), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_181), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
XOR2xp5_ASAP7_75t_L g233 ( .A(n_195), .B(n_178), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_181), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_199), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_190), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_206), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_181), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_190), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_179), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_181), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_176), .B(n_151), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_179), .Y(n_246) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_220), .A2(n_163), .B(n_162), .Y(n_247) );
XNOR2xp5_ASAP7_75t_L g248 ( .A(n_195), .B(n_5), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_176), .Y(n_249) );
XOR2xp5_ASAP7_75t_L g250 ( .A(n_178), .B(n_8), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_176), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_206), .B(n_161), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
NOR2xp33_ASAP7_75t_SL g255 ( .A(n_216), .B(n_157), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_183), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_185), .B(n_161), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_209), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_209), .B(n_161), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_178), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_178), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_182), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_187), .B(n_151), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_188), .Y(n_267) );
BUFx8_ASAP7_75t_L g268 ( .A(n_188), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_179), .B(n_162), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_191), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_214), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_191), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_189), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_221), .Y(n_274) );
NOR2xp67_ASAP7_75t_L g275 ( .A(n_207), .B(n_151), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_175), .A2(n_155), .B(n_162), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_189), .Y(n_278) );
XOR2xp5_ASAP7_75t_L g279 ( .A(n_189), .B(n_9), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_218), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_201), .B(n_161), .Y(n_281) );
BUFx2_ASAP7_75t_R g282 ( .A(n_213), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_218), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_200), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_215), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_234), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_234), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_226), .B(n_177), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
INVx3_ASAP7_75t_SL g292 ( .A(n_269), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_269), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_222), .B(n_221), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_269), .B(n_213), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_227), .B(n_213), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_245), .B(n_204), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_284), .B(n_198), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_245), .B(n_213), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_247), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_236), .B(n_207), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_230), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_247), .Y(n_303) );
AND2x2_ASAP7_75t_SL g304 ( .A(n_242), .B(n_154), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_259), .B(n_211), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_280), .B(n_211), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_283), .B(n_203), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_268), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_228), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_263), .B(n_203), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_242), .B(n_184), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_223), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_277), .A2(n_212), .B(n_186), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_265), .B(n_161), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_236), .B(n_151), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_228), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_249), .B(n_151), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_251), .B(n_151), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_252), .B(n_151), .Y(n_319) );
AND2x6_ASAP7_75t_L g320 ( .A(n_244), .B(n_154), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_240), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_279), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_240), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_244), .B(n_151), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_237), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_246), .B(n_151), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_261), .B(n_157), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_246), .B(n_151), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_237), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_267), .B(n_155), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_270), .B(n_155), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_272), .B(n_155), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_262), .B(n_275), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_222), .B(n_9), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_241), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_286), .B(n_157), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_241), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_230), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_260), .A2(n_193), .B(n_186), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_266), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_292), .B(n_233), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_326), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_326), .Y(n_345) );
BUFx5_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
BUFx5_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_301), .B(n_229), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_291), .B(n_231), .Y(n_350) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_292), .B(n_291), .Y(n_351) );
NAND2x1_ASAP7_75t_L g352 ( .A(n_320), .B(n_157), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_292), .B(n_233), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_301), .B(n_250), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_301), .B(n_250), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_320), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_330), .B(n_232), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_338), .B(n_235), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_330), .B(n_268), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_300), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_336), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_291), .B(n_273), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_291), .Y(n_364) );
BUFx4f_ASAP7_75t_L g365 ( .A(n_320), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_300), .Y(n_367) );
INVx6_ASAP7_75t_L g368 ( .A(n_321), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_321), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_320), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_293), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_338), .B(n_235), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_373), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_373), .B(n_293), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_349), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_354), .A2(n_279), .B1(n_243), .B2(n_225), .Y(n_379) );
NOR2xp67_ASAP7_75t_SL g380 ( .A(n_349), .B(n_293), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_354), .A2(n_225), .B1(n_335), .B2(n_323), .Y(n_381) );
BUFx2_ASAP7_75t_R g382 ( .A(n_360), .Y(n_382) );
INVx6_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g384 ( .A(n_351), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_368), .Y(n_385) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_342), .Y(n_386) );
BUFx12f_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_365), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
INVx6_ASAP7_75t_L g390 ( .A(n_368), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_351), .B(n_308), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
BUFx2_ASAP7_75t_SL g393 ( .A(n_342), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_344), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_359), .B(n_338), .Y(n_395) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_358), .Y(n_396) );
AO21x1_ASAP7_75t_L g397 ( .A1(n_358), .A2(n_295), .B(n_296), .Y(n_397) );
NOR2x1_ASAP7_75t_SL g398 ( .A(n_349), .B(n_295), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_358), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_359), .B(n_297), .Y(n_401) );
INVx8_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_349), .Y(n_403) );
BUFx8_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_375), .B(n_295), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_376), .B(n_358), .Y(n_406) );
INVx6_ASAP7_75t_L g407 ( .A(n_404), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_395), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_386), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_404), .A2(n_355), .B1(n_354), .B2(n_323), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_379), .A2(n_282), .B1(n_335), .B2(n_355), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_396), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_404), .A2(n_355), .B1(n_335), .B2(n_294), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_404), .A2(n_353), .B1(n_343), .B2(n_243), .Y(n_414) );
INVx4_ASAP7_75t_L g415 ( .A(n_384), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_395), .B(n_388), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_402), .A2(n_294), .B1(n_353), .B2(n_343), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_386), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_402), .A2(n_343), .B1(n_353), .B2(n_375), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_396), .B(n_400), .Y(n_424) );
INVx6_ASAP7_75t_L g425 ( .A(n_402), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_386), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_387), .Y(n_428) );
BUFx8_ASAP7_75t_SL g429 ( .A(n_387), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_379), .A2(n_248), .B(n_296), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_395), .A2(n_367), .B1(n_294), .B2(n_365), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_378), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_402), .A2(n_367), .B1(n_365), .B2(n_248), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_382), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_402), .A2(n_311), .B1(n_299), .B2(n_296), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_402), .Y(n_439) );
OAI22x1_ASAP7_75t_L g440 ( .A1(n_377), .A2(n_274), .B1(n_361), .B2(n_308), .Y(n_440) );
BUFx12f_ASAP7_75t_L g441 ( .A(n_377), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_378), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_381), .A2(n_311), .B1(n_299), .B2(n_348), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_388), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_401), .A2(n_365), .B1(n_299), .B2(n_348), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_401), .A2(n_334), .B1(n_360), .B2(n_297), .Y(n_447) );
INVx8_ASAP7_75t_L g448 ( .A(n_385), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_378), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_378), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_424), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_411), .A2(n_405), .B1(n_397), .B2(n_334), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_411), .A2(n_274), .B1(n_306), .B2(n_305), .C1(n_307), .C2(n_310), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_430), .A2(n_405), .B1(n_397), .B2(n_334), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_421), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_407), .A2(n_393), .B1(n_398), .B2(n_405), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_430), .A2(n_334), .B1(n_350), .B2(n_391), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_413), .A2(n_334), .B1(n_350), .B2(n_363), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_444), .B(n_344), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_413), .A2(n_350), .B1(n_363), .B2(n_393), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_421), .B(n_388), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_436), .A2(n_350), .B1(n_363), .B2(n_268), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_424), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_441), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_432), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_441), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_432), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_424), .B(n_398), .Y(n_470) );
CKINVDCx11_ASAP7_75t_R g471 ( .A(n_439), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_409), .B(n_382), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_406), .B(n_361), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_436), .A2(n_350), .B1(n_363), .B2(n_347), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_444), .B(n_345), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_443), .B(n_345), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_423), .A2(n_363), .B1(n_346), .B2(n_347), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_443), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_439), .A2(n_239), .B1(n_377), .B2(n_219), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_423), .A2(n_347), .B1(n_346), .B2(n_297), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_410), .A2(n_347), .B1(n_346), .B2(n_297), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_412), .B(n_361), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_410), .A2(n_347), .B1(n_346), .B2(n_297), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_412), .Y(n_484) );
INVx1_ASAP7_75t_SL g485 ( .A(n_429), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_414), .A2(n_239), .B1(n_377), .B2(n_219), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_418), .A2(n_407), .B1(n_425), .B2(n_446), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_418), .A2(n_347), .B1(n_346), .B2(n_364), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_407), .A2(n_347), .B1(n_346), .B2(n_364), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g491 ( .A1(n_437), .A2(n_302), .B1(n_339), .B2(n_389), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_407), .A2(n_339), .B1(n_302), .B2(n_346), .Y(n_492) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_415), .B(n_388), .Y(n_493) );
OAI21xp5_ASAP7_75t_SL g494 ( .A1(n_417), .A2(n_328), .B(n_349), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_407), .A2(n_389), .B1(n_352), .B2(n_364), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g496 ( .A1(n_407), .A2(n_389), .B1(n_352), .B2(n_362), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_420), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_427), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_427), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_441), .A2(n_346), .B1(n_347), .B2(n_389), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_426), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_427), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_406), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_406), .Y(n_504) );
OAI21xp33_ASAP7_75t_L g505 ( .A1(n_426), .A2(n_163), .B(n_162), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_425), .A2(n_374), .B1(n_372), .B2(n_362), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_433), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_425), .A2(n_346), .B1(n_347), .B2(n_374), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_433), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_426), .Y(n_510) );
AOI22xp5_ASAP7_75t_SL g511 ( .A1(n_428), .A2(n_356), .B1(n_371), .B2(n_349), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_425), .A2(n_347), .B1(n_346), .B2(n_374), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_425), .A2(n_347), .B1(n_346), .B2(n_341), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_408), .B(n_361), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_425), .A2(n_372), .B1(n_304), .B2(n_356), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_433), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_435), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_428), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_447), .A2(n_304), .B1(n_366), .B2(n_371), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_428), .Y(n_520) );
INVx4_ASAP7_75t_L g521 ( .A(n_434), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_434), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_454), .A2(n_415), .B1(n_419), .B2(n_431), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_486), .A2(n_446), .B1(n_431), .B2(n_438), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_479), .A2(n_438), .B1(n_440), .B2(n_434), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_451), .B(n_408), .Y(n_526) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_468), .A2(n_419), .B1(n_415), .B2(n_445), .Y(n_527) );
OAI221xp5_ASAP7_75t_L g528 ( .A1(n_464), .A2(n_306), .B1(n_307), .B2(n_305), .C(n_310), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_487), .A2(n_419), .B1(n_415), .B2(n_440), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_456), .A2(n_419), .B1(n_416), .B2(n_408), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_468), .A2(n_417), .B1(n_416), .B2(n_408), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_481), .A2(n_408), .B1(n_416), .B2(n_429), .Y(n_532) );
OAI222xp33_ASAP7_75t_L g533 ( .A1(n_468), .A2(n_417), .B1(n_416), .B2(n_445), .C1(n_380), .C2(n_352), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_483), .A2(n_416), .B1(n_417), .B2(n_445), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_455), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_459), .A2(n_445), .B1(n_390), .B2(n_383), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_480), .A2(n_445), .B1(n_448), .B2(n_390), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_470), .A2(n_448), .B1(n_390), .B2(n_383), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_451), .B(n_448), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_470), .A2(n_448), .B1(n_390), .B2(n_383), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_467), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_470), .A2(n_448), .B1(n_390), .B2(n_383), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_465), .A2(n_474), .B1(n_462), .B2(n_477), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_455), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_465), .B(n_448), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_460), .A2(n_399), .B1(n_385), .B2(n_347), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_488), .A2(n_399), .B1(n_385), .B2(n_347), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_499), .B(n_435), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_453), .B(n_341), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_503), .B(n_341), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_492), .A2(n_493), .B1(n_475), .B2(n_461), .Y(n_551) );
OAI221xp5_ASAP7_75t_SL g552 ( .A1(n_485), .A2(n_298), .B1(n_163), .B2(n_290), .C(n_278), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_491), .A2(n_346), .B1(n_368), .B2(n_369), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_463), .A2(n_370), .B1(n_369), .B2(n_312), .Y(n_554) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_466), .A2(n_356), .B1(n_366), .B2(n_371), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_458), .A2(n_370), .B1(n_369), .B2(n_312), .Y(n_556) );
OAI222xp33_ASAP7_75t_L g557 ( .A1(n_520), .A2(n_521), .B1(n_466), .B2(n_510), .C1(n_457), .C2(n_518), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_520), .A2(n_356), .B1(n_366), .B2(n_371), .Y(n_558) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_499), .A2(n_442), .B(n_435), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_506), .A2(n_369), .B1(n_370), .B2(n_312), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_467), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_471), .A2(n_370), .B1(n_369), .B2(n_285), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_469), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_520), .A2(n_357), .B1(n_276), .B2(n_285), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_471), .A2(n_370), .B1(n_157), .B2(n_357), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_522), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_503), .A2(n_157), .B1(n_271), .B2(n_264), .Y(n_567) );
OAI221xp5_ASAP7_75t_SL g568 ( .A1(n_494), .A2(n_298), .B1(n_163), .B2(n_290), .C(n_238), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_521), .A2(n_371), .B1(n_356), .B2(n_366), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_521), .A2(n_366), .B1(n_356), .B2(n_371), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_504), .B(n_442), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_501), .A2(n_371), .B1(n_356), .B2(n_366), .Y(n_572) );
OAI221xp5_ASAP7_75t_SL g573 ( .A1(n_505), .A2(n_472), .B1(n_513), .B2(n_489), .C(n_501), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_504), .A2(n_157), .B1(n_271), .B2(n_264), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_502), .B(n_442), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_511), .A2(n_403), .B1(n_392), .B2(n_378), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_469), .B(n_449), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_478), .B(n_10), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_500), .A2(n_449), .B1(n_300), .B2(n_303), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_508), .A2(n_303), .B1(n_449), .B2(n_392), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_478), .B(n_11), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_496), .A2(n_403), .B1(n_392), .B2(n_450), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_473), .A2(n_403), .B1(n_392), .B2(n_450), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_484), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_490), .A2(n_157), .B1(n_328), .B2(n_450), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_495), .B(n_392), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_484), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_512), .A2(n_303), .B1(n_420), .B2(n_450), .Y(n_588) );
AOI21xp5_ASAP7_75t_SL g589 ( .A1(n_515), .A2(n_403), .B(n_392), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_502), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_490), .B(n_11), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_476), .B(n_12), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_519), .A2(n_157), .B1(n_328), .B2(n_450), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_514), .A2(n_157), .B1(n_328), .B2(n_450), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_473), .A2(n_238), .B1(n_303), .B2(n_328), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_482), .B(n_167), .C(n_168), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_514), .A2(n_157), .B1(n_420), .B2(n_450), .Y(n_597) );
AND2x2_ASAP7_75t_SL g598 ( .A(n_498), .B(n_420), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_498), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_482), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_507), .B(n_12), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_507), .A2(n_157), .B1(n_420), .B2(n_403), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_509), .A2(n_516), .B1(n_157), .B2(n_517), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_509), .A2(n_420), .B1(n_403), .B2(n_380), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_516), .A2(n_403), .B1(n_223), .B2(n_314), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_517), .A2(n_167), .B1(n_321), .B2(n_315), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_497), .A2(n_320), .B1(n_154), .B2(n_158), .Y(n_607) );
OAI22xp5_ASAP7_75t_SL g608 ( .A1(n_497), .A2(n_337), .B1(n_287), .B2(n_288), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_497), .A2(n_167), .B1(n_315), .B2(n_329), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_497), .A2(n_167), .B1(n_315), .B2(n_329), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_497), .B(n_13), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_454), .A2(n_167), .B1(n_288), .B2(n_287), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_454), .A2(n_167), .B1(n_320), .B2(n_257), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_467), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_455), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_451), .B(n_13), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_454), .A2(n_167), .B1(n_320), .B2(n_309), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_452), .A2(n_316), .B1(n_253), .B2(n_332), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_454), .A2(n_167), .B1(n_320), .B2(n_316), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g620 ( .A1(n_551), .A2(n_331), .B1(n_332), .B2(n_333), .C(n_319), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_566), .B(n_14), .Y(n_621) );
AND2x2_ASAP7_75t_SL g622 ( .A(n_590), .B(n_255), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_600), .B(n_15), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_573), .A2(n_167), .B1(n_158), .B2(n_168), .C(n_171), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_557), .A2(n_168), .B(n_171), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_527), .B(n_158), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_600), .B(n_15), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_526), .B(n_167), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_526), .B(n_158), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_541), .B(n_16), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_541), .B(n_561), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_561), .B(n_16), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_548), .B(n_158), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_523), .A2(n_158), .B1(n_168), .B2(n_171), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_578), .B(n_17), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_563), .B(n_17), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_563), .B(n_18), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_614), .B(n_18), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_614), .B(n_19), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_575), .B(n_158), .Y(n_641) );
OA21x2_ASAP7_75t_L g642 ( .A1(n_586), .A2(n_313), .B(n_340), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_592), .B(n_158), .C(n_168), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_590), .B(n_19), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_524), .B(n_23), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_539), .B(n_23), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_545), .B(n_24), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_524), .B(n_24), .Y(n_648) );
OAI221xp5_ASAP7_75t_SL g649 ( .A1(n_525), .A2(n_331), .B1(n_333), .B2(n_317), .C(n_318), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_616), .B(n_25), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_525), .A2(n_110), .B1(n_128), .B2(n_119), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_582), .B(n_168), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_575), .B(n_25), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_599), .B(n_26), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_599), .B(n_26), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g656 ( .A1(n_533), .A2(n_281), .B(n_28), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_576), .B(n_168), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_571), .B(n_27), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_535), .B(n_27), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_535), .B(n_28), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_581), .B(n_29), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_529), .B(n_29), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_596), .B(n_168), .C(n_171), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_544), .B(n_30), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_591), .B(n_30), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_544), .B(n_32), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_543), .B(n_32), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_584), .B(n_33), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g669 ( .A(n_552), .B(n_313), .C(n_114), .Y(n_669) );
AOI21xp5_ASAP7_75t_SL g670 ( .A1(n_531), .A2(n_33), .B(n_35), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_584), .B(n_36), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_587), .B(n_36), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_568), .B(n_37), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_587), .B(n_37), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g675 ( .A1(n_612), .A2(n_317), .B1(n_319), .B2(n_318), .C(n_316), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_615), .B(n_168), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_534), .A2(n_168), .B1(n_171), .B2(n_316), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_618), .A2(n_171), .B1(n_327), .B2(n_325), .Y(n_678) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_598), .B(n_289), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_615), .B(n_171), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g681 ( .A1(n_530), .A2(n_340), .B(n_327), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_601), .B(n_171), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_550), .B(n_171), .Y(n_683) );
OA21x2_ASAP7_75t_L g684 ( .A1(n_604), .A2(n_193), .B(n_205), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_577), .B(n_325), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_611), .A2(n_319), .B(n_318), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_549), .B(n_317), .Y(n_687) );
OAI21xp33_ASAP7_75t_SL g688 ( .A1(n_598), .A2(n_224), .B(n_42), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_596), .B(n_324), .C(n_322), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_564), .B(n_41), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_559), .B(n_43), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_532), .B(n_46), .Y(n_692) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_556), .A2(n_324), .B(n_322), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_559), .B(n_47), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_559), .B(n_48), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_559), .B(n_53), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_603), .B(n_324), .C(n_322), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_565), .B(n_324), .C(n_322), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_583), .B(n_54), .Y(n_699) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_553), .B(n_324), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_560), .B(n_58), .Y(n_701) );
NOR2xp33_ASAP7_75t_SL g702 ( .A(n_608), .B(n_324), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_538), .B(n_59), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_589), .B(n_60), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_608), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_589), .B(n_61), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_540), .B(n_63), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_542), .B(n_64), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_536), .A2(n_324), .B(n_322), .C(n_289), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_537), .B(n_65), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_562), .B(n_254), .C(n_217), .D(n_210), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_597), .B(n_322), .C(n_289), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_580), .B(n_67), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_617), .B(n_546), .C(n_619), .D(n_594), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_605), .B(n_68), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_585), .B(n_322), .C(n_289), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_605), .B(n_69), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_595), .B(n_580), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_602), .B(n_289), .C(n_208), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_632), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_656), .B(n_593), .C(n_579), .Y(n_721) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_670), .A2(n_554), .B(n_613), .C(n_558), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_624), .B(n_588), .Y(n_723) );
AO21x2_ASAP7_75t_L g724 ( .A1(n_694), .A2(n_555), .B(n_570), .Y(n_724) );
NAND4xp75_ASAP7_75t_L g725 ( .A(n_667), .B(n_595), .C(n_569), .D(n_547), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_705), .A2(n_528), .B1(n_567), .B2(n_574), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_653), .Y(n_727) );
AO21x2_ASAP7_75t_L g728 ( .A1(n_696), .A2(n_572), .B(n_205), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_667), .A2(n_606), .B1(n_609), .B2(n_610), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_653), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_624), .B(n_607), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_630), .B(n_70), .Y(n_732) );
AND2x4_ASAP7_75t_SL g733 ( .A(n_630), .B(n_289), .Y(n_733) );
NAND4xp75_ASAP7_75t_L g734 ( .A(n_688), .B(n_72), .C(n_73), .D(n_74), .Y(n_734) );
AO21x2_ASAP7_75t_L g735 ( .A1(n_644), .A2(n_208), .B(n_258), .Y(n_735) );
AND2x4_ASAP7_75t_L g736 ( .A(n_704), .B(n_76), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_655), .B(n_77), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_714), .A2(n_240), .B1(n_256), .B2(n_258), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_627), .A2(n_240), .B(n_83), .Y(n_739) );
BUFx3_ASAP7_75t_L g740 ( .A(n_634), .Y(n_740) );
OAI211xp5_ASAP7_75t_SL g741 ( .A1(n_645), .A2(n_79), .B(n_87), .C(n_88), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_655), .B(n_93), .Y(n_742) );
OAI21xp33_ASAP7_75t_SL g743 ( .A1(n_679), .A2(n_94), .B(n_95), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_625), .B(n_648), .C(n_621), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_659), .Y(n_745) );
AO21x2_ASAP7_75t_L g746 ( .A1(n_691), .A2(n_96), .B(n_97), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_643), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_651), .B(n_102), .C(n_103), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_704), .B(n_104), .Y(n_749) );
NAND4xp75_ASAP7_75t_L g750 ( .A(n_622), .B(n_700), .C(n_662), .D(n_652), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_620), .B(n_649), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_659), .B(n_660), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_642), .B(n_691), .Y(n_753) );
AO21x2_ASAP7_75t_L g754 ( .A1(n_695), .A2(n_668), .B(n_672), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_642), .B(n_695), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_660), .Y(n_756) );
OAI211xp5_ASAP7_75t_SL g757 ( .A1(n_650), .A2(n_665), .B(n_635), .C(n_636), .Y(n_757) );
INVx2_ASAP7_75t_SL g758 ( .A(n_679), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_661), .B(n_702), .C(n_709), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g760 ( .A(n_661), .B(n_636), .C(n_693), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_658), .B(n_623), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_634), .B(n_641), .Y(n_762) );
NAND4xp25_ASAP7_75t_L g763 ( .A(n_673), .B(n_626), .C(n_718), .D(n_646), .Y(n_763) );
NAND4xp75_ASAP7_75t_L g764 ( .A(n_622), .B(n_700), .C(n_652), .D(n_657), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_628), .B(n_631), .C(n_633), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_664), .B(n_671), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_641), .B(n_671), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_647), .A2(n_637), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_654), .B(n_692), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_674), .B(n_686), .Y(n_770) );
AOI211xp5_ASAP7_75t_SL g771 ( .A1(n_706), .A2(n_699), .B(n_675), .C(n_681), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g772 ( .A(n_657), .B(n_689), .C(n_663), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_664), .Y(n_773) );
NAND4xp75_ASAP7_75t_L g774 ( .A(n_706), .B(n_699), .C(n_710), .D(n_666), .Y(n_774) );
NAND4xp75_ASAP7_75t_L g775 ( .A(n_666), .B(n_713), .C(n_680), .D(n_690), .Y(n_775) );
AO21x2_ASAP7_75t_L g776 ( .A1(n_715), .A2(n_717), .B(n_713), .Y(n_776) );
AO21x2_ASAP7_75t_L g777 ( .A1(n_676), .A2(n_682), .B(n_707), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_676), .B(n_684), .Y(n_778) );
INVx3_ASAP7_75t_L g779 ( .A(n_684), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_712), .B(n_698), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_669), .A2(n_677), .B1(n_708), .B2(n_703), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_711), .B(n_701), .C(n_683), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_685), .B(n_687), .Y(n_783) );
OA211x2_ASAP7_75t_L g784 ( .A1(n_716), .A2(n_697), .B(n_719), .C(n_678), .Y(n_784) );
NOR3xp33_ASAP7_75t_L g785 ( .A(n_656), .B(n_667), .C(n_625), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_632), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_656), .B(n_667), .C(n_705), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_632), .B(n_451), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_629), .B(n_653), .Y(n_789) );
AO21x2_ASAP7_75t_L g790 ( .A1(n_694), .A2(n_696), .B(n_644), .Y(n_790) );
NAND4xp75_ASAP7_75t_L g791 ( .A(n_784), .B(n_743), .C(n_751), .D(n_768), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_740), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_720), .Y(n_793) );
INVxp67_ASAP7_75t_L g794 ( .A(n_761), .Y(n_794) );
NAND3xp33_ASAP7_75t_L g795 ( .A(n_787), .B(n_771), .C(n_760), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_740), .Y(n_796) );
BUFx2_ASAP7_75t_L g797 ( .A(n_762), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_786), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_788), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_727), .B(n_730), .Y(n_800) );
NOR4xp25_ASAP7_75t_L g801 ( .A(n_757), .B(n_761), .C(n_763), .D(n_759), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_751), .A2(n_785), .B1(n_725), .B2(n_774), .Y(n_802) );
NAND4xp75_ASAP7_75t_L g803 ( .A(n_769), .B(n_731), .C(n_753), .D(n_755), .Y(n_803) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_780), .Y(n_804) );
XNOR2x2_ASAP7_75t_L g805 ( .A(n_764), .B(n_750), .Y(n_805) );
NAND4xp75_ASAP7_75t_L g806 ( .A(n_769), .B(n_731), .C(n_755), .D(n_753), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_744), .A2(n_721), .B1(n_782), .B2(n_770), .Y(n_807) );
AND2x4_ASAP7_75t_L g808 ( .A(n_758), .B(n_723), .Y(n_808) );
XOR2x2_ASAP7_75t_L g809 ( .A(n_775), .B(n_734), .Y(n_809) );
NAND4xp75_ASAP7_75t_L g810 ( .A(n_758), .B(n_770), .C(n_723), .D(n_780), .Y(n_810) );
CKINVDCx8_ASAP7_75t_R g811 ( .A(n_736), .Y(n_811) );
INVx2_ASAP7_75t_SL g812 ( .A(n_733), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_733), .Y(n_813) );
BUFx2_ASAP7_75t_L g814 ( .A(n_767), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_789), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_745), .B(n_773), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_756), .Y(n_817) );
AND2x4_ASAP7_75t_L g818 ( .A(n_790), .B(n_754), .Y(n_818) );
XOR2x2_ASAP7_75t_L g819 ( .A(n_783), .B(n_765), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_752), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_754), .B(n_790), .Y(n_821) );
AND2x4_ASAP7_75t_L g822 ( .A(n_790), .B(n_754), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_777), .B(n_766), .Y(n_823) );
XOR2x2_ASAP7_75t_L g824 ( .A(n_736), .B(n_749), .Y(n_824) );
INVx2_ASAP7_75t_SL g825 ( .A(n_778), .Y(n_825) );
NAND4xp75_ASAP7_75t_L g826 ( .A(n_737), .B(n_742), .C(n_739), .D(n_722), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_777), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g828 ( .A(n_726), .B(n_781), .Y(n_828) );
XOR2x2_ASAP7_75t_L g829 ( .A(n_749), .B(n_772), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_797), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_808), .B(n_777), .Y(n_831) );
XOR2x2_ASAP7_75t_L g832 ( .A(n_802), .B(n_748), .Y(n_832) );
XOR2x2_ASAP7_75t_L g833 ( .A(n_805), .B(n_746), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_793), .Y(n_834) );
XNOR2xp5_ASAP7_75t_L g835 ( .A(n_824), .B(n_738), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_798), .Y(n_836) );
XOR2x2_ASAP7_75t_L g837 ( .A(n_791), .B(n_776), .Y(n_837) );
XNOR2xp5_ASAP7_75t_L g838 ( .A(n_824), .B(n_729), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_816), .Y(n_839) );
XNOR2x1_ASAP7_75t_L g840 ( .A(n_828), .B(n_732), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_792), .Y(n_841) );
XOR2x2_ASAP7_75t_L g842 ( .A(n_819), .B(n_776), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_808), .B(n_724), .Y(n_843) );
XNOR2x1_ASAP7_75t_L g844 ( .A(n_795), .B(n_779), .Y(n_844) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_827), .Y(n_845) );
XNOR2x1_ASAP7_75t_L g846 ( .A(n_819), .B(n_776), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_807), .A2(n_735), .B1(n_741), .B2(n_724), .Y(n_847) );
INVx1_ASAP7_75t_SL g848 ( .A(n_792), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_808), .B(n_735), .Y(n_849) );
INVx1_ASAP7_75t_SL g850 ( .A(n_796), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_800), .Y(n_851) );
INVxp67_ASAP7_75t_L g852 ( .A(n_804), .Y(n_852) );
XNOR2xp5_ASAP7_75t_L g853 ( .A(n_829), .B(n_747), .Y(n_853) );
XOR2x2_ASAP7_75t_L g854 ( .A(n_829), .B(n_735), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_817), .Y(n_855) );
XOR2x2_ASAP7_75t_L g856 ( .A(n_809), .B(n_728), .Y(n_856) );
INVx2_ASAP7_75t_SL g857 ( .A(n_796), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_834), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_836), .Y(n_859) );
OA22x2_ASAP7_75t_L g860 ( .A1(n_838), .A2(n_804), .B1(n_794), .B2(n_825), .Y(n_860) );
INVxp67_ASAP7_75t_SL g861 ( .A(n_852), .Y(n_861) );
INVxp67_ASAP7_75t_L g862 ( .A(n_832), .Y(n_862) );
INVx2_ASAP7_75t_SL g863 ( .A(n_841), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_851), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_846), .A2(n_811), .B1(n_806), .B2(n_803), .Y(n_865) );
OA22x2_ASAP7_75t_L g866 ( .A1(n_853), .A2(n_794), .B1(n_818), .B2(n_822), .Y(n_866) );
OA22x2_ASAP7_75t_L g867 ( .A1(n_853), .A2(n_818), .B1(n_822), .B2(n_801), .Y(n_867) );
OA22x2_ASAP7_75t_L g868 ( .A1(n_835), .A2(n_822), .B1(n_818), .B2(n_812), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_841), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_855), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_857), .Y(n_871) );
XOR2x2_ASAP7_75t_L g872 ( .A(n_840), .B(n_809), .Y(n_872) );
AND2x4_ASAP7_75t_L g873 ( .A(n_857), .B(n_813), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_861), .Y(n_874) );
INVxp33_ASAP7_75t_SL g875 ( .A(n_867), .Y(n_875) );
XNOR2xp5_ASAP7_75t_L g876 ( .A(n_872), .B(n_840), .Y(n_876) );
XNOR2xp5_ASAP7_75t_L g877 ( .A(n_867), .B(n_837), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_864), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_858), .Y(n_879) );
AOI322xp5_ASAP7_75t_L g880 ( .A1(n_862), .A2(n_843), .A3(n_830), .B1(n_831), .B2(n_842), .C1(n_839), .C2(n_847), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_859), .Y(n_881) );
OAI322xp33_ASAP7_75t_L g882 ( .A1(n_866), .A2(n_846), .A3(n_844), .B1(n_821), .B2(n_842), .C1(n_850), .C2(n_848), .Y(n_882) );
AOI22x1_ASAP7_75t_L g883 ( .A1(n_877), .A2(n_860), .B1(n_866), .B2(n_871), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_874), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_875), .A2(n_860), .B1(n_868), .B2(n_865), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_875), .A2(n_837), .B1(n_832), .B2(n_833), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_878), .Y(n_887) );
A2O1A1Ixp33_ASAP7_75t_L g888 ( .A1(n_886), .A2(n_880), .B(n_865), .C(n_863), .Y(n_888) );
NAND4xp75_ASAP7_75t_L g889 ( .A(n_883), .B(n_877), .C(n_882), .D(n_876), .Y(n_889) );
INVx2_ASAP7_75t_SL g890 ( .A(n_884), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_890), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_888), .B(n_885), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_889), .A2(n_833), .B1(n_868), .B2(n_844), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_893), .A2(n_856), .B1(n_887), .B2(n_854), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_891), .Y(n_895) );
AND4x1_ASAP7_75t_L g896 ( .A(n_895), .B(n_892), .C(n_883), .D(n_881), .Y(n_896) );
AND4x1_ASAP7_75t_L g897 ( .A(n_894), .B(n_879), .C(n_843), .D(n_856), .Y(n_897) );
XNOR2xp5_ASAP7_75t_L g898 ( .A(n_896), .B(n_854), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_897), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_899), .A2(n_873), .B1(n_869), .B2(n_826), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_900), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g902 ( .A1(n_901), .A2(n_898), .B1(n_873), .B2(n_810), .Y(n_902) );
INVxp67_ASAP7_75t_L g903 ( .A(n_902), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_903), .A2(n_870), .B1(n_845), .B2(n_831), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_904), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_905), .A2(n_823), .B1(n_820), .B2(n_849), .C(n_815), .Y(n_906) );
AOI211xp5_ASAP7_75t_L g907 ( .A1(n_906), .A2(n_799), .B(n_814), .C(n_849), .Y(n_907) );
endmodule