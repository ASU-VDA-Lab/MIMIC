module real_aes_6422_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
NOR4xp25_ASAP7_75t_SL g22 ( .A(n_0), .B(n_7), .C(n_9), .D(n_23), .Y(n_22) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_1), .B(n_9), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_2), .Y(n_20) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_3), .B(n_6), .C(n_19), .Y(n_18) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_4), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_5), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_8), .Y(n_21) );
AOI31xp33_ASAP7_75t_R g10 ( .A1(n_11), .A2(n_12), .A3(n_13), .B(n_22), .Y(n_10) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_14), .B(n_16), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_16), .Y(n_24) );
NAND2xp33_ASAP7_75t_SL g16 ( .A(n_17), .B(n_21), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_18), .B(n_20), .Y(n_17) );
NAND2xp33_ASAP7_75t_SL g23 ( .A(n_24), .B(n_25), .Y(n_23) );
endmodule