module fake_jpeg_12602_n_117 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_117);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_117;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_7),
.B(n_0),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_9),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_49),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_25),
.C(n_21),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_49),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_19),
.B1(n_25),
.B2(n_11),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_53),
.B1(n_58),
.B2(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_19),
.B1(n_11),
.B2(n_13),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_13),
.B1(n_21),
.B2(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_29),
.A2(n_2),
.B1(n_15),
.B2(n_43),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_2),
.B(n_36),
.C(n_15),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_35),
.B(n_15),
.C(n_48),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_51),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_65),
.B1(n_59),
.B2(n_70),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_68),
.B1(n_58),
.B2(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_68),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_66),
.C(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_55),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_81),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_74),
.C(n_77),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_54),
.B1(n_69),
.B2(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_93),
.A2(n_76),
.B1(n_82),
.B2(n_79),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_97),
.B1(n_94),
.B2(n_71),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_SL g103 ( 
.A1(n_95),
.A2(n_86),
.A3(n_92),
.B1(n_87),
.B2(n_74),
.C1(n_88),
.C2(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_96),
.C(n_98),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_106),
.A2(n_97),
.B1(n_89),
.B2(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_102),
.C(n_104),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_106),
.B1(n_105),
.B2(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.Y(n_114)
);

AOI321xp33_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_113),
.A3(n_109),
.B1(n_89),
.B2(n_66),
.C(n_57),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_115),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_57),
.Y(n_117)
);


endmodule