module fake_netlist_6_1525_n_2329 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2329);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2329;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_2292;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_89),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_80),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_52),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_226),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_145),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_202),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_111),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_118),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_89),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_162),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_123),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_132),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_148),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_69),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_140),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_102),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_114),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_186),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_116),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_110),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_39),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_176),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_119),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_81),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_52),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_72),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_53),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_85),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_87),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_232),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_101),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_212),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_96),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_135),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_168),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_19),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_4),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_25),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_190),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_20),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_199),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_197),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_153),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_196),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_223),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_28),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_27),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_90),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_171),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_65),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_170),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_82),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_205),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_25),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_38),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_174),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_181),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_136),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_56),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_79),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_178),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_156),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_146),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_194),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_17),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_120),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_231),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_29),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_155),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_195),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_10),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_34),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_1),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_8),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_203),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_185),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_14),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_213),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_97),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_103),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_201),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_46),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_210),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_144),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_177),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_30),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_126),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_40),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_159),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_138),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_109),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_66),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_22),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_53),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_14),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_129),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_106),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_10),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_6),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_49),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_228),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_161),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_16),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_227),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_115),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_11),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_125),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_217),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_61),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_165),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_7),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_92),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_90),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_39),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_23),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_54),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_63),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_36),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_164),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_37),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_63),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_9),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_86),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_204),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_26),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_38),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_28),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_163),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_95),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_160),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_40),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_216),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_57),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_33),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_78),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_184),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_220),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_200),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_219),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_62),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_55),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_51),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_141),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_137),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_4),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_180),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_61),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_51),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_46),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_108),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_211),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_175),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_215),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_173),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_70),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_87),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_167),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_158),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_27),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_7),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_43),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_44),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_76),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_208),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_139),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_6),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_214),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_66),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_59),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_92),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_188),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_166),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_172),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_154),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_37),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_3),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_21),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_131),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_79),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_78),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_30),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_209),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_68),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_122),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_64),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_12),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_151),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_36),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_99),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_206),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_74),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_48),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_187),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_35),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_31),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_23),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_58),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_45),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_59),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_67),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_124),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_43),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_19),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_9),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_182),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_130),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_50),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_26),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_113),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_133),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_41),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_80),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_112),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_95),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_83),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_143),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_443),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_293),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_443),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_235),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_240),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_290),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_363),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_235),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_348),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_255),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_255),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_256),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_242),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_237),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_256),
.Y(n_475)
);

INVxp33_ASAP7_75t_SL g476 ( 
.A(n_290),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_248),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_278),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_258),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_233),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_354),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_354),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_233),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_259),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_363),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_263),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_363),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_265),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_268),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_233),
.B(n_0),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_363),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_353),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_308),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_363),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_266),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_388),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_278),
.B(n_0),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_284),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_R g500 ( 
.A(n_327),
.B(n_98),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_350),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_282),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_288),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_282),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_353),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_283),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_400),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_283),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_416),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_304),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_236),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_292),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_425),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_348),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_294),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_304),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_306),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_310),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_306),
.B(n_1),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_313),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_323),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_323),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_334),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_388),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_353),
.B(n_2),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_314),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_261),
.B(n_2),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_334),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_316),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_377),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_351),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_351),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_449),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_328),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_380),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_335),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_380),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_336),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_388),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_338),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_341),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_342),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_396),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_396),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_388),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_377),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_238),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_244),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_343),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_414),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_349),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_245),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_414),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_415),
.B(n_3),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_427),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_427),
.B(n_5),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_430),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_430),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_236),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_234),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_234),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_377),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_234),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_253),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_388),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_352),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_246),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_253),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_247),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_253),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_276),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_250),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_276),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_276),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_R g578 ( 
.A(n_459),
.B(n_5),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_357),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_377),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_361),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_418),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_364),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_249),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_239),
.B(n_326),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_241),
.B(n_8),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_251),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_460),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_461),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_553),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_575),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_480),
.B(n_432),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_461),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_575),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_483),
.B(n_418),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_545),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_467),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_492),
.B(n_456),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_467),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_575),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_485),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_485),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_487),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_585),
.B(n_418),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_487),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_567),
.Y(n_610)
);

OA21x2_ASAP7_75t_L g611 ( 
.A1(n_491),
.A2(n_301),
.B(n_279),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_505),
.B(n_418),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_490),
.B(n_418),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_567),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_553),
.B(n_456),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_494),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_573),
.B(n_456),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_573),
.B(n_324),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_494),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_496),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_562),
.B(n_563),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_496),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_497),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_497),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_524),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_565),
.B(n_324),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_518),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_539),
.B(n_582),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_469),
.B(n_514),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_463),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_539),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_582),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_464),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_468),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_470),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_463),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_471),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_472),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_418),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_475),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_525),
.B(n_299),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_478),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_502),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_504),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_506),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_508),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_465),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

XOR2x2_ASAP7_75t_L g651 ( 
.A(n_527),
.B(n_243),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_516),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_566),
.B(n_324),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_517),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_570),
.B(n_445),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_521),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_572),
.B(n_445),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_474),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_530),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_522),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_523),
.Y(n_661)
);

OA21x2_ASAP7_75t_L g662 ( 
.A1(n_528),
.A2(n_301),
.B(n_279),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_574),
.B(n_360),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

BUFx8_ASAP7_75t_L g665 ( 
.A(n_576),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_532),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_535),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_544),
.B(n_340),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_500),
.B(n_445),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_550),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_554),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_556),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_557),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_474),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_559),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_560),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_577),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_511),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_561),
.B(n_360),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_498),
.B(n_445),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_462),
.B(n_445),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_519),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_555),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_662),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_685),
.A2(n_476),
.B1(n_333),
.B2(n_358),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_662),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_593),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_591),
.B(n_477),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_662),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_659),
.B(n_546),
.Y(n_693)
);

INVxp33_ASAP7_75t_L g694 ( 
.A(n_651),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_594),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_593),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_643),
.B(n_241),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_619),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_593),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_686),
.B(n_241),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_684),
.B(n_595),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_662),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_662),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_684),
.B(n_547),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_684),
.A2(n_476),
.B1(n_481),
.B2(n_466),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_591),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_686),
.B(n_393),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_631),
.A2(n_580),
.B1(n_564),
.B2(n_359),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_684),
.B(n_548),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_595),
.B(n_482),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_594),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_662),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_643),
.B(n_393),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_611),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_611),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_594),
.Y(n_716)
);

CKINVDCx6p67_ASAP7_75t_R g717 ( 
.A(n_659),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_611),
.Y(n_718)
);

INVxp33_ASAP7_75t_L g719 ( 
.A(n_651),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_598),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_685),
.B(n_552),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_593),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_591),
.B(n_477),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_623),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_594),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_608),
.A2(n_402),
.B1(n_403),
.B2(n_289),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_594),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_594),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_594),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_599),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_659),
.B(n_479),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_611),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_686),
.B(n_479),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_686),
.B(n_407),
.C(n_393),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_686),
.B(n_407),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_686),
.B(n_486),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_588),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_630),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_588),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_599),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_630),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_619),
.B(n_486),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_686),
.B(n_488),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_619),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_630),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_623),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_629),
.B(n_569),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_686),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_599),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_659),
.B(n_488),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_598),
.B(n_407),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_630),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_608),
.B(n_495),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_669),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_595),
.B(n_436),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_630),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_659),
.B(n_495),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_594),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_601),
.B(n_499),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_669),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_669),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_601),
.B(n_499),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_682),
.B(n_453),
.C(n_436),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_617),
.Y(n_764)
);

INVx6_ASAP7_75t_L g765 ( 
.A(n_665),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_616),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_617),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_682),
.A2(n_445),
.B1(n_301),
.B2(n_307),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_617),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_667),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_617),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_629),
.B(n_571),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_L g773 ( 
.A(n_680),
.B(n_360),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_667),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_667),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_601),
.B(n_503),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_641),
.A2(n_307),
.B1(n_355),
.B2(n_279),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_590),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_612),
.B(n_503),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_659),
.B(n_512),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_640),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_649),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_659),
.B(n_512),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_641),
.A2(n_307),
.B1(n_356),
.B2(n_355),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_683),
.B(n_584),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_640),
.Y(n_786)
);

BUFx10_ASAP7_75t_L g787 ( 
.A(n_683),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_613),
.B(n_453),
.C(n_436),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_625),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_610),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_667),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_613),
.A2(n_612),
.B1(n_670),
.B2(n_671),
.Y(n_792)
);

INVx4_ASAP7_75t_SL g793 ( 
.A(n_610),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_625),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_667),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_590),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_610),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_616),
.B(n_587),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_589),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_640),
.Y(n_800)
);

AND2x6_ASAP7_75t_L g801 ( 
.A(n_616),
.B(n_453),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_610),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_589),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_625),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_625),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_627),
.Y(n_806)
);

BUFx4f_ASAP7_75t_L g807 ( 
.A(n_640),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_592),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_610),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_627),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_618),
.B(n_515),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_596),
.Y(n_812)
);

XOR2x2_ASAP7_75t_SL g813 ( 
.A(n_651),
.B(n_527),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_618),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_618),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_627),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_649),
.Y(n_817)
);

AO21x2_ASAP7_75t_L g818 ( 
.A1(n_671),
.A2(n_371),
.B(n_340),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_596),
.B(n_515),
.Y(n_819)
);

HAxp5_ASAP7_75t_SL g820 ( 
.A(n_680),
.B(n_267),
.CON(n_820),
.SN(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_681),
.Y(n_821)
);

AND2x6_ASAP7_75t_L g822 ( 
.A(n_670),
.B(n_250),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_600),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_600),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_627),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_634),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_602),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_588),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_634),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_670),
.A2(n_355),
.B1(n_398),
.B2(n_356),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_634),
.Y(n_831)
);

AND3x2_ASAP7_75t_L g832 ( 
.A(n_631),
.B(n_371),
.C(n_356),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_602),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_592),
.Y(n_834)
);

AND2x6_ASAP7_75t_L g835 ( 
.A(n_670),
.B(n_250),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_605),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_622),
.B(n_520),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_605),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_638),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_606),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_610),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_658),
.B(n_520),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_606),
.B(n_526),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_623),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_622),
.B(n_628),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_720),
.B(n_640),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_817),
.Y(n_847)
);

AO221x1_ASAP7_75t_L g848 ( 
.A1(n_778),
.A2(n_658),
.B1(n_676),
.B2(n_638),
.C(n_250),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_730),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_744),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_742),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_701),
.B(n_733),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_821),
.A2(n_635),
.B(n_637),
.C(n_636),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_744),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_738),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_762),
.B(n_658),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_748),
.B(n_676),
.Y(n_857)
);

INVx5_ASAP7_75t_L g858 ( 
.A(n_707),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_701),
.B(n_640),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_753),
.B(n_676),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_748),
.B(n_250),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_748),
.B(n_250),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_742),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_821),
.A2(n_670),
.B(n_681),
.C(n_635),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_738),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_741),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_704),
.A2(n_632),
.B1(n_638),
.B2(n_484),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_740),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_762),
.B(n_681),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_736),
.B(n_640),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_817),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_779),
.B(n_526),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_743),
.A2(n_489),
.B1(n_493),
.B2(n_473),
.Y(n_873)
);

XOR2xp5_ASAP7_75t_L g874 ( 
.A(n_782),
.B(n_501),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_706),
.B(n_622),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_698),
.B(n_628),
.Y(n_876)
);

NOR2x1p5_ASAP7_75t_L g877 ( 
.A(n_759),
.B(n_529),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_740),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_748),
.B(n_665),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_749),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_749),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_700),
.B(n_665),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_741),
.Y(n_883)
);

BUFx6f_ASAP7_75t_SL g884 ( 
.A(n_697),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_700),
.B(n_665),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_700),
.B(n_665),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_706),
.B(n_640),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_766),
.B(n_644),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_776),
.B(n_529),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_709),
.B(n_534),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_766),
.A2(n_632),
.B1(n_509),
.B2(n_513),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_745),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_L g893 ( 
.A(n_755),
.B(n_269),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_787),
.B(n_269),
.Y(n_894)
);

OAI22xp33_ASAP7_75t_L g895 ( 
.A1(n_697),
.A2(n_413),
.B1(n_434),
.B2(n_398),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_787),
.B(n_269),
.Y(n_896)
);

CKINVDCx11_ASAP7_75t_R g897 ( 
.A(n_828),
.Y(n_897)
);

INVx8_ASAP7_75t_L g898 ( 
.A(n_755),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_745),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_710),
.B(n_534),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_814),
.B(n_815),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_737),
.B(n_628),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_721),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_814),
.A2(n_533),
.B1(n_507),
.B2(n_536),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_815),
.B(n_644),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_698),
.B(n_644),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_752),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_756),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_687),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_754),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_752),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_787),
.B(n_269),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_811),
.B(n_536),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_787),
.B(n_269),
.Y(n_914)
);

NOR2xp67_ASAP7_75t_L g915 ( 
.A(n_747),
.B(n_538),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_845),
.B(n_653),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_792),
.B(n_644),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_756),
.B(n_269),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_772),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_785),
.B(n_687),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_754),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_845),
.B(n_644),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_689),
.B(n_692),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_799),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_764),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_737),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_692),
.B(n_644),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_760),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_702),
.B(n_269),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_799),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_702),
.B(n_644),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_819),
.B(n_538),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_760),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_703),
.B(n_269),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_703),
.B(n_269),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_761),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_739),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_803),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_712),
.B(n_648),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_712),
.A2(n_637),
.B(n_642),
.C(n_636),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_770),
.B(n_648),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_739),
.Y(n_942)
);

BUFx6f_ASAP7_75t_SL g943 ( 
.A(n_697),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_764),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_714),
.B(n_648),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_697),
.A2(n_454),
.B1(n_458),
.B2(n_419),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_714),
.B(n_648),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_808),
.A2(n_657),
.B(n_655),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_715),
.B(n_648),
.Y(n_949)
);

BUFx8_ASAP7_75t_L g950 ( 
.A(n_839),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_715),
.B(n_648),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_812),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_770),
.B(n_648),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_812),
.Y(n_954)
);

INVxp67_ASAP7_75t_SL g955 ( 
.A(n_718),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_823),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_823),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_755),
.A2(n_541),
.B1(n_542),
.B2(n_540),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_774),
.B(n_648),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_843),
.B(n_541),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_718),
.B(n_652),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_763),
.A2(n_398),
.B1(n_434),
.B2(n_413),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_767),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_774),
.B(n_652),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_767),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_824),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_755),
.A2(n_549),
.B1(n_551),
.B2(n_542),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_839),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_SL g969 ( 
.A(n_798),
.B(n_549),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_824),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_773),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_827),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_691),
.B(n_551),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_827),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_732),
.B(n_652),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_769),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_761),
.B(n_642),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_833),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_763),
.B(n_568),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_833),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_769),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_697),
.A2(n_389),
.B1(n_387),
.B2(n_568),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_771),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_836),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_732),
.B(n_652),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_723),
.B(n_579),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_775),
.A2(n_791),
.B(n_795),
.C(n_710),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_796),
.B(n_837),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_705),
.B(n_726),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_836),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_837),
.B(n_579),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_L g992 ( 
.A1(n_726),
.A2(n_262),
.B1(n_264),
.B2(n_366),
.C(n_319),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_773),
.B(n_581),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_775),
.B(n_654),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_832),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_791),
.B(n_654),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_838),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_755),
.A2(n_581),
.B1(n_583),
.B2(n_578),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_838),
.Y(n_999)
);

OR2x6_ASAP7_75t_L g1000 ( 
.A(n_842),
.B(n_653),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_795),
.B(n_690),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_L g1002 ( 
.A(n_693),
.B(n_708),
.C(n_731),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_840),
.B(n_654),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_713),
.A2(n_583),
.B1(n_254),
.B2(n_257),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_688),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_789),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_713),
.B(n_653),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_921),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_852),
.A2(n_713),
.B1(n_765),
.B2(n_751),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_L g1010 ( 
.A(n_898),
.B(n_801),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_920),
.A2(n_940),
.B(n_895),
.C(n_987),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_860),
.B(n_713),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_908),
.Y(n_1013)
);

AOI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_890),
.A2(n_719),
.B(n_694),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_846),
.A2(n_807),
.B(n_834),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_917),
.A2(n_807),
.B(n_800),
.Y(n_1016)
);

NOR2x1p5_ASAP7_75t_L g1017 ( 
.A(n_989),
.B(n_820),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_870),
.A2(n_807),
.B(n_800),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_858),
.B(n_690),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_897),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_856),
.B(n_688),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_859),
.A2(n_800),
.B(n_724),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_890),
.B(n_757),
.C(n_750),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_860),
.B(n_713),
.Y(n_1024)
);

OAI321xp33_ASAP7_75t_L g1025 ( 
.A1(n_992),
.A2(n_982),
.A3(n_903),
.B1(n_1005),
.B2(n_895),
.C(n_919),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_923),
.A2(n_947),
.B(n_945),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_955),
.B(n_840),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_894),
.A2(n_699),
.B(n_696),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_955),
.B(n_751),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_949),
.A2(n_961),
.B(n_951),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_855),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_921),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_909),
.B(n_751),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_865),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_909),
.B(n_751),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_872),
.B(n_751),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_920),
.A2(n_783),
.B(n_780),
.C(n_647),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_929),
.A2(n_734),
.B(n_707),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_857),
.A2(n_864),
.B(n_934),
.C(n_929),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_894),
.A2(n_699),
.B(n_696),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1002),
.A2(n_801),
.B1(n_735),
.B2(n_707),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_872),
.B(n_801),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_850),
.B(n_801),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_900),
.B(n_663),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_850),
.B(n_801),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_858),
.B(n_722),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_962),
.A2(n_768),
.B1(n_784),
.B2(n_777),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_901),
.B(n_801),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_924),
.B(n_801),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_930),
.B(n_722),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_938),
.B(n_818),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_975),
.A2(n_985),
.B(n_927),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_896),
.A2(n_794),
.B(n_789),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_952),
.B(n_818),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_934),
.A2(n_734),
.B(n_707),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_889),
.B(n_302),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_935),
.A2(n_735),
.B(n_707),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_931),
.A2(n_844),
.B(n_746),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_866),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_926),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_954),
.B(n_707),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_956),
.B(n_707),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_939),
.A2(n_922),
.B(n_887),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_935),
.A2(n_735),
.B(n_788),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_869),
.A2(n_788),
.B(n_830),
.C(n_820),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_921),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_883),
.A2(n_765),
.B1(n_717),
.B2(n_725),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_858),
.B(n_790),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_957),
.B(n_966),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_892),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_847),
.B(n_765),
.Y(n_1071)
);

AOI33xp33_ASAP7_75t_L g1072 ( 
.A1(n_946),
.A2(n_267),
.A3(n_273),
.B1(n_275),
.B2(n_277),
.B3(n_440),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_899),
.A2(n_663),
.B(n_434),
.C(n_450),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_970),
.B(n_735),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_907),
.Y(n_1075)
);

AOI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_889),
.A2(n_370),
.B(n_365),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_991),
.B(n_663),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_950),
.Y(n_1078)
);

AOI33xp33_ASAP7_75t_L g1079 ( 
.A1(n_851),
.A2(n_368),
.A3(n_273),
.B1(n_275),
.B2(n_277),
.B3(n_297),
.Y(n_1079)
);

OR2x2_ASAP7_75t_SL g1080 ( 
.A(n_969),
.B(n_813),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_911),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_972),
.B(n_735),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_974),
.B(n_735),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_916),
.B(n_679),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_L g1085 ( 
.A(n_904),
.B(n_679),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_916),
.B(n_647),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_978),
.B(n_735),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_980),
.B(n_716),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_857),
.A2(n_765),
.B1(n_717),
.B2(n_725),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_984),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_913),
.B(n_863),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_990),
.B(n_716),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_997),
.B(n_716),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1002),
.A2(n_450),
.B(n_413),
.C(n_297),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1007),
.A2(n_728),
.B1(n_729),
.B2(n_725),
.Y(n_1095)
);

NOR2x2_ASAP7_75t_L g1096 ( 
.A(n_988),
.B(n_813),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_896),
.A2(n_729),
.B(n_728),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_999),
.B(n_728),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_888),
.A2(n_711),
.B(n_695),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_858),
.B(n_695),
.Y(n_1100)
);

NOR2x1p5_ASAP7_75t_L g1101 ( 
.A(n_968),
.B(n_369),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_876),
.B(n_650),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_876),
.B(n_650),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_932),
.B(n_729),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_905),
.A2(n_906),
.B(n_898),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_932),
.B(n_758),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_SL g1107 ( 
.A(n_871),
.B(n_299),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_921),
.B(n_928),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_928),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_854),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_898),
.A2(n_711),
.B(n_695),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_861),
.A2(n_711),
.B(n_695),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_913),
.B(n_656),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_873),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_861),
.A2(n_711),
.B(n_695),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_862),
.A2(n_727),
.B(n_781),
.Y(n_1116)
);

NOR3xp33_ASAP7_75t_L g1117 ( 
.A(n_960),
.B(n_660),
.C(n_656),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_960),
.A2(n_986),
.B(n_973),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_L g1119 ( 
.A1(n_912),
.A2(n_804),
.B(n_794),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_973),
.B(n_758),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1001),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_862),
.A2(n_948),
.B(n_1001),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_849),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_986),
.B(n_758),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_995),
.A2(n_664),
.B(n_666),
.C(n_660),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_928),
.B(n_727),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_902),
.B(n_664),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_912),
.A2(n_727),
.B(n_781),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_914),
.A2(n_727),
.B(n_781),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_902),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_875),
.B(n_790),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_928),
.B(n_727),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_937),
.B(n_666),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_875),
.B(n_797),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_936),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_971),
.B(n_668),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_853),
.A2(n_673),
.B(n_674),
.C(n_668),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_914),
.A2(n_786),
.B(n_781),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_918),
.A2(n_786),
.B(n_781),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_936),
.B(n_797),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_979),
.B(n_797),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_918),
.A2(n_786),
.B(n_802),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_868),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1007),
.A2(n_809),
.B1(n_841),
.B2(n_802),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1003),
.A2(n_786),
.B(n_802),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_878),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_942),
.B(n_673),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_936),
.B(n_809),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_867),
.B(n_674),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_893),
.A2(n_786),
.B(n_809),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_882),
.A2(n_678),
.B(n_655),
.C(n_657),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_941),
.A2(n_959),
.B(n_953),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_880),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_882),
.A2(n_678),
.B(n_639),
.C(n_646),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_885),
.A2(n_841),
.B(n_592),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_936),
.B(n_841),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_902),
.B(n_372),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_962),
.A2(n_998),
.B(n_885),
.C(n_886),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_886),
.A2(n_953),
.B(n_941),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_910),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_910),
.B(n_804),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_933),
.B(n_805),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_L g1163 ( 
.A(n_915),
.B(n_385),
.C(n_378),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1004),
.A2(n_639),
.B(n_646),
.C(n_645),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_958),
.B(n_805),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_848),
.A2(n_450),
.B1(n_374),
.B2(n_383),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_933),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_988),
.B(n_390),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_959),
.A2(n_592),
.B(n_806),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_993),
.B(n_806),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_964),
.A2(n_592),
.B(n_810),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_964),
.A2(n_816),
.B(n_810),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_977),
.B(n_881),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_994),
.A2(n_825),
.B(n_816),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_925),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_977),
.B(n_825),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_944),
.Y(n_1177)
);

AOI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1000),
.A2(n_406),
.B(n_399),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_988),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1007),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_994),
.A2(n_829),
.B(n_826),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1006),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_996),
.A2(n_829),
.B(n_826),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_963),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_965),
.B(n_976),
.Y(n_1185)
);

CKINVDCx10_ASAP7_75t_R g1186 ( 
.A(n_874),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_967),
.B(n_831),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_996),
.A2(n_831),
.B(n_603),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_981),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_891),
.B(n_793),
.Y(n_1190)
);

BUFx12f_ASAP7_75t_L g1191 ( 
.A(n_1078),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_1020),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1180),
.B(n_1000),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1060),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1031),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1113),
.B(n_877),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1113),
.B(n_1000),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1026),
.A2(n_879),
.B(n_983),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1118),
.A2(n_639),
.B(n_646),
.C(n_645),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1056),
.B(n_645),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_1066),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1056),
.B(n_645),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1030),
.A2(n_603),
.B(n_597),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1052),
.A2(n_603),
.B(n_597),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1091),
.B(n_950),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1091),
.B(n_646),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1066),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1179),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1096),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1025),
.B(n_252),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1044),
.B(n_661),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1063),
.A2(n_1105),
.B(n_1042),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_R g1213 ( 
.A(n_1114),
.B(n_884),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1066),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1066),
.Y(n_1215)
);

NOR2x1_ASAP7_75t_L g1216 ( 
.A(n_1135),
.B(n_369),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1031),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1076),
.A2(n_315),
.B(n_337),
.C(n_330),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1017),
.A2(n_1024),
.B1(n_1012),
.B2(n_1021),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_1107),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1130),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1014),
.B(n_884),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1122),
.A2(n_1039),
.B(n_1048),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1158),
.A2(n_374),
.B(n_383),
.C(n_369),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1010),
.A2(n_603),
.B(n_597),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1158),
.A2(n_604),
.B(n_597),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1077),
.B(n_661),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1180),
.Y(n_1228)
);

NOR2xp67_ASAP7_75t_L g1229 ( 
.A(n_1110),
.B(n_260),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_1180),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1094),
.A2(n_315),
.B(n_337),
.C(n_330),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1127),
.B(n_661),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_R g1233 ( 
.A(n_1071),
.B(n_943),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1086),
.B(n_661),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1070),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1070),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1016),
.A2(n_604),
.B(n_675),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1160),
.B(n_607),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1180),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1034),
.B(n_675),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1036),
.A2(n_392),
.B(n_437),
.C(n_405),
.Y(n_1241)
);

INVxp33_ASAP7_75t_L g1242 ( 
.A(n_1168),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1059),
.B(n_675),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1186),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1102),
.B(n_270),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1081),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1081),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1104),
.A2(n_604),
.B(n_675),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1106),
.A2(n_604),
.B(n_615),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1015),
.A2(n_615),
.B(n_634),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1135),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1018),
.A2(n_615),
.B(n_654),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1080),
.B(n_411),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1120),
.A2(n_615),
.B(n_654),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1053),
.A2(n_609),
.B(n_607),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1102),
.B(n_271),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1103),
.B(n_272),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1069),
.B(n_609),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1029),
.A2(n_943),
.B1(n_367),
.B2(n_362),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1130),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1103),
.B(n_274),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1033),
.A2(n_295),
.B1(n_285),
.B2(n_281),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1101),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_SL g1264 ( 
.A1(n_1023),
.A2(n_614),
.B(n_620),
.C(n_633),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1167),
.B(n_1075),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1035),
.A2(n_298),
.B1(n_286),
.B2(n_287),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1094),
.A2(n_620),
.B(n_614),
.Y(n_1267)
);

AND2x6_ASAP7_75t_L g1268 ( 
.A(n_1041),
.B(n_346),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1168),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1090),
.B(n_621),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1027),
.A2(n_280),
.B1(n_291),
.B2(n_300),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1065),
.A2(n_440),
.B(n_424),
.C(n_412),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1149),
.B(n_420),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1167),
.B(n_303),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1084),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1124),
.A2(n_672),
.B(n_654),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1008),
.B(n_374),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1157),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1051),
.A2(n_633),
.B(n_624),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1136),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1011),
.A2(n_677),
.B(n_672),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_SL g1282 ( 
.A(n_1163),
.B(n_426),
.C(n_423),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1149),
.B(n_429),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1170),
.A2(n_677),
.B(n_672),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1013),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1175),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1117),
.A2(n_835),
.B1(n_822),
.B2(n_299),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1160),
.B(n_305),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1136),
.B(n_309),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1157),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1065),
.A2(n_437),
.B(n_405),
.C(n_392),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1133),
.B(n_624),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1178),
.B(n_431),
.Y(n_1293)
);

BUFx4f_ASAP7_75t_L g1294 ( 
.A(n_1032),
.Y(n_1294)
);

NOR3xp33_ASAP7_75t_L g1295 ( 
.A(n_1133),
.B(n_441),
.C(n_438),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1147),
.B(n_442),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1147),
.B(n_672),
.Y(n_1297)
);

AOI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1054),
.A2(n_368),
.B(n_346),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1028),
.A2(n_384),
.B(n_376),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1047),
.A2(n_397),
.B1(n_311),
.B2(n_317),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1032),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1190),
.A2(n_384),
.B(n_435),
.C(n_376),
.Y(n_1302)
);

INVx5_ASAP7_75t_L g1303 ( 
.A(n_1109),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1037),
.A2(n_1159),
.B(n_1085),
.C(n_1121),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1165),
.A2(n_677),
.B(n_672),
.Y(n_1305)
);

BUFx8_ASAP7_75t_L g1306 ( 
.A(n_1123),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1050),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1109),
.B(n_672),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1177),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_SL g1310 ( 
.A(n_1190),
.B(n_447),
.C(n_446),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1072),
.B(n_439),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1008),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1153),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1072),
.B(n_677),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1165),
.A2(n_677),
.B(n_610),
.Y(n_1315)
);

OAI21xp33_ASAP7_75t_L g1316 ( 
.A1(n_1079),
.A2(n_455),
.B(n_451),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1184),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1143),
.B(n_822),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_L g1319 ( 
.A(n_1125),
.B(n_457),
.C(n_321),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1189),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1108),
.B(n_391),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1146),
.B(n_320),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1049),
.A2(n_437),
.B(n_383),
.C(n_405),
.Y(n_1323)
);

NAND2xp33_ASAP7_75t_L g1324 ( 
.A(n_1182),
.B(n_822),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1043),
.A2(n_339),
.B1(n_322),
.B2(n_325),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1182),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1182),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1182),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1173),
.B(n_329),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1079),
.B(n_822),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1137),
.B(n_822),
.Y(n_1331)
);

INVx5_ASAP7_75t_L g1332 ( 
.A(n_1068),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1187),
.A2(n_610),
.B(n_623),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1185),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1009),
.B(n_331),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1045),
.B(n_332),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1187),
.A2(n_623),
.B(n_626),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1088),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1108),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1161),
.B(n_344),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1151),
.A2(n_392),
.B(n_391),
.C(n_404),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1064),
.A2(n_422),
.B(n_404),
.C(n_409),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1152),
.Y(n_1343)
);

NOR3xp33_ASAP7_75t_SL g1344 ( 
.A(n_1073),
.B(n_408),
.C(n_448),
.Y(n_1344)
);

O2A1O1Ixp5_ASAP7_75t_L g1345 ( 
.A1(n_1067),
.A2(n_296),
.B(n_412),
.C(n_428),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1166),
.B(n_822),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1148),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1166),
.B(n_822),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1022),
.A2(n_623),
.B(n_626),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1176),
.B(n_345),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1092),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1304),
.A2(n_1089),
.B(n_1111),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1194),
.Y(n_1353)
);

BUFx10_ASAP7_75t_L g1354 ( 
.A(n_1205),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1219),
.B(n_1307),
.Y(n_1355)
);

AND2x6_ASAP7_75t_L g1356 ( 
.A(n_1228),
.B(n_1131),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1224),
.A2(n_1073),
.A3(n_1144),
.B(n_1095),
.Y(n_1357)
);

AO21x1_ASAP7_75t_L g1358 ( 
.A1(n_1335),
.A2(n_1154),
.B(n_1164),
.Y(n_1358)
);

NOR2xp67_ASAP7_75t_L g1359 ( 
.A(n_1196),
.B(n_1141),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1195),
.Y(n_1360)
);

AOI221x1_ASAP7_75t_L g1361 ( 
.A1(n_1273),
.A2(n_1155),
.B1(n_1038),
.B2(n_1055),
.C(n_1057),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1283),
.B(n_1162),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1279),
.A2(n_1040),
.B(n_1119),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1208),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1255),
.A2(n_1099),
.B(n_1145),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1252),
.A2(n_1129),
.B(n_1128),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1252),
.A2(n_1138),
.B(n_1058),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1197),
.A2(n_1126),
.B1(n_1132),
.B2(n_1098),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1296),
.A2(n_1342),
.B1(n_1292),
.B2(n_1291),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1293),
.A2(n_1061),
.B(n_1083),
.C(n_1062),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1244),
.Y(n_1371)
);

AOI221x1_ASAP7_75t_L g1372 ( 
.A1(n_1341),
.A2(n_1097),
.B1(n_1134),
.B2(n_1087),
.C(n_1082),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1281),
.A2(n_1174),
.B(n_1172),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1281),
.A2(n_1183),
.B(n_1181),
.Y(n_1374)
);

BUFx10_ASAP7_75t_L g1375 ( 
.A(n_1222),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1236),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1193),
.B(n_1156),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_1280),
.B(n_1074),
.Y(n_1378)
);

BUFx12f_ASAP7_75t_L g1379 ( 
.A(n_1191),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1272),
.A2(n_409),
.B(n_422),
.C(n_424),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1218),
.A2(n_428),
.B(n_435),
.C(n_296),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1217),
.Y(n_1382)
);

NAND2x1_ASAP7_75t_L g1383 ( 
.A(n_1201),
.B(n_1093),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1235),
.A2(n_1132),
.B1(n_1126),
.B2(n_1140),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1295),
.A2(n_1140),
.B(n_1046),
.C(n_1019),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1349),
.A2(n_1237),
.B(n_1204),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1269),
.B(n_1068),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1221),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1334),
.B(n_1019),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1226),
.A2(n_1188),
.B(n_1150),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1198),
.A2(n_1116),
.A3(n_1115),
.B(n_1112),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1220),
.A2(n_410),
.B1(n_347),
.B2(n_386),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1310),
.A2(n_1142),
.B(n_1139),
.C(n_1171),
.Y(n_1393)
);

BUFx2_ASAP7_75t_SL g1394 ( 
.A(n_1230),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1198),
.A2(n_1046),
.B(n_1100),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1206),
.B(n_1100),
.Y(n_1396)
);

AOI221x1_ASAP7_75t_L g1397 ( 
.A1(n_1241),
.A2(n_1169),
.B1(n_626),
.B2(n_623),
.C(n_394),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1286),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1246),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1226),
.A2(n_835),
.A3(n_793),
.B(n_417),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1305),
.A2(n_395),
.B(n_375),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1338),
.B(n_835),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1247),
.Y(n_1403)
);

AOI221xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1210),
.A2(n_439),
.B1(n_373),
.B2(n_417),
.C(n_394),
.Y(n_1404)
);

AO31x2_ASAP7_75t_L g1405 ( 
.A1(n_1323),
.A2(n_835),
.A3(n_793),
.B(n_417),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1275),
.Y(n_1406)
);

BUFx4f_ASAP7_75t_L g1407 ( 
.A(n_1251),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1336),
.A2(n_421),
.B(n_381),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1297),
.A2(n_433),
.B(n_401),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1242),
.B(n_299),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1260),
.Y(n_1411)
);

AO32x2_ASAP7_75t_L g1412 ( 
.A1(n_1259),
.A2(n_439),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1351),
.B(n_835),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1313),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1200),
.B(n_379),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1202),
.A2(n_452),
.B(n_444),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1258),
.B(n_382),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1209),
.B(n_439),
.Y(n_1418)
);

AOI22x1_ASAP7_75t_L g1419 ( 
.A1(n_1339),
.A2(n_626),
.B1(n_417),
.B2(n_394),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1309),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1306),
.Y(n_1421)
);

AOI221xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1302),
.A2(n_1316),
.B1(n_1231),
.B2(n_1311),
.C(n_1314),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1211),
.A2(n_626),
.B(n_179),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1290),
.B(n_312),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1193),
.B(n_626),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_SL g1426 ( 
.A(n_1278),
.B(n_394),
.C(n_373),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1227),
.B(n_626),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1199),
.A2(n_312),
.B(n_373),
.Y(n_1428)
);

BUFx8_ASAP7_75t_L g1429 ( 
.A(n_1263),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1192),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1288),
.A2(n_626),
.B(n_169),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1193),
.B(n_100),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1251),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1350),
.A2(n_1324),
.B(n_1340),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1345),
.A2(n_373),
.B(n_318),
.C(n_312),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_SL g1436 ( 
.A1(n_1330),
.A2(n_318),
.B(n_312),
.C(n_230),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1248),
.A2(n_318),
.B(n_229),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1322),
.A2(n_318),
.B(n_13),
.C(n_15),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_1251),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1317),
.Y(n_1440)
);

AO31x2_ASAP7_75t_L g1441 ( 
.A1(n_1343),
.A2(n_11),
.A3(n_16),
.B(n_18),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1203),
.A2(n_222),
.B(n_221),
.Y(n_1442)
);

AO31x2_ASAP7_75t_L g1443 ( 
.A1(n_1305),
.A2(n_22),
.A3(n_24),
.B(n_29),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1276),
.A2(n_24),
.A3(n_31),
.B(n_32),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_SL g1445 ( 
.A1(n_1264),
.A2(n_207),
.B(n_198),
.C(n_193),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1319),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1214),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1232),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1329),
.A2(n_192),
.B(n_191),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1204),
.A2(n_152),
.B(n_150),
.Y(n_1450)
);

AOI221x1_ASAP7_75t_L g1451 ( 
.A1(n_1276),
.A2(n_1248),
.B1(n_1254),
.B2(n_1315),
.C(n_1284),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1250),
.A2(n_149),
.B(n_147),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1232),
.B(n_35),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1344),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1213),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1285),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1320),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_SL g1458 ( 
.A(n_1230),
.B(n_47),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1331),
.A2(n_142),
.B(n_134),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1240),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1243),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1284),
.A2(n_128),
.B(n_127),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_SL g1463 ( 
.A1(n_1346),
.A2(n_121),
.B(n_117),
.C(n_107),
.Y(n_1463)
);

NOR2xp67_ASAP7_75t_L g1464 ( 
.A(n_1282),
.B(n_105),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1234),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1250),
.A2(n_104),
.B(n_50),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1253),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1234),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1321),
.B(n_57),
.Y(n_1469)
);

AO31x2_ASAP7_75t_L g1470 ( 
.A1(n_1315),
.A2(n_58),
.A3(n_60),
.B(n_62),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1333),
.A2(n_60),
.B(n_64),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_SL g1472 ( 
.A1(n_1298),
.A2(n_1299),
.B(n_1326),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1233),
.B(n_65),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1214),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1289),
.B(n_67),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1265),
.A2(n_68),
.B(n_70),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_SL g1477 ( 
.A1(n_1348),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1300),
.B(n_71),
.C(n_74),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1254),
.A2(n_75),
.B(n_76),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1216),
.B(n_75),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1333),
.A2(n_77),
.B(n_81),
.Y(n_1481)
);

AOI211x1_ASAP7_75t_L g1482 ( 
.A1(n_1245),
.A2(n_77),
.B(n_82),
.C(n_83),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1337),
.A2(n_84),
.B(n_85),
.Y(n_1483)
);

AOI221x1_ASAP7_75t_L g1484 ( 
.A1(n_1249),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.C(n_91),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1306),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1268),
.B(n_88),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1337),
.A2(n_91),
.B(n_93),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1225),
.A2(n_94),
.B(n_1308),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1270),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1271),
.B(n_1262),
.C(n_1266),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_SL g1491 ( 
.A1(n_1274),
.A2(n_1318),
.B(n_1261),
.C(n_1257),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1321),
.B(n_1277),
.Y(n_1492)
);

AOI221x1_ASAP7_75t_L g1493 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1327),
.B2(n_1215),
.C(n_1207),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1214),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1267),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1228),
.Y(n_1496)
);

A2O1A1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1229),
.A2(n_1347),
.B(n_1256),
.C(n_1287),
.Y(n_1497)
);

AO31x2_ASAP7_75t_L g1498 ( 
.A1(n_1267),
.A2(n_1201),
.A3(n_1268),
.B(n_1238),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1268),
.A2(n_1277),
.B1(n_1228),
.B2(n_1301),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1332),
.A2(n_1294),
.B(n_1303),
.Y(n_1500)
);

BUFx8_ASAP7_75t_L g1501 ( 
.A(n_1268),
.Y(n_1501)
);

NOR2x1_ASAP7_75t_SL g1502 ( 
.A(n_1230),
.B(n_1239),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1303),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1230),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1268),
.B(n_1312),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1294),
.A2(n_1277),
.B(n_1215),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1332),
.A2(n_1303),
.B(n_1239),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1239),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1239),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1332),
.A2(n_1212),
.B(n_1223),
.Y(n_1510)
);

AO32x2_ASAP7_75t_L g1511 ( 
.A1(n_1303),
.A2(n_1259),
.A3(n_1300),
.B1(n_1009),
.B2(n_1144),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1332),
.A2(n_1118),
.B(n_1056),
.C(n_903),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1212),
.A2(n_1223),
.B(n_852),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1273),
.A2(n_1283),
.B1(n_1017),
.B2(n_1056),
.Y(n_1514)
);

AOI221x1_ASAP7_75t_L g1515 ( 
.A1(n_1273),
.A2(n_1118),
.B1(n_1283),
.B2(n_890),
.C(n_1212),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1219),
.B(n_1118),
.Y(n_1516)
);

NAND2x1_ASAP7_75t_L g1517 ( 
.A(n_1201),
.B(n_1008),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1251),
.Y(n_1518)
);

NOR4xp25_ASAP7_75t_L g1519 ( 
.A(n_1272),
.B(n_1118),
.C(n_1291),
.D(n_1218),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1217),
.Y(n_1520)
);

BUFx2_ASAP7_75t_R g1521 ( 
.A(n_1371),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1514),
.A2(n_1478),
.B1(n_1516),
.B2(n_1467),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1411),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1407),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1514),
.A2(n_1478),
.B1(n_1362),
.B2(n_1369),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1453),
.B(n_1448),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1456),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1369),
.A2(n_1487),
.B1(n_1475),
.B2(n_1457),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.B(n_1480),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1407),
.Y(n_1530)
);

BUFx10_ASAP7_75t_L g1531 ( 
.A(n_1455),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1487),
.A2(n_1457),
.B1(n_1426),
.B2(n_1355),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1355),
.A2(n_1489),
.B1(n_1458),
.B2(n_1490),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1424),
.A2(n_1497),
.B1(n_1388),
.B2(n_1359),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1382),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1406),
.Y(n_1537)
);

INVx6_ASAP7_75t_L g1538 ( 
.A(n_1504),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1430),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1353),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1360),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1458),
.A2(n_1501),
.B1(n_1490),
.B2(n_1419),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1376),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1486),
.A2(n_1437),
.B1(n_1473),
.B2(n_1469),
.Y(n_1544)
);

INVx8_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1417),
.B(n_1515),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1398),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1399),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1486),
.A2(n_1437),
.B1(n_1501),
.B2(n_1479),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1484),
.A2(n_1505),
.B1(n_1417),
.B2(n_1361),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1403),
.Y(n_1551)
);

BUFx2_ASAP7_75t_SL g1552 ( 
.A(n_1364),
.Y(n_1552)
);

CKINVDCx11_ASAP7_75t_R g1553 ( 
.A(n_1379),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1410),
.A2(n_1418),
.B1(n_1432),
.B2(n_1464),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1518),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1476),
.A2(n_1375),
.B1(n_1354),
.B2(n_1432),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1495),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1465),
.B(n_1468),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1375),
.A2(n_1354),
.B1(n_1460),
.B2(n_1461),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1520),
.A2(n_1377),
.B1(n_1358),
.B2(n_1414),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1485),
.A2(n_1421),
.B1(n_1394),
.B2(n_1506),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1420),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1440),
.Y(n_1563)
);

CKINVDCx11_ASAP7_75t_R g1564 ( 
.A(n_1518),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1441),
.Y(n_1565)
);

CKINVDCx11_ASAP7_75t_R g1566 ( 
.A(n_1518),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1472),
.Y(n_1567)
);

BUFx2_ASAP7_75t_SL g1568 ( 
.A(n_1509),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1377),
.A2(n_1415),
.B1(n_1387),
.B2(n_1488),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1429),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1503),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1392),
.A2(n_1378),
.B1(n_1491),
.B2(n_1422),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1433),
.B(n_1439),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1433),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1389),
.A2(n_1368),
.B1(n_1434),
.B2(n_1449),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1512),
.A2(n_1499),
.B1(n_1506),
.B2(n_1425),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1429),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1441),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1496),
.Y(n_1579)
);

INVx6_ASAP7_75t_L g1580 ( 
.A(n_1447),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1508),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1438),
.B(n_1454),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1425),
.A2(n_1500),
.B1(n_1396),
.B2(n_1368),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1502),
.A2(n_1459),
.B1(n_1450),
.B2(n_1483),
.Y(n_1584)
);

BUFx4_ASAP7_75t_SL g1585 ( 
.A(n_1425),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1396),
.A2(n_1462),
.B1(n_1471),
.B2(n_1481),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1397),
.A2(n_1412),
.B1(n_1413),
.B2(n_1402),
.Y(n_1587)
);

CKINVDCx6p67_ASAP7_75t_R g1588 ( 
.A(n_1447),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1517),
.B(n_1446),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1380),
.A2(n_1381),
.B(n_1435),
.Y(n_1590)
);

BUFx8_ASAP7_75t_L g1591 ( 
.A(n_1412),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1519),
.B(n_1404),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1447),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1519),
.A2(n_1412),
.B1(n_1416),
.B2(n_1428),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1404),
.B(n_1422),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1474),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_SL g1597 ( 
.A1(n_1431),
.A2(n_1356),
.B1(n_1466),
.B2(n_1452),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1474),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1352),
.A2(n_1413),
.B1(n_1402),
.B2(n_1370),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1470),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1494),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1470),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1385),
.A2(n_1510),
.B1(n_1384),
.B2(n_1409),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1356),
.A2(n_1384),
.B1(n_1373),
.B2(n_1374),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1356),
.A2(n_1373),
.B1(n_1374),
.B2(n_1427),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1494),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1383),
.A2(n_1482),
.B1(n_1393),
.B2(n_1408),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1494),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1427),
.A2(n_1423),
.B1(n_1390),
.B2(n_1395),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1470),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1390),
.A2(n_1395),
.B1(n_1401),
.B2(n_1442),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1507),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1477),
.B(n_1436),
.Y(n_1613)
);

CKINVDCx6p67_ASAP7_75t_R g1614 ( 
.A(n_1443),
.Y(n_1614)
);

CKINVDCx11_ASAP7_75t_R g1615 ( 
.A(n_1444),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1443),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1463),
.A2(n_1445),
.B1(n_1367),
.B2(n_1366),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1363),
.A2(n_1511),
.B1(n_1493),
.B2(n_1372),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1451),
.A2(n_1511),
.B1(n_1444),
.B2(n_1357),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1365),
.A2(n_1357),
.B1(n_1405),
.B2(n_1400),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1357),
.A2(n_1405),
.B1(n_1400),
.B2(n_1498),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1498),
.B(n_1405),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1400),
.A2(n_1514),
.B1(n_1118),
.B2(n_1017),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1391),
.A2(n_1514),
.B1(n_1118),
.B2(n_1017),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1391),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1391),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1456),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1504),
.Y(n_1629)
);

BUFx2_ASAP7_75t_SL g1630 ( 
.A(n_1430),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1411),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1504),
.Y(n_1632)
);

INVx5_ASAP7_75t_L g1633 ( 
.A(n_1504),
.Y(n_1633)
);

BUFx10_ASAP7_75t_L g1634 ( 
.A(n_1371),
.Y(n_1634)
);

CKINVDCx11_ASAP7_75t_R g1635 ( 
.A(n_1430),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1453),
.B(n_856),
.Y(n_1636)
);

INVx6_ASAP7_75t_L g1637 ( 
.A(n_1504),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1456),
.Y(n_1638)
);

OAI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1514),
.A2(n_1458),
.B1(n_1118),
.B2(n_989),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1360),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1514),
.A2(n_1273),
.B1(n_1283),
.B2(n_1056),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1514),
.A2(n_1118),
.B(n_1273),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1411),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1456),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1456),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1362),
.B(n_903),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1456),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1407),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_SL g1652 ( 
.A1(n_1458),
.A2(n_1273),
.B1(n_1283),
.B2(n_1056),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1514),
.A2(n_1458),
.B1(n_1118),
.B2(n_989),
.Y(n_1654)
);

OA21x2_ASAP7_75t_L g1655 ( 
.A1(n_1451),
.A2(n_1386),
.B(n_1513),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1456),
.Y(n_1656)
);

BUFx12f_ASAP7_75t_L g1657 ( 
.A(n_1379),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1411),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1456),
.Y(n_1661)
);

BUFx4f_ASAP7_75t_SL g1662 ( 
.A(n_1379),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1456),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1514),
.A2(n_903),
.B1(n_1118),
.B2(n_1056),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1362),
.B(n_903),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1406),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1362),
.B(n_903),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1504),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1504),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1504),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1504),
.Y(n_1675)
);

CKINVDCx11_ASAP7_75t_R g1676 ( 
.A(n_1430),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1514),
.A2(n_1273),
.B1(n_1283),
.B2(n_1056),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1456),
.Y(n_1678)
);

NAND2x1p5_ASAP7_75t_L g1679 ( 
.A(n_1507),
.B(n_1230),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1680)
);

BUFx8_ASAP7_75t_L g1681 ( 
.A(n_1379),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1504),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1514),
.A2(n_1273),
.B1(n_1283),
.B2(n_1056),
.Y(n_1684)
);

CKINVDCx11_ASAP7_75t_R g1685 ( 
.A(n_1430),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1475),
.A2(n_1283),
.B1(n_1273),
.B2(n_1056),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1456),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1411),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1456),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1406),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1456),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1514),
.A2(n_1118),
.B(n_1273),
.Y(n_1694)
);

CKINVDCx6p67_ASAP7_75t_R g1695 ( 
.A(n_1379),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1456),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1458),
.A2(n_1273),
.B1(n_1283),
.B2(n_1056),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1371),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1430),
.Y(n_1699)
);

CKINVDCx6p67_ASAP7_75t_R g1700 ( 
.A(n_1379),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1514),
.A2(n_1118),
.B1(n_1017),
.B2(n_1273),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1514),
.A2(n_1458),
.B1(n_1118),
.B2(n_989),
.Y(n_1702)
);

INVx6_ASAP7_75t_L g1703 ( 
.A(n_1504),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1371),
.Y(n_1704)
);

BUFx8_ASAP7_75t_L g1705 ( 
.A(n_1379),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1612),
.Y(n_1706)
);

OAI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1642),
.A2(n_1684),
.B1(n_1677),
.B2(n_1643),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1624),
.B(n_1546),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1612),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1557),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1686),
.B(n_1694),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1557),
.B(n_1625),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1565),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1527),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1614),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1627),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1626),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1624),
.B(n_1600),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1635),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1536),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1602),
.B(n_1610),
.Y(n_1722)
);

NAND2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1567),
.B(n_1589),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1578),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1616),
.B(n_1592),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1622),
.B(n_1595),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1623),
.B(n_1529),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1669),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1524),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1631),
.Y(n_1730)
);

BUFx12f_ASAP7_75t_L g1731 ( 
.A(n_1676),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1638),
.Y(n_1732)
);

OAI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1641),
.A2(n_1653),
.B1(n_1647),
.B2(n_1659),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1619),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1685),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1619),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1649),
.B(n_1668),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1652),
.A2(n_1697),
.B1(n_1680),
.B2(n_1682),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1658),
.A2(n_1667),
.B(n_1663),
.C(n_1666),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1591),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1604),
.B(n_1645),
.Y(n_1742)
);

AO31x2_ASAP7_75t_L g1743 ( 
.A1(n_1618),
.A2(n_1603),
.A3(n_1583),
.B(n_1599),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1646),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1650),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1656),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1661),
.B(n_1665),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1670),
.B(n_1523),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1678),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1539),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1644),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1687),
.B(n_1689),
.Y(n_1752)
);

BUFx4f_ASAP7_75t_SL g1753 ( 
.A(n_1657),
.Y(n_1753)
);

AO21x2_ASAP7_75t_L g1754 ( 
.A1(n_1617),
.A2(n_1587),
.B(n_1550),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1692),
.B(n_1696),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1690),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1698),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1628),
.B(n_1648),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1537),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1562),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1655),
.Y(n_1761)
);

CKINVDCx8_ASAP7_75t_R g1762 ( 
.A(n_1630),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1591),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1581),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1563),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1621),
.B(n_1560),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1541),
.Y(n_1767)
);

AO21x2_ASAP7_75t_L g1768 ( 
.A1(n_1587),
.A2(n_1550),
.B(n_1613),
.Y(n_1768)
);

CKINVDCx9p33_ASAP7_75t_R g1769 ( 
.A(n_1660),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1543),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1628),
.B(n_1648),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1538),
.Y(n_1772)
);

AO21x2_ASAP7_75t_L g1773 ( 
.A1(n_1607),
.A2(n_1572),
.B(n_1576),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1547),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1538),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1640),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1664),
.B(n_1673),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1679),
.Y(n_1778)
);

CKINVDCx12_ASAP7_75t_R g1779 ( 
.A(n_1636),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1655),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1571),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1621),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1620),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1620),
.Y(n_1784)
);

AO21x2_ASAP7_75t_L g1785 ( 
.A1(n_1639),
.A2(n_1654),
.B(n_1702),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1573),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1615),
.Y(n_1787)
);

AO21x2_ASAP7_75t_L g1788 ( 
.A1(n_1639),
.A2(n_1702),
.B(n_1654),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1582),
.A2(n_1535),
.B1(n_1682),
.B2(n_1680),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1574),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1688),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1558),
.Y(n_1792)
);

AOI21xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1664),
.A2(n_1701),
.B(n_1673),
.Y(n_1793)
);

OR2x6_ASAP7_75t_L g1794 ( 
.A(n_1590),
.B(n_1577),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1524),
.Y(n_1795)
);

BUFx3_ASAP7_75t_L g1796 ( 
.A(n_1579),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1585),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1552),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1559),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1691),
.A2(n_1693),
.B(n_1701),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1691),
.B(n_1693),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1605),
.B(n_1534),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1559),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1585),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1629),
.Y(n_1805)
);

OAI21xp33_ASAP7_75t_SL g1806 ( 
.A1(n_1528),
.A2(n_1525),
.B(n_1532),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1629),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1629),
.Y(n_1808)
);

BUFx2_ASAP7_75t_SL g1809 ( 
.A(n_1633),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1605),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1632),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1632),
.Y(n_1812)
);

CKINVDCx8_ASAP7_75t_R g1813 ( 
.A(n_1704),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1534),
.B(n_1525),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1609),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1611),
.Y(n_1816)
);

OAI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1586),
.A2(n_1575),
.B(n_1549),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1528),
.B(n_1594),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1549),
.A2(n_1532),
.B(n_1544),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1594),
.B(n_1544),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1575),
.Y(n_1821)
);

AO21x2_ASAP7_75t_L g1822 ( 
.A1(n_1554),
.A2(n_1586),
.B(n_1597),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1671),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1633),
.B(n_1533),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1522),
.B(n_1526),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1545),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1569),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1671),
.Y(n_1828)
);

OR2x6_ASAP7_75t_L g1829 ( 
.A(n_1577),
.B(n_1568),
.Y(n_1829)
);

OAI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1569),
.A2(n_1556),
.B(n_1522),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1584),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1556),
.A2(n_1542),
.B(n_1561),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1672),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1672),
.B(n_1674),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1672),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1540),
.B(n_1633),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1674),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1577),
.A2(n_1570),
.B1(n_1662),
.B2(n_1700),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1538),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1674),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1699),
.A2(n_1695),
.B1(n_1662),
.B2(n_1651),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1588),
.A2(n_1545),
.B(n_1637),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1674),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1606),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1606),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1545),
.A2(n_1637),
.B(n_1703),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1596),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1596),
.Y(n_1848)
);

OAI21xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1675),
.A2(n_1683),
.B(n_1530),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1606),
.Y(n_1850)
);

INVx4_ASAP7_75t_L g1851 ( 
.A(n_1675),
.Y(n_1851)
);

NAND2x1_ASAP7_75t_L g1852 ( 
.A(n_1637),
.B(n_1703),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1598),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1598),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1593),
.B(n_1608),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1703),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1580),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1580),
.Y(n_1858)
);

INVx4_ASAP7_75t_L g1859 ( 
.A(n_1564),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1555),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1555),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1707),
.A2(n_1705),
.B1(n_1681),
.B2(n_1553),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1737),
.B(n_1601),
.Y(n_1863)
);

AO21x2_ASAP7_75t_L g1864 ( 
.A1(n_1819),
.A2(n_1566),
.B(n_1521),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1720),
.Y(n_1865)
);

INVxp67_ASAP7_75t_SL g1866 ( 
.A(n_1728),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1769),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1806),
.A2(n_1634),
.B(n_1531),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1706),
.B(n_1634),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1738),
.A2(n_1681),
.B1(n_1705),
.B2(n_1531),
.Y(n_1870)
);

INVxp67_ASAP7_75t_SL g1871 ( 
.A(n_1756),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1748),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1792),
.B(n_1759),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1720),
.Y(n_1874)
);

AO32x2_ASAP7_75t_L g1875 ( 
.A1(n_1706),
.A2(n_1768),
.A3(n_1754),
.B1(n_1726),
.B2(n_1725),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1709),
.B(n_1721),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1744),
.Y(n_1877)
);

O2A1O1Ixp33_ASAP7_75t_SL g1878 ( 
.A1(n_1800),
.A2(n_1793),
.B(n_1733),
.C(n_1801),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1709),
.B(n_1721),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1825),
.B(n_1799),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1718),
.B(n_1742),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1744),
.Y(n_1882)
);

A2O1A1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1740),
.A2(n_1789),
.B(n_1830),
.C(n_1711),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1742),
.B(n_1815),
.Y(n_1884)
);

AND2x2_ASAP7_75t_SL g1885 ( 
.A(n_1741),
.B(n_1763),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1726),
.B(n_1710),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1745),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1745),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1815),
.B(n_1708),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1709),
.B(n_1721),
.Y(n_1890)
);

O2A1O1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1758),
.A2(n_1777),
.B(n_1771),
.C(n_1814),
.Y(n_1891)
);

AOI221xp5_ASAP7_75t_L g1892 ( 
.A1(n_1820),
.A2(n_1739),
.B1(n_1818),
.B2(n_1803),
.C(n_1827),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1782),
.B(n_1734),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1782),
.B(n_1736),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1825),
.B(n_1781),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1831),
.A2(n_1773),
.B(n_1827),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1785),
.A2(n_1788),
.B1(n_1739),
.B2(n_1802),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1747),
.B(n_1752),
.Y(n_1898)
);

OAI221xp5_ASAP7_75t_L g1899 ( 
.A1(n_1794),
.A2(n_1831),
.B1(n_1838),
.B2(n_1798),
.C(n_1802),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1820),
.B(n_1783),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1785),
.A2(n_1788),
.B(n_1773),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1730),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1794),
.B(n_1727),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1783),
.B(n_1784),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1784),
.B(n_1810),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1747),
.B(n_1752),
.Y(n_1906)
);

AOI22x1_ASAP7_75t_SL g1907 ( 
.A1(n_1735),
.A2(n_1719),
.B1(n_1787),
.B2(n_1859),
.Y(n_1907)
);

INVx4_ASAP7_75t_L g1908 ( 
.A(n_1829),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1727),
.B(n_1741),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1763),
.B(n_1786),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1760),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1810),
.B(n_1754),
.Y(n_1912)
);

BUFx4f_ASAP7_75t_SL g1913 ( 
.A(n_1731),
.Y(n_1913)
);

OA21x2_ASAP7_75t_L g1914 ( 
.A1(n_1761),
.A2(n_1780),
.B(n_1817),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1829),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1821),
.B(n_1830),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1816),
.B(n_1746),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1818),
.A2(n_1821),
.B1(n_1768),
.B2(n_1816),
.C(n_1773),
.Y(n_1918)
);

O2A1O1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1794),
.A2(n_1836),
.B(n_1788),
.C(n_1785),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1729),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1760),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1751),
.A2(n_1791),
.B1(n_1822),
.B2(n_1766),
.C(n_1714),
.Y(n_1922)
);

AO32x2_ASAP7_75t_L g1923 ( 
.A1(n_1772),
.A2(n_1839),
.A3(n_1775),
.B1(n_1712),
.B2(n_1722),
.Y(n_1923)
);

AO32x2_ASAP7_75t_L g1924 ( 
.A1(n_1772),
.A2(n_1839),
.A3(n_1775),
.B1(n_1712),
.B2(n_1722),
.Y(n_1924)
);

NAND3xp33_ASAP7_75t_L g1925 ( 
.A(n_1794),
.B(n_1849),
.C(n_1765),
.Y(n_1925)
);

AO32x2_ASAP7_75t_L g1926 ( 
.A1(n_1764),
.A2(n_1859),
.A3(n_1851),
.B1(n_1761),
.B2(n_1780),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1749),
.B(n_1743),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1749),
.B(n_1743),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1743),
.B(n_1755),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1755),
.B(n_1834),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1832),
.B(n_1829),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1716),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1743),
.B(n_1732),
.Y(n_1933)
);

AO32x2_ASAP7_75t_L g1934 ( 
.A1(n_1764),
.A2(n_1859),
.A3(n_1851),
.B1(n_1743),
.B2(n_1724),
.Y(n_1934)
);

AO21x2_ASAP7_75t_L g1935 ( 
.A1(n_1817),
.A2(n_1822),
.B(n_1713),
.Y(n_1935)
);

OA21x2_ASAP7_75t_L g1936 ( 
.A1(n_1717),
.A2(n_1832),
.B(n_1715),
.Y(n_1936)
);

AOI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1822),
.A2(n_1774),
.B1(n_1776),
.B2(n_1770),
.C(n_1767),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1796),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1762),
.A2(n_1804),
.B1(n_1797),
.B2(n_1841),
.Y(n_1939)
);

OAI21xp33_ASAP7_75t_SL g1940 ( 
.A1(n_1842),
.A2(n_1846),
.B(n_1851),
.Y(n_1940)
);

OA21x2_ASAP7_75t_L g1941 ( 
.A1(n_1844),
.A2(n_1843),
.B(n_1835),
.Y(n_1941)
);

OA21x2_ASAP7_75t_L g1942 ( 
.A1(n_1844),
.A2(n_1843),
.B(n_1835),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1790),
.B(n_1723),
.Y(n_1943)
);

A2O1A1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1809),
.A2(n_1842),
.B(n_1846),
.C(n_1729),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1723),
.B(n_1796),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1778),
.B(n_1731),
.Y(n_1946)
);

AO21x2_ASAP7_75t_L g1947 ( 
.A1(n_1853),
.A2(n_1854),
.B(n_1860),
.Y(n_1947)
);

AND2x4_ASAP7_75t_SL g1948 ( 
.A(n_1869),
.B(n_1908),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1920),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1929),
.B(n_1853),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1866),
.B(n_1847),
.Y(n_1951)
);

BUFx3_ASAP7_75t_L g1952 ( 
.A(n_1920),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1876),
.B(n_1823),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1876),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1929),
.B(n_1854),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1886),
.B(n_1848),
.Y(n_1956)
);

INVx4_ASAP7_75t_L g1957 ( 
.A(n_1946),
.Y(n_1957)
);

AOI221x1_ASAP7_75t_SL g1958 ( 
.A1(n_1896),
.A2(n_1855),
.B1(n_1858),
.B2(n_1857),
.C(n_1856),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1877),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1912),
.B(n_1808),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1912),
.B(n_1808),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1871),
.B(n_1807),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1895),
.B(n_1833),
.Y(n_1963)
);

NAND2x1p5_ASAP7_75t_L g1964 ( 
.A(n_1908),
.B(n_1861),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1917),
.Y(n_1965)
);

NOR2xp67_ASAP7_75t_L g1966 ( 
.A(n_1925),
.B(n_1719),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1882),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1872),
.B(n_1762),
.Y(n_1968)
);

AND2x4_ASAP7_75t_SL g1969 ( 
.A(n_1869),
.B(n_1735),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1941),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1881),
.B(n_1833),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1887),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1888),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_1869),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1942),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1880),
.B(n_1840),
.Y(n_1976)
);

AND2x2_ASAP7_75t_SL g1977 ( 
.A(n_1897),
.B(n_1824),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1942),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1906),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1881),
.B(n_1840),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1927),
.B(n_1812),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1889),
.B(n_1837),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1873),
.B(n_1837),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1899),
.A2(n_1753),
.B1(n_1795),
.B2(n_1750),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1889),
.B(n_1845),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1942),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1900),
.B(n_1930),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1900),
.B(n_1906),
.Y(n_1988)
);

OAI222xp33_ASAP7_75t_L g1989 ( 
.A1(n_1862),
.A2(n_1856),
.B1(n_1858),
.B2(n_1857),
.C1(n_1813),
.C2(n_1850),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1892),
.A2(n_1750),
.B1(n_1861),
.B2(n_1824),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1884),
.B(n_1811),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1928),
.B(n_1933),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1911),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1921),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1879),
.Y(n_1995)
);

BUFx3_ASAP7_75t_L g1996 ( 
.A(n_1946),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1916),
.B(n_1805),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1865),
.Y(n_1998)
);

NOR2x1_ASAP7_75t_L g1999 ( 
.A(n_1947),
.B(n_1828),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1902),
.B(n_1779),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1916),
.B(n_1811),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1874),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1868),
.B(n_1757),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1874),
.Y(n_2004)
);

INVx3_ASAP7_75t_L g2005 ( 
.A(n_1890),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1938),
.Y(n_2006)
);

AND2x2_ASAP7_75t_SL g2007 ( 
.A(n_1977),
.B(n_1922),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1959),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1950),
.B(n_1935),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1960),
.Y(n_2010)
);

AOI31xp33_ASAP7_75t_L g2011 ( 
.A1(n_2003),
.A2(n_1878),
.A3(n_1939),
.B(n_1931),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1959),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1954),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1954),
.Y(n_2014)
);

INVxp67_ASAP7_75t_L g2015 ( 
.A(n_1956),
.Y(n_2015)
);

AO21x2_ASAP7_75t_L g2016 ( 
.A1(n_1970),
.A2(n_1901),
.B(n_1944),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1977),
.A2(n_1931),
.B1(n_1897),
.B2(n_1864),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1983),
.B(n_1918),
.Y(n_2018)
);

OAI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_1984),
.A2(n_1878),
.B1(n_1883),
.B2(n_1870),
.C(n_1891),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1998),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1957),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1966),
.A2(n_1883),
.B(n_1919),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1960),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1992),
.B(n_1988),
.Y(n_2024)
);

OAI221xp5_ASAP7_75t_L g2025 ( 
.A1(n_1958),
.A2(n_1867),
.B1(n_1944),
.B2(n_1945),
.C(n_1946),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1998),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1992),
.B(n_1923),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2002),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1988),
.B(n_1923),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2002),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1954),
.B(n_1890),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1989),
.A2(n_1937),
.B(n_1864),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1950),
.B(n_1955),
.Y(n_2033)
);

INVx1_ASAP7_75t_SL g2034 ( 
.A(n_1969),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1995),
.B(n_2005),
.Y(n_2035)
);

AND4x1_ASAP7_75t_L g2036 ( 
.A(n_1968),
.B(n_1945),
.C(n_1903),
.D(n_1907),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1976),
.B(n_1898),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1995),
.B(n_1923),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1969),
.B(n_1946),
.Y(n_2039)
);

INVxp67_ASAP7_75t_SL g2040 ( 
.A(n_1999),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2004),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_SL g2042 ( 
.A(n_1957),
.B(n_1913),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1951),
.B(n_1963),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_L g2044 ( 
.A(n_1957),
.B(n_1940),
.C(n_2000),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1995),
.B(n_1923),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1967),
.Y(n_2046)
);

NOR2x1_ASAP7_75t_L g2047 ( 
.A(n_1999),
.B(n_1947),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1972),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_2005),
.Y(n_2049)
);

OAI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_1990),
.A2(n_1885),
.B1(n_1903),
.B2(n_1915),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1962),
.B(n_1987),
.Y(n_2051)
);

AOI33xp33_ASAP7_75t_L g2052 ( 
.A1(n_1972),
.A2(n_1904),
.A3(n_1905),
.B1(n_1932),
.B2(n_1994),
.B3(n_1993),
.Y(n_2052)
);

NOR2x1_ASAP7_75t_L g2053 ( 
.A(n_1949),
.B(n_1952),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1961),
.B(n_1935),
.Y(n_2054)
);

INVx4_ASAP7_75t_L g2055 ( 
.A(n_1996),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2005),
.B(n_1924),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1973),
.Y(n_2057)
);

AND2x4_ASAP7_75t_SL g2058 ( 
.A(n_1953),
.B(n_1908),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1979),
.B(n_1924),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_L g2060 ( 
.A(n_1997),
.B(n_1936),
.C(n_1943),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1997),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1979),
.B(n_1924),
.Y(n_2062)
);

INVxp67_ASAP7_75t_SL g2063 ( 
.A(n_2001),
.Y(n_2063)
);

AOI31xp33_ASAP7_75t_L g2064 ( 
.A1(n_1964),
.A2(n_1909),
.A3(n_1910),
.B(n_1863),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_1974),
.Y(n_2065)
);

AOI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2006),
.A2(n_1905),
.B1(n_1894),
.B2(n_1893),
.C(n_1943),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_1965),
.B(n_1914),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2018),
.B(n_1987),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_2007),
.B(n_2022),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2009),
.B(n_1975),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2020),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2009),
.B(n_1975),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2052),
.B(n_2063),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2027),
.B(n_1875),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2027),
.B(n_2038),
.Y(n_2075)
);

BUFx3_ASAP7_75t_L g2076 ( 
.A(n_2016),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_2067),
.B(n_1978),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2015),
.B(n_1982),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_2020),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2045),
.B(n_1875),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2026),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_2045),
.B(n_1978),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2056),
.B(n_1875),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_2040),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2056),
.B(n_1934),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2067),
.B(n_1986),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2029),
.B(n_1934),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2026),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2054),
.B(n_1986),
.Y(n_2089)
);

NAND2x1p5_ASAP7_75t_L g2090 ( 
.A(n_2047),
.B(n_1936),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_2028),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2029),
.B(n_1934),
.Y(n_2092)
);

NOR2xp67_ASAP7_75t_L g2093 ( 
.A(n_2060),
.B(n_2001),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2028),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2046),
.B(n_2048),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2059),
.B(n_1934),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2059),
.B(n_1977),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2048),
.B(n_2057),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2054),
.B(n_1981),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2030),
.Y(n_2100)
);

AND2x2_ASAP7_75t_SL g2101 ( 
.A(n_2007),
.B(n_1936),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2062),
.B(n_1971),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2062),
.B(n_1971),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2030),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2024),
.B(n_1980),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2008),
.B(n_1985),
.Y(n_2106)
);

BUFx2_ASAP7_75t_L g2107 ( 
.A(n_2021),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2024),
.B(n_1980),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2035),
.B(n_1926),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_2041),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_2064),
.B(n_1885),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2035),
.B(n_2061),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2041),
.Y(n_2113)
);

AOI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2069),
.A2(n_2019),
.B(n_2032),
.C(n_2025),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2079),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2068),
.B(n_2066),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2068),
.B(n_2043),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2073),
.B(n_2033),
.Y(n_2118)
);

OAI21xp33_ASAP7_75t_L g2119 ( 
.A1(n_2069),
.A2(n_2017),
.B(n_2011),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_2111),
.A2(n_2044),
.B1(n_2101),
.B2(n_2050),
.Y(n_2120)
);

OAI22xp33_ASAP7_75t_R g2121 ( 
.A1(n_2101),
.A2(n_2036),
.B1(n_2039),
.B2(n_2034),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2076),
.Y(n_2122)
);

O2A1O1Ixp33_ASAP7_75t_SL g2123 ( 
.A1(n_2111),
.A2(n_2065),
.B(n_2013),
.C(n_2014),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2079),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2097),
.B(n_2031),
.Y(n_2125)
);

HB1xp67_ASAP7_75t_L g2126 ( 
.A(n_2084),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2084),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2091),
.Y(n_2128)
);

INVx4_ASAP7_75t_L g2129 ( 
.A(n_2107),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2097),
.B(n_2031),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2091),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2097),
.B(n_2031),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2110),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_2084),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2110),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2073),
.B(n_2051),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_2107),
.B(n_2053),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2107),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2076),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2099),
.B(n_2033),
.Y(n_2140)
);

NAND4xp25_ASAP7_75t_L g2141 ( 
.A(n_2093),
.B(n_2042),
.C(n_2021),
.D(n_2055),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2112),
.B(n_2013),
.Y(n_2142)
);

INVx1_ASAP7_75t_SL g2143 ( 
.A(n_2101),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2076),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2081),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2112),
.B(n_2075),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2105),
.B(n_2037),
.Y(n_2147)
);

NAND3xp33_ASAP7_75t_SL g2148 ( 
.A(n_2090),
.B(n_2055),
.C(n_2021),
.Y(n_2148)
);

INVxp67_ASAP7_75t_L g2149 ( 
.A(n_2101),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2112),
.B(n_2014),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2081),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2093),
.B(n_2055),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2105),
.B(n_2010),
.Y(n_2153)
);

OAI21xp33_ASAP7_75t_SL g2154 ( 
.A1(n_2087),
.A2(n_2049),
.B(n_2065),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2081),
.Y(n_2155)
);

NOR2x1_ASAP7_75t_L g2156 ( 
.A(n_2076),
.B(n_1996),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2075),
.B(n_2049),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2075),
.B(n_2023),
.Y(n_2158)
);

NOR2x1_ASAP7_75t_L g2159 ( 
.A(n_2095),
.B(n_1949),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2082),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2094),
.Y(n_2161)
);

AND2x4_ASAP7_75t_L g2162 ( 
.A(n_2094),
.B(n_2016),
.Y(n_2162)
);

AOI32xp33_ASAP7_75t_L g2163 ( 
.A1(n_2087),
.A2(n_1948),
.A3(n_2058),
.B1(n_1974),
.B2(n_1991),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2094),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2102),
.B(n_2058),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2136),
.B(n_2087),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2146),
.B(n_2109),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_2129),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2116),
.B(n_2092),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2146),
.B(n_2109),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2125),
.B(n_2130),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2125),
.B(n_2096),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2114),
.B(n_2092),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2130),
.B(n_2132),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2132),
.B(n_2109),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2145),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2145),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2158),
.B(n_2102),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2162),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2156),
.B(n_2096),
.Y(n_2180)
);

INVxp67_ASAP7_75t_SL g2181 ( 
.A(n_2126),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2151),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2151),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2117),
.B(n_2092),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2118),
.B(n_2099),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2158),
.B(n_2157),
.Y(n_2186)
);

NOR2x1_ASAP7_75t_L g2187 ( 
.A(n_2129),
.B(n_2100),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2155),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2162),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2155),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2118),
.B(n_2085),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2159),
.B(n_2096),
.Y(n_2192)
);

NAND2x1_ASAP7_75t_SL g2193 ( 
.A(n_2120),
.B(n_2085),
.Y(n_2193)
);

OA211x2_ASAP7_75t_L g2194 ( 
.A1(n_2119),
.A2(n_1852),
.B(n_2095),
.C(n_2098),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2161),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2157),
.B(n_2102),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2138),
.B(n_2085),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2147),
.B(n_2099),
.Y(n_2198)
);

AOI331xp33_ASAP7_75t_L g2199 ( 
.A1(n_2115),
.A2(n_2100),
.A3(n_2088),
.B1(n_2071),
.B2(n_2104),
.B3(n_2113),
.C1(n_2012),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2165),
.B(n_2103),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2153),
.B(n_2098),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2162),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2127),
.B(n_2074),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_2140),
.B(n_2078),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2161),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2164),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2134),
.B(n_2074),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2173),
.B(n_2129),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2173),
.B(n_2115),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2171),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2181),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2193),
.B(n_2143),
.Y(n_2212)
);

INVx1_ASAP7_75t_SL g2213 ( 
.A(n_2193),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2181),
.B(n_2124),
.Y(n_2214)
);

AOI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2169),
.A2(n_2149),
.B1(n_2152),
.B2(n_2123),
.C(n_2141),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2176),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2194),
.A2(n_2121),
.B1(n_2148),
.B2(n_2154),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2176),
.Y(n_2218)
);

AOI32xp33_ASAP7_75t_L g2219 ( 
.A1(n_2180),
.A2(n_2137),
.A3(n_2121),
.B1(n_2142),
.B2(n_2150),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2171),
.B(n_2137),
.Y(n_2220)
);

AOI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2194),
.A2(n_2137),
.B1(n_2142),
.B2(n_2150),
.Y(n_2221)
);

OAI221xp5_ASAP7_75t_L g2222 ( 
.A1(n_2169),
.A2(n_2163),
.B1(n_2090),
.B2(n_2135),
.C(n_2131),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2191),
.B(n_2140),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2177),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2177),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_2180),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2182),
.Y(n_2227)
);

AOI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_2199),
.A2(n_2163),
.B(n_2139),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2199),
.B(n_2124),
.Y(n_2229)
);

OAI321xp33_ASAP7_75t_L g2230 ( 
.A1(n_2180),
.A2(n_2122),
.A3(n_2139),
.B1(n_2144),
.B2(n_2135),
.C(n_2133),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2182),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2183),
.Y(n_2232)
);

OAI21xp5_ASAP7_75t_SL g2233 ( 
.A1(n_2192),
.A2(n_2090),
.B(n_2165),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2174),
.B(n_2105),
.Y(n_2234)
);

AOI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2192),
.A2(n_2122),
.B1(n_2144),
.B2(n_2128),
.C(n_2133),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2183),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2174),
.B(n_2108),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2213),
.B(n_2186),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_2217),
.B(n_2192),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2211),
.B(n_2186),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2216),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2208),
.B(n_2200),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2219),
.A2(n_2166),
.B1(n_2191),
.B2(n_2187),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2230),
.A2(n_2228),
.B(n_2212),
.Y(n_2244)
);

NOR3xp33_ASAP7_75t_SL g2245 ( 
.A(n_2222),
.B(n_2166),
.C(n_2197),
.Y(n_2245)
);

OAI21xp33_ASAP7_75t_L g2246 ( 
.A1(n_2215),
.A2(n_2197),
.B(n_2185),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2210),
.B(n_2208),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2226),
.B(n_2200),
.Y(n_2248)
);

INVxp67_ASAP7_75t_L g2249 ( 
.A(n_2209),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_2209),
.B(n_2204),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2229),
.A2(n_2187),
.B(n_2168),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_2223),
.B(n_2204),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2220),
.B(n_2178),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2220),
.B(n_2178),
.Y(n_2254)
);

O2A1O1Ixp5_ASAP7_75t_L g2255 ( 
.A1(n_2229),
.A2(n_2168),
.B(n_2179),
.C(n_2202),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2235),
.A2(n_2185),
.B1(n_2201),
.B2(n_2207),
.C(n_2203),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2234),
.B(n_2172),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2214),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2237),
.B(n_2172),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2214),
.B(n_2172),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2240),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2238),
.B(n_2175),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2253),
.B(n_2175),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_L g2264 ( 
.A(n_2258),
.B(n_2233),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2254),
.Y(n_2265)
);

XNOR2x2_ASAP7_75t_L g2266 ( 
.A(n_2244),
.B(n_2221),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2247),
.B(n_2168),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2248),
.Y(n_2268)
);

O2A1O1Ixp33_ASAP7_75t_L g2269 ( 
.A1(n_2239),
.A2(n_2168),
.B(n_2232),
.C(n_2231),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2251),
.B(n_2218),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2260),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2251),
.B(n_2224),
.Y(n_2272)
);

XOR2xp5_ASAP7_75t_L g2273 ( 
.A(n_2243),
.B(n_1757),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_2246),
.A2(n_2236),
.B1(n_2227),
.B2(n_2225),
.Y(n_2274)
);

OAI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2255),
.A2(n_2207),
.B(n_2203),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2250),
.B(n_2196),
.Y(n_2276)
);

XOR2xp5_ASAP7_75t_L g2277 ( 
.A(n_2273),
.B(n_2242),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2265),
.B(n_2249),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2263),
.B(n_2252),
.Y(n_2279)
);

CKINVDCx20_ASAP7_75t_L g2280 ( 
.A(n_2266),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2267),
.B(n_2245),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2267),
.Y(n_2282)
);

INVx2_ASAP7_75t_SL g2283 ( 
.A(n_2270),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2268),
.B(n_2257),
.Y(n_2284)
);

OAI31xp33_ASAP7_75t_SL g2285 ( 
.A1(n_2264),
.A2(n_2256),
.A3(n_2241),
.B(n_2189),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2269),
.B(n_2259),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2262),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2264),
.B(n_2196),
.Y(n_2288)
);

NOR2x1_ASAP7_75t_SL g2289 ( 
.A(n_2272),
.B(n_2179),
.Y(n_2289)
);

AOI221x1_ASAP7_75t_L g2290 ( 
.A1(n_2282),
.A2(n_2261),
.B1(n_2271),
.B2(n_2275),
.C(n_2276),
.Y(n_2290)
);

AO22x2_ASAP7_75t_L g2291 ( 
.A1(n_2282),
.A2(n_2286),
.B1(n_2283),
.B2(n_2277),
.Y(n_2291)
);

AOI211xp5_ASAP7_75t_L g2292 ( 
.A1(n_2285),
.A2(n_2269),
.B(n_2274),
.C(n_2206),
.Y(n_2292)
);

NAND4xp25_ASAP7_75t_L g2293 ( 
.A(n_2288),
.B(n_2274),
.C(n_2189),
.D(n_2179),
.Y(n_2293)
);

NAND5xp2_ASAP7_75t_L g2294 ( 
.A(n_2279),
.B(n_2206),
.C(n_2190),
.D(n_2205),
.E(n_2195),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2280),
.A2(n_2189),
.B1(n_2202),
.B2(n_2131),
.Y(n_2295)
);

OA22x2_ASAP7_75t_L g2296 ( 
.A1(n_2286),
.A2(n_2202),
.B1(n_2205),
.B2(n_2188),
.Y(n_2296)
);

AOI221x1_ASAP7_75t_L g2297 ( 
.A1(n_2278),
.A2(n_2188),
.B1(n_2195),
.B2(n_2190),
.C(n_2128),
.Y(n_2297)
);

AOI311xp33_ASAP7_75t_L g2298 ( 
.A1(n_2287),
.A2(n_2184),
.A3(n_2164),
.B(n_2100),
.C(n_2088),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2292),
.B(n_2283),
.Y(n_2299)
);

AOI211xp5_ASAP7_75t_L g2300 ( 
.A1(n_2293),
.A2(n_2281),
.B(n_2278),
.C(n_2284),
.Y(n_2300)
);

AOI221xp5_ASAP7_75t_L g2301 ( 
.A1(n_2291),
.A2(n_2289),
.B1(n_2184),
.B2(n_2201),
.C(n_2170),
.Y(n_2301)
);

AOI221x1_ASAP7_75t_L g2302 ( 
.A1(n_2294),
.A2(n_2170),
.B1(n_2167),
.B2(n_2160),
.C(n_2104),
.Y(n_2302)
);

AO22x1_ASAP7_75t_L g2303 ( 
.A1(n_2296),
.A2(n_2167),
.B1(n_1813),
.B2(n_2160),
.Y(n_2303)
);

NAND4xp25_ASAP7_75t_L g2304 ( 
.A(n_2290),
.B(n_2198),
.C(n_1826),
.D(n_2078),
.Y(n_2304)
);

OAI211xp5_ASAP7_75t_SL g2305 ( 
.A1(n_2295),
.A2(n_2198),
.B(n_2106),
.C(n_2086),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2297),
.A2(n_2090),
.B(n_2086),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2300),
.B(n_2298),
.Y(n_2307)
);

NAND4xp75_ASAP7_75t_L g2308 ( 
.A(n_2299),
.B(n_2074),
.C(n_2083),
.D(n_2080),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2303),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2306),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2301),
.B(n_2304),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2302),
.Y(n_2312)
);

OAI211xp5_ASAP7_75t_SL g2313 ( 
.A1(n_2309),
.A2(n_2305),
.B(n_2106),
.C(n_2086),
.Y(n_2313)
);

NAND3xp33_ASAP7_75t_L g2314 ( 
.A(n_2312),
.B(n_2077),
.C(n_2070),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_2311),
.B(n_2082),
.Y(n_2315)
);

NOR2x1p5_ASAP7_75t_L g2316 ( 
.A(n_2310),
.B(n_1826),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2315),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2317),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2318),
.A2(n_2308),
.B1(n_2314),
.B2(n_2310),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2318),
.Y(n_2320)
);

OAI31xp67_ASAP7_75t_SL g2321 ( 
.A1(n_2320),
.A2(n_2316),
.A3(n_2311),
.B(n_2307),
.Y(n_2321)
);

AOI22x1_ASAP7_75t_L g2322 ( 
.A1(n_2319),
.A2(n_2307),
.B1(n_2313),
.B2(n_2090),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2322),
.Y(n_2323)
);

AOI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2321),
.A2(n_2082),
.B1(n_2080),
.B2(n_2083),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2323),
.Y(n_2325)
);

OAI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2325),
.A2(n_2324),
.B(n_2077),
.Y(n_2326)
);

XNOR2xp5_ASAP7_75t_L g2327 ( 
.A(n_2326),
.B(n_1852),
.Y(n_2327)
);

OAI221xp5_ASAP7_75t_R g2328 ( 
.A1(n_2327),
.A2(n_2077),
.B1(n_2070),
.B2(n_2072),
.C(n_2089),
.Y(n_2328)
);

AOI211xp5_ASAP7_75t_L g2329 ( 
.A1(n_2328),
.A2(n_2070),
.B(n_2072),
.C(n_2089),
.Y(n_2329)
);


endmodule