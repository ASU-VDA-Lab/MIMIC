module fake_netlist_5_2453_n_1428 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1428);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1428;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_159),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_166),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_195),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_144),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_102),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_26),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_212),
.B(n_223),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_160),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_192),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_207),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_11),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_146),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_145),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_53),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_269),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_342),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_229),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_288),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_176),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_190),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_44),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_316),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_209),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_108),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_307),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_167),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_304),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_85),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_134),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_367),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_188),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_327),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_20),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_161),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_257),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_48),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_148),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_164),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_114),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_41),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_72),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_25),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_291),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_0),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_163),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_136),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_371),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_353),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_306),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_208),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_149),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_118),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_9),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_197),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_97),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_61),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_278),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_273),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_81),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_279),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_54),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_328),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_4),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_178),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_191),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_251),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_244),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_4),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_294),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_247),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_84),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_369),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_143),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_222),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_350),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_334),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_21),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_153),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_250),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_115),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_182),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_87),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_339),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_147),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_183),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_337),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_201),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_346),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_93),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_245),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_354),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_35),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_71),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_100),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_165),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_315),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_171),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_59),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_226),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_335),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_243),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_45),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_88),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_103),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_276),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_293),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_74),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_170),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_198),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_55),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_366),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_60),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_124),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_362),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_216),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_280),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_26),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_141),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_206),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_289),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_186),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_101),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_256),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_372),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_125),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_285),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_368),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_365),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_248),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_96),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_59),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_53),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_173),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_263),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_189),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_336),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_363),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_30),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_24),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_238),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_129),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_14),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_87),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_314),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_3),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_203),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_94),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_277),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_272),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_31),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_0),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g539 ( 
.A(n_33),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_138),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_230),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_234),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_98),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_155),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_109),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_539),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_448),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_460),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_460),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_448),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_457),
.B(n_476),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_532),
.Y(n_553)
);

OAI22x1_ASAP7_75t_SL g554 ( 
.A1(n_383),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_475),
.B(n_1),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_532),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_485),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_391),
.B(n_2),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_483),
.B(n_5),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_488),
.B(n_5),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_491),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_532),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_467),
.B(n_6),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_394),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_520),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_478),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_542),
.Y(n_569)
);

OAI22x1_ASAP7_75t_R g570 ( 
.A1(n_453),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_403),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_478),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_478),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_410),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_478),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_416),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_513),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_462),
.B(n_7),
.Y(n_579)
);

AOI22x1_ASAP7_75t_SL g580 ( 
.A1(n_480),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_475),
.A2(n_91),
.B(n_90),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_513),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_378),
.B(n_10),
.Y(n_583)
);

BUFx12f_ASAP7_75t_L g584 ( 
.A(n_542),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_418),
.B(n_12),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_513),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_399),
.B(n_13),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_380),
.A2(n_13),
.B(n_14),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_426),
.B(n_15),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_389),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_423),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_382),
.Y(n_593)
);

BUFx12f_ASAP7_75t_L g594 ( 
.A(n_419),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_446),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_525),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_447),
.B(n_386),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_456),
.Y(n_598)
);

INVx6_ASAP7_75t_L g599 ( 
.A(n_433),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_425),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_463),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_433),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_468),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_433),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_404),
.B(n_16),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_526),
.B(n_17),
.Y(n_607)
);

BUFx12f_ASAP7_75t_L g608 ( 
.A(n_427),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_502),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_497),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_388),
.B(n_397),
.Y(n_611)
);

BUFx8_ASAP7_75t_SL g612 ( 
.A(n_393),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_424),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_517),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_412),
.B(n_18),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_384),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_612),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_612),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_602),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_599),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_599),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_600),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_553),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_600),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_556),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_584),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_547),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_613),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_590),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_594),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_547),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_608),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_567),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_563),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_567),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_569),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_569),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_602),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_555),
.B(n_422),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_558),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_546),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_548),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_562),
.B(n_454),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_546),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_562),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_552),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_604),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_551),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_604),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_R g651 ( 
.A(n_579),
.B(n_396),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_551),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_605),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_595),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_606),
.B(n_434),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_555),
.B(n_516),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_605),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_552),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_549),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_597),
.B(n_458),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_605),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_613),
.Y(n_662)
);

CKINVDCx16_ASAP7_75t_R g663 ( 
.A(n_615),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_616),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_593),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_616),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_640),
.B(n_559),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_639),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_640),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_643),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_623),
.B(n_461),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_656),
.A2(n_581),
.B(n_564),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_659),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_659),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_644),
.B(n_609),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_629),
.B(n_583),
.C(n_561),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_647),
.B(n_583),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_625),
.Y(n_679)
);

OAI21xp33_ASAP7_75t_L g680 ( 
.A1(n_629),
.A2(n_561),
.B(n_587),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_665),
.B(n_589),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_654),
.Y(n_682)
);

INVxp67_ASAP7_75t_SL g683 ( 
.A(n_660),
.Y(n_683)
);

BUFx6f_ASAP7_75t_SL g684 ( 
.A(n_662),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_650),
.B(n_614),
.Y(n_685)
);

NOR2x1p5_ASAP7_75t_L g686 ( 
.A(n_642),
.B(n_424),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_646),
.B(n_589),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_653),
.B(n_614),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_648),
.Y(n_689)
);

AND2x2_ASAP7_75t_SL g690 ( 
.A(n_663),
.B(n_588),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_634),
.B(n_587),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_659),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_636),
.B(n_585),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_664),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_657),
.B(n_550),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_651),
.B(n_528),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_658),
.B(n_585),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_661),
.B(n_550),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_637),
.A2(n_464),
.B1(n_560),
.B2(n_459),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_666),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_624),
.B(n_550),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_621),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_658),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_654),
.B(n_597),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_593),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_626),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_622),
.Y(n_707)
);

INVxp33_ASAP7_75t_L g708 ( 
.A(n_655),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_635),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_645),
.B(n_617),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_655),
.B(n_379),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_649),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_630),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_631),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_633),
.B(n_550),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_627),
.B(n_611),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_628),
.B(n_565),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_652),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_632),
.B(n_565),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_641),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_618),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_619),
.B(n_611),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_640),
.B(n_381),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_639),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_640),
.B(n_565),
.Y(n_725)
);

INVx5_ASAP7_75t_L g726 ( 
.A(n_659),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_640),
.B(n_409),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_640),
.B(n_466),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_640),
.B(n_387),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_640),
.B(n_565),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_709),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_668),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_SL g733 ( 
.A1(n_727),
.A2(n_489),
.B1(n_570),
.B2(n_537),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_706),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_720),
.A2(n_596),
.B1(n_518),
.B2(n_489),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_674),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_706),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_667),
.A2(n_385),
.B(n_607),
.C(n_401),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_724),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_703),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_675),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_R g742 ( 
.A(n_721),
.B(n_390),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_728),
.B(n_683),
.Y(n_743)
);

BUFx8_ASAP7_75t_L g744 ( 
.A(n_684),
.Y(n_744)
);

NOR2xp67_ASAP7_75t_L g745 ( 
.A(n_669),
.B(n_595),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_677),
.A2(n_523),
.B1(n_545),
.B2(n_492),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_699),
.A2(n_596),
.B1(n_607),
.B2(n_402),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_683),
.B(n_392),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_712),
.Y(n_749)
);

INVx5_ASAP7_75t_L g750 ( 
.A(n_704),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_718),
.B(n_610),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_687),
.B(n_437),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_700),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_671),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_679),
.Y(n_755)
);

BUFx8_ASAP7_75t_L g756 ( 
.A(n_684),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_710),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_725),
.B(n_414),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_702),
.B(n_566),
.Y(n_759)
);

NOR2x1p5_ASAP7_75t_L g760 ( 
.A(n_713),
.B(n_441),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_677),
.B(n_395),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_691),
.B(n_398),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_682),
.B(n_708),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_693),
.B(n_400),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_689),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_682),
.B(n_572),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_730),
.B(n_417),
.Y(n_767)
);

AND3x1_ASAP7_75t_L g768 ( 
.A(n_680),
.B(n_554),
.C(n_580),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_678),
.A2(n_406),
.B1(n_407),
.B2(n_405),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_670),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_694),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_707),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_692),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_712),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_705),
.B(n_408),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_686),
.B(n_575),
.Y(n_776)
);

AND2x6_ASAP7_75t_SL g777 ( 
.A(n_722),
.B(n_577),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_717),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_690),
.A2(n_588),
.B1(n_509),
.B2(n_500),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_697),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_673),
.A2(n_429),
.B(n_420),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_690),
.B(n_436),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_723),
.A2(n_413),
.B1(n_415),
.B2(n_411),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_697),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_676),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_719),
.Y(n_786)
);

INVxp33_ASAP7_75t_L g787 ( 
.A(n_716),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_714),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_729),
.A2(n_440),
.B1(n_445),
.B2(n_439),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_685),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_688),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_711),
.B(n_455),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_696),
.B(n_479),
.Y(n_793)
);

CKINVDCx8_ASAP7_75t_R g794 ( 
.A(n_716),
.Y(n_794)
);

BUFx8_ASAP7_75t_SL g795 ( 
.A(n_715),
.Y(n_795)
);

INVx5_ASAP7_75t_L g796 ( 
.A(n_726),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_701),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_672),
.B(n_421),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_695),
.A2(n_472),
.B1(n_474),
.B2(n_470),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_698),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_726),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_670),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_667),
.B(n_477),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_667),
.B(n_493),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_681),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_667),
.B(n_501),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_709),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_702),
.B(n_592),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_667),
.A2(n_601),
.B(n_603),
.C(n_598),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_709),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_703),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_R g812 ( 
.A(n_721),
.B(n_428),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_674),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_679),
.Y(n_814)
);

BUFx4f_ASAP7_75t_L g815 ( 
.A(n_713),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_667),
.B(n_505),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_709),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_667),
.B(n_508),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_679),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_709),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_709),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_681),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_709),
.Y(n_823)
);

BUFx4f_ASAP7_75t_SL g824 ( 
.A(n_670),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_727),
.A2(n_431),
.B1(n_432),
.B2(n_430),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_677),
.A2(n_531),
.B1(n_540),
.B2(n_533),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_709),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_727),
.B(n_490),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_SL g829 ( 
.A(n_742),
.B(n_435),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_781),
.A2(n_582),
.B(n_576),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_743),
.A2(n_442),
.B1(n_443),
.B2(n_438),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_749),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_753),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_734),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_779),
.A2(n_582),
.B(n_576),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_770),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_SL g837 ( 
.A(n_746),
.B(n_499),
.C(n_494),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_750),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_737),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_822),
.B(n_757),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_748),
.A2(n_800),
.B(n_790),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_752),
.B(n_449),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_SL g843 ( 
.A(n_787),
.B(n_519),
.C(n_504),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_763),
.B(n_529),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_803),
.B(n_450),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_804),
.B(n_451),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_744),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_791),
.A2(n_557),
.B(n_549),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_774),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_824),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_785),
.A2(n_782),
.B(n_767),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_758),
.A2(n_557),
.B(n_549),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_731),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_814),
.B(n_517),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_806),
.B(n_452),
.Y(n_855)
);

BUFx12f_ASAP7_75t_L g856 ( 
.A(n_744),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_802),
.Y(n_857)
);

INVx6_ASAP7_75t_L g858 ( 
.A(n_756),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_816),
.B(n_818),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_776),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_810),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_772),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_780),
.B(n_465),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_761),
.A2(n_571),
.B(n_471),
.C(n_473),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_784),
.B(n_469),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_750),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_745),
.B(n_571),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_793),
.A2(n_482),
.B1(n_484),
.B2(n_481),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_766),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_740),
.B(n_530),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_794),
.B(n_538),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_738),
.A2(n_487),
.B(n_495),
.C(n_486),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_826),
.A2(n_498),
.B(n_503),
.C(n_496),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_786),
.B(n_762),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_817),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_759),
.B(n_92),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_SL g877 ( 
.A1(n_768),
.A2(n_507),
.B1(n_510),
.B2(n_506),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_SL g878 ( 
.A(n_819),
.B(n_511),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_776),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_755),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_821),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_792),
.A2(n_823),
.B1(n_827),
.B2(n_820),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_797),
.B(n_512),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_751),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_778),
.B(n_514),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_812),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_759),
.B(n_95),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_795),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_796),
.A2(n_573),
.B(n_568),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_751),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_825),
.B(n_732),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_809),
.A2(n_521),
.B(n_522),
.C(n_515),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_739),
.B(n_524),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_775),
.B(n_527),
.Y(n_894)
);

NAND2xp33_ASAP7_75t_SL g895 ( 
.A(n_760),
.B(n_534),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_815),
.B(n_535),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_788),
.B(n_536),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_811),
.B(n_541),
.Y(n_898)
);

BUFx12f_ASAP7_75t_L g899 ( 
.A(n_756),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_754),
.B(n_543),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_808),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_SL g902 ( 
.A1(n_764),
.A2(n_544),
.B(n_20),
.C(n_18),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_796),
.A2(n_574),
.B(n_573),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_765),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_736),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_798),
.B(n_19),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_789),
.A2(n_616),
.B(n_578),
.C(n_586),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_769),
.B(n_574),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_771),
.B(n_574),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_808),
.B(n_99),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_736),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_799),
.A2(n_22),
.B(n_19),
.C(n_21),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_733),
.B(n_22),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_SL g914 ( 
.A(n_735),
.B(n_23),
.C(n_24),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_783),
.B(n_591),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_741),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_741),
.A2(n_105),
.B1(n_106),
.B2(n_104),
.Y(n_917)
);

INVx6_ASAP7_75t_L g918 ( 
.A(n_777),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_741),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_SL g920 ( 
.A(n_773),
.B(n_27),
.C(n_28),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_813),
.Y(n_921)
);

OR2x4_ASAP7_75t_L g922 ( 
.A(n_801),
.B(n_29),
.Y(n_922)
);

AOI21xp33_ASAP7_75t_L g923 ( 
.A1(n_801),
.A2(n_30),
.B(n_31),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_805),
.B(n_32),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_750),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_743),
.A2(n_110),
.B1(n_111),
.B2(n_107),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_743),
.B(n_32),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_743),
.B(n_33),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_753),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_781),
.A2(n_113),
.B(n_112),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_743),
.Y(n_931)
);

BUFx12f_ASAP7_75t_L g932 ( 
.A(n_744),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_770),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_805),
.B(n_34),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_753),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_L g936 ( 
.A1(n_828),
.A2(n_34),
.B(n_36),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_R g937 ( 
.A(n_755),
.B(n_116),
.Y(n_937)
);

OAI22x1_ASAP7_75t_L g938 ( 
.A1(n_805),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_743),
.B(n_38),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_781),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_782),
.A2(n_43),
.B(n_40),
.C(n_42),
.Y(n_941)
);

AO21x1_ASAP7_75t_L g942 ( 
.A1(n_781),
.A2(n_42),
.B(n_43),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_781),
.A2(n_119),
.B(n_117),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_743),
.A2(n_121),
.B1(n_122),
.B2(n_120),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_770),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_807),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_781),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_750),
.B(n_123),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_749),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_782),
.A2(n_49),
.B(n_46),
.C(n_47),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_781),
.A2(n_127),
.B(n_126),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_753),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_807),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_743),
.B(n_47),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_781),
.A2(n_130),
.B(n_128),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_805),
.B(n_49),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_805),
.B(n_50),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_749),
.Y(n_958)
);

BUFx12f_ASAP7_75t_L g959 ( 
.A(n_744),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_743),
.B(n_50),
.Y(n_960)
);

NAND2x1p5_ASAP7_75t_L g961 ( 
.A(n_750),
.B(n_131),
.Y(n_961)
);

AOI221xp5_ASAP7_75t_L g962 ( 
.A1(n_747),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.C(n_55),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_743),
.B(n_51),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_743),
.B(n_56),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_828),
.A2(n_133),
.B1(n_135),
.B2(n_132),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_743),
.B(n_56),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_805),
.B(n_57),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_840),
.B(n_58),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_836),
.B(n_58),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_906),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_857),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_933),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_850),
.Y(n_973)
);

BUFx6f_ASAP7_75t_SL g974 ( 
.A(n_880),
.Y(n_974)
);

NOR2x1_ASAP7_75t_R g975 ( 
.A(n_847),
.B(n_856),
.Y(n_975)
);

INVx8_ASAP7_75t_L g976 ( 
.A(n_876),
.Y(n_976)
);

AOI22x1_ASAP7_75t_L g977 ( 
.A1(n_851),
.A2(n_841),
.B1(n_931),
.B2(n_930),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_945),
.Y(n_978)
);

BUFx24_ASAP7_75t_L g979 ( 
.A(n_876),
.Y(n_979)
);

NOR2xp67_ASAP7_75t_L g980 ( 
.A(n_886),
.B(n_137),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_860),
.B(n_879),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_859),
.A2(n_140),
.B(n_139),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_862),
.B(n_142),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_832),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_849),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_833),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_905),
.Y(n_987)
);

BUFx8_ASAP7_75t_L g988 ( 
.A(n_899),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_862),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_905),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_949),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_862),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_929),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_949),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_935),
.Y(n_995)
);

INVx6_ASAP7_75t_L g996 ( 
.A(n_858),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_869),
.B(n_63),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_916),
.Y(n_998)
);

AO21x2_ASAP7_75t_L g999 ( 
.A1(n_943),
.A2(n_151),
.B(n_150),
.Y(n_999)
);

OAI21x1_ASAP7_75t_SL g1000 ( 
.A1(n_942),
.A2(n_154),
.B(n_152),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_842),
.B(n_63),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_951),
.A2(n_157),
.B(n_156),
.Y(n_1002)
);

BUFx2_ASAP7_75t_R g1003 ( 
.A(n_888),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_901),
.B(n_158),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_927),
.B(n_64),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_884),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_844),
.B(n_64),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_834),
.B(n_162),
.Y(n_1008)
);

AOI22x1_ASAP7_75t_L g1009 ( 
.A1(n_955),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_838),
.B(n_168),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_867),
.B(n_65),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_830),
.A2(n_172),
.B(n_169),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_925),
.B(n_174),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_958),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_839),
.B(n_887),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_932),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_875),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_887),
.B(n_910),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_952),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_881),
.Y(n_1020)
);

INVx8_ASAP7_75t_L g1021 ( 
.A(n_910),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_904),
.Y(n_1022)
);

AOI22x1_ASAP7_75t_L g1023 ( 
.A1(n_938),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_835),
.A2(n_177),
.B(n_175),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_921),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_853),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_928),
.A2(n_180),
.B(n_179),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_909),
.A2(n_184),
.B(n_181),
.Y(n_1028)
);

BUFx2_ASAP7_75t_SL g1029 ( 
.A(n_925),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_911),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_861),
.Y(n_1031)
);

AO21x2_ASAP7_75t_L g1032 ( 
.A1(n_939),
.A2(n_187),
.B(n_185),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_890),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_946),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_922),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_954),
.A2(n_194),
.B(n_193),
.Y(n_1036)
);

OA21x2_ASAP7_75t_L g1037 ( 
.A1(n_960),
.A2(n_199),
.B(n_196),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_858),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_963),
.A2(n_202),
.B(n_200),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_870),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_953),
.Y(n_1041)
);

OR3x4_ASAP7_75t_SL g1042 ( 
.A(n_914),
.B(n_918),
.C(n_962),
.Y(n_1042)
);

AOI22x1_ASAP7_75t_L g1043 ( 
.A1(n_848),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_866),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_864),
.A2(n_205),
.B(n_204),
.Y(n_1045)
);

AO21x1_ASAP7_75t_L g1046 ( 
.A1(n_964),
.A2(n_69),
.B(n_70),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_911),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_966),
.B(n_71),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_882),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_959),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_924),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_891),
.A2(n_211),
.B(n_210),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_854),
.Y(n_1053)
);

AO21x2_ASAP7_75t_L g1054 ( 
.A1(n_872),
.A2(n_214),
.B(n_213),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_898),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_961),
.Y(n_1056)
);

AO21x2_ASAP7_75t_L g1057 ( 
.A1(n_894),
.A2(n_217),
.B(n_215),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_871),
.B(n_72),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_915),
.A2(n_219),
.B(n_218),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_948),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_893),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_845),
.B(n_846),
.Y(n_1062)
);

AO21x1_ASAP7_75t_L g1063 ( 
.A1(n_926),
.A2(n_73),
.B(n_74),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_919),
.A2(n_221),
.B(n_220),
.Y(n_1064)
);

AO21x1_ASAP7_75t_L g1065 ( 
.A1(n_944),
.A2(n_73),
.B(n_75),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_918),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_934),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_900),
.Y(n_1068)
);

BUFx2_ASAP7_75t_SL g1069 ( 
.A(n_917),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_913),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_863),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_937),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_883),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_865),
.Y(n_1074)
);

AOI22x1_ASAP7_75t_L g1075 ( 
.A1(n_852),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_837),
.A2(n_897),
.B1(n_843),
.B2(n_885),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_940),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_855),
.A2(n_225),
.B(n_224),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_947),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_936),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_956),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_L g1082 ( 
.A(n_854),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_957),
.B(n_76),
.Y(n_1083)
);

INVx5_ASAP7_75t_SL g1084 ( 
.A(n_878),
.Y(n_1084)
);

BUFx2_ASAP7_75t_R g1085 ( 
.A(n_874),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_941),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_829),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_967),
.B(n_77),
.Y(n_1088)
);

OA21x2_ASAP7_75t_L g1089 ( 
.A1(n_892),
.A2(n_228),
.B(n_227),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_920),
.Y(n_1090)
);

AO21x1_ASAP7_75t_SL g1091 ( 
.A1(n_965),
.A2(n_923),
.B(n_868),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_908),
.Y(n_1092)
);

INVx3_ASAP7_75t_SL g1093 ( 
.A(n_896),
.Y(n_1093)
);

BUFx12f_ASAP7_75t_L g1094 ( 
.A(n_895),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_877),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_831),
.B(n_231),
.Y(n_1096)
);

INVx8_ASAP7_75t_L g1097 ( 
.A(n_902),
.Y(n_1097)
);

BUFx2_ASAP7_75t_R g1098 ( 
.A(n_950),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_912),
.B(n_78),
.C(n_79),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_873),
.A2(n_233),
.B(n_232),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_907),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_889),
.Y(n_1102)
);

AO21x2_ASAP7_75t_L g1103 ( 
.A1(n_903),
.A2(n_236),
.B(n_235),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_850),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1070),
.B(n_78),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1022),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_992),
.Y(n_1107)
);

BUFx2_ASAP7_75t_R g1108 ( 
.A(n_1016),
.Y(n_1108)
);

BUFx10_ASAP7_75t_L g1109 ( 
.A(n_996),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_986),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_1038),
.B(n_237),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_993),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_1066),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_1014),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_995),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_972),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_978),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1019),
.Y(n_1118)
);

BUFx2_ASAP7_75t_R g1119 ( 
.A(n_1050),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1026),
.Y(n_1120)
);

CKINVDCx14_ASAP7_75t_R g1121 ( 
.A(n_991),
.Y(n_1121)
);

AO21x1_ASAP7_75t_L g1122 ( 
.A1(n_1001),
.A2(n_79),
.B(n_80),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_1038),
.B(n_1025),
.Y(n_1123)
);

CKINVDCx11_ASAP7_75t_R g1124 ( 
.A(n_994),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1030),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1058),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1005),
.A2(n_1048),
.B(n_1012),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1031),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1034),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1007),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_971),
.Y(n_1131)
);

INVx6_ASAP7_75t_L g1132 ( 
.A(n_1038),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1067),
.B(n_86),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_973),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_988),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1083),
.A2(n_89),
.B1(n_239),
.B2(n_240),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1081),
.B(n_89),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1051),
.B(n_241),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_1025),
.B(n_989),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1104),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1017),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1088),
.A2(n_242),
.B1(n_246),
.B2(n_249),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_976),
.B(n_252),
.Y(n_1143)
);

CKINVDCx6p67_ASAP7_75t_R g1144 ( 
.A(n_979),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1077),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_984),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1084),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_985),
.Y(n_1148)
);

BUFx2_ASAP7_75t_R g1149 ( 
.A(n_1095),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_992),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1079),
.Y(n_1151)
);

AO21x1_ASAP7_75t_L g1152 ( 
.A1(n_1027),
.A2(n_258),
.B(n_259),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_SL g1153 ( 
.A1(n_982),
.A2(n_260),
.B(n_261),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1020),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_968),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1071),
.B(n_266),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1018),
.B(n_376),
.Y(n_1157)
);

CKINVDCx6p67_ASAP7_75t_R g1158 ( 
.A(n_974),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1030),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_989),
.B(n_267),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1074),
.B(n_268),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1041),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1076),
.A2(n_270),
.B1(n_271),
.B2(n_274),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_992),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_SL g1165 ( 
.A(n_1003),
.B(n_275),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1049),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_1033),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_SL g1168 ( 
.A1(n_1000),
.A2(n_281),
.B(n_282),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1040),
.B(n_283),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_988),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1011),
.B(n_997),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_1084),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1006),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1055),
.A2(n_290),
.B1(n_292),
.B2(n_295),
.Y(n_1174)
);

AOI222xp33_ASAP7_75t_L g1175 ( 
.A1(n_970),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.C1(n_299),
.C2(n_300),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1101),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1047),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1080),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_1087),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1090),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1072),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1091),
.A2(n_305),
.B1(n_308),
.B2(n_309),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1068),
.B(n_310),
.Y(n_1183)
);

OAI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1073),
.A2(n_1062),
.B1(n_1093),
.B2(n_1061),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1015),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_987),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1091),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1044),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1035),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_998),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1099),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1086),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_976),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1069),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_990),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1094),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1069),
.A2(n_324),
.B1(n_325),
.B2(n_329),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_981),
.B(n_1056),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1063),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1021),
.A2(n_1053),
.B1(n_1023),
.B2(n_1082),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1004),
.B(n_333),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1008),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1092),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1059),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_969),
.A2(n_338),
.B1(n_340),
.B2(n_343),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1056),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_981),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1146),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_SL g1209 ( 
.A1(n_1183),
.A2(n_983),
.B(n_1039),
.C(n_1078),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1204),
.A2(n_1065),
.A3(n_1046),
.B(n_1064),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1166),
.B(n_1060),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1109),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1171),
.B(n_1085),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_1113),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1132),
.B(n_1029),
.Y(n_1215)
);

AOI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_1130),
.A2(n_1097),
.B1(n_1042),
.B2(n_1053),
.C(n_1060),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1170),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_R g1218 ( 
.A(n_1181),
.B(n_1056),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1184),
.A2(n_1096),
.B(n_977),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1148),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1106),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1132),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1133),
.B(n_980),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_R g1224 ( 
.A(n_1179),
.B(n_1102),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1137),
.B(n_1098),
.Y(n_1225)
);

INVxp33_ASAP7_75t_SL g1226 ( 
.A(n_1131),
.Y(n_1226)
);

INVx5_ASAP7_75t_SL g1227 ( 
.A(n_1144),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1116),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1112),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1188),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1110),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_SL g1233 ( 
.A(n_1200),
.B(n_975),
.C(n_1009),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_R g1234 ( 
.A(n_1121),
.B(n_1097),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1175),
.A2(n_1075),
.B1(n_1043),
.B2(n_1054),
.Y(n_1235)
);

BUFx4f_ASAP7_75t_SL g1236 ( 
.A(n_1158),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1105),
.B(n_1029),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1173),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1191),
.A2(n_1075),
.B1(n_1043),
.B2(n_1002),
.Y(n_1239)
);

NAND2xp33_ASAP7_75t_R g1240 ( 
.A(n_1117),
.B(n_1089),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1134),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1115),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1167),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1201),
.B(n_1013),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1118),
.Y(n_1245)
);

XNOR2xp5_ASAP7_75t_L g1246 ( 
.A(n_1135),
.B(n_1010),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1120),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1136),
.A2(n_1199),
.B1(n_1152),
.B2(n_1126),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1192),
.B(n_1202),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1122),
.A2(n_999),
.B1(n_1100),
.B2(n_1089),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1138),
.B(n_1032),
.Y(n_1251)
);

INVx3_ASAP7_75t_SL g1252 ( 
.A(n_1140),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1114),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1108),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_1165),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1193),
.B(n_1024),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1128),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1123),
.B(n_1052),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1206),
.B(n_1045),
.Y(n_1259)
);

NOR2x1p5_ASAP7_75t_L g1260 ( 
.A(n_1196),
.B(n_1057),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1207),
.B(n_1036),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_R g1262 ( 
.A(n_1125),
.B(n_344),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1189),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_R g1264 ( 
.A(n_1124),
.B(n_1103),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1141),
.B(n_1037),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1149),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1203),
.B(n_1028),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1129),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1206),
.B(n_345),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1178),
.B(n_373),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1154),
.B(n_347),
.Y(n_1271)
);

XOR2xp5_ASAP7_75t_L g1272 ( 
.A(n_1119),
.B(n_348),
.Y(n_1272)
);

NOR3xp33_ASAP7_75t_SL g1273 ( 
.A(n_1156),
.B(n_351),
.C(n_352),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1164),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_R g1275 ( 
.A(n_1159),
.B(n_1177),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1107),
.Y(n_1276)
);

CKINVDCx16_ASAP7_75t_R g1277 ( 
.A(n_1143),
.Y(n_1277)
);

NOR3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1161),
.B(n_356),
.C(n_357),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1163),
.A2(n_358),
.B1(n_360),
.B2(n_361),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1107),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1159),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1230),
.B(n_1154),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1229),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1222),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1242),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1221),
.Y(n_1286)
);

OAI211xp5_ASAP7_75t_L g1287 ( 
.A1(n_1248),
.A2(n_1205),
.B(n_1182),
.C(n_1187),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1268),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1208),
.B(n_1162),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1245),
.B(n_1151),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1247),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1257),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1249),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1219),
.B(n_1153),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1220),
.B(n_1243),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1215),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1265),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1232),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1259),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1228),
.B(n_1162),
.Y(n_1300)
);

AOI221xp5_ASAP7_75t_L g1301 ( 
.A1(n_1235),
.A2(n_1155),
.B1(n_1142),
.B2(n_1180),
.C(n_1168),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1237),
.B(n_1195),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1267),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1275),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1251),
.B(n_1145),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1216),
.A2(n_1147),
.B1(n_1172),
.B2(n_1174),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1253),
.B(n_1169),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1280),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1211),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1240),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1225),
.A2(n_1279),
.B1(n_1239),
.B2(n_1255),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1226),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1210),
.B(n_1176),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1258),
.B(n_1260),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1218),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1223),
.B(n_1190),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1244),
.B(n_1186),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1213),
.B(n_1198),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1256),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1261),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1231),
.B(n_1127),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1286),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1320),
.B(n_1277),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1299),
.B(n_1256),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1293),
.B(n_1270),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1317),
.B(n_1266),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1315),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1299),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1305),
.B(n_1274),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1283),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1320),
.B(n_1271),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1285),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1305),
.B(n_1250),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1299),
.B(n_1258),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1297),
.B(n_1303),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1302),
.B(n_1233),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1291),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1288),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1311),
.B(n_1278),
.C(n_1273),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1304),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1291),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1292),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1292),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1309),
.B(n_1281),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1311),
.B(n_1316),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1297),
.B(n_1263),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1290),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1296),
.B(n_1264),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1335),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1322),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1337),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1323),
.B(n_1303),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1345),
.B(n_1310),
.Y(n_1353)
);

NAND2xp33_ASAP7_75t_SL g1354 ( 
.A(n_1345),
.B(n_1262),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1333),
.B(n_1347),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1333),
.B(n_1313),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1330),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1337),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1332),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1342),
.B(n_1319),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1338),
.B(n_1321),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1342),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1331),
.B(n_1321),
.Y(n_1363)
);

OAI21xp33_ASAP7_75t_L g1364 ( 
.A1(n_1339),
.A2(n_1306),
.B(n_1287),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1343),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1329),
.B(n_1319),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1327),
.B(n_1319),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1343),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1340),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1349),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1364),
.B(n_1340),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1350),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1358),
.Y(n_1373)
);

OAI322xp33_ASAP7_75t_L g1374 ( 
.A1(n_1353),
.A2(n_1325),
.A3(n_1289),
.B1(n_1282),
.B2(n_1300),
.C1(n_1348),
.C2(n_1307),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1369),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1363),
.B(n_1346),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1351),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_1351),
.B(n_1328),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1357),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1353),
.A2(n_1294),
.B1(n_1348),
.B2(n_1314),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1365),
.Y(n_1381)
);

NOR2xp67_ASAP7_75t_R g1382 ( 
.A(n_1369),
.B(n_1328),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1361),
.B(n_1341),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1352),
.B(n_1312),
.Y(n_1384)
);

NAND2x1_ASAP7_75t_L g1385 ( 
.A(n_1362),
.B(n_1314),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1365),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1372),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1374),
.A2(n_1336),
.B(n_1294),
.C(n_1344),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1371),
.A2(n_1246),
.B(n_1272),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1380),
.A2(n_1301),
.B(n_1354),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1375),
.Y(n_1391)
);

NOR3xp33_ASAP7_75t_L g1392 ( 
.A(n_1374),
.B(n_1354),
.C(n_1295),
.Y(n_1392)
);

OAI21xp33_ASAP7_75t_L g1393 ( 
.A1(n_1370),
.A2(n_1356),
.B(n_1355),
.Y(n_1393)
);

AOI21xp33_ASAP7_75t_L g1394 ( 
.A1(n_1385),
.A2(n_1294),
.B(n_1314),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1389),
.B(n_1214),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1391),
.Y(n_1396)
);

OAI211xp5_ASAP7_75t_L g1397 ( 
.A1(n_1390),
.A2(n_1392),
.B(n_1388),
.C(n_1394),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1387),
.B(n_1355),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1393),
.B(n_1356),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1397),
.B(n_1379),
.Y(n_1400)
);

NOR3x1_ASAP7_75t_L g1401 ( 
.A(n_1396),
.B(n_1308),
.C(n_1382),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1395),
.A2(n_1252),
.B(n_1209),
.C(n_1241),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1399),
.A2(n_1334),
.B1(n_1367),
.B2(n_1324),
.Y(n_1403)
);

OAI322xp33_ASAP7_75t_L g1404 ( 
.A1(n_1398),
.A2(n_1384),
.A3(n_1359),
.B1(n_1383),
.B2(n_1376),
.C1(n_1368),
.C2(n_1377),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1397),
.B(n_1373),
.Y(n_1405)
);

AOI211x1_ASAP7_75t_L g1406 ( 
.A1(n_1405),
.A2(n_1382),
.B(n_1326),
.C(n_1366),
.Y(n_1406)
);

OR2x6_ASAP7_75t_L g1407 ( 
.A(n_1402),
.B(n_1212),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1400),
.B(n_1360),
.Y(n_1408)
);

NOR3xp33_ASAP7_75t_L g1409 ( 
.A(n_1408),
.B(n_1404),
.C(n_1254),
.Y(n_1409)
);

O2A1O1Ixp5_ASAP7_75t_L g1410 ( 
.A1(n_1406),
.A2(n_1401),
.B(n_1386),
.C(n_1381),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1410),
.Y(n_1411)
);

NAND4xp25_ASAP7_75t_L g1412 ( 
.A(n_1411),
.B(n_1409),
.C(n_1403),
.D(n_1238),
.Y(n_1412)
);

INVxp33_ASAP7_75t_L g1413 ( 
.A(n_1412),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1412),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1414),
.A2(n_1236),
.B1(n_1217),
.B2(n_1407),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1413),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1416),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1415),
.B(n_1378),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1417),
.A2(n_1227),
.B1(n_1284),
.B2(n_1222),
.Y(n_1419)
);

NAND5xp2_ASAP7_75t_L g1420 ( 
.A(n_1418),
.B(n_1111),
.C(n_1227),
.D(n_1139),
.E(n_1234),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1419),
.B(n_1222),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1420),
.A2(n_1269),
.B(n_1318),
.Y(n_1422)
);

AOI21xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1421),
.A2(n_1160),
.B(n_1269),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1422),
.A2(n_1150),
.B(n_1276),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1424),
.A2(n_1284),
.B1(n_1107),
.B2(n_1224),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1423),
.A2(n_1197),
.B(n_1194),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1425),
.B(n_1298),
.Y(n_1427)
);

AOI21xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1427),
.A2(n_1426),
.B(n_364),
.Y(n_1428)
);


endmodule