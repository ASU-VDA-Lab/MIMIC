module real_jpeg_4087_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_57;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_50;
wire n_33;
wire n_29;
wire n_55;
wire n_58;
wire n_10;
wire n_31;
wire n_9;
wire n_49;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_60;
wire n_44;
wire n_46;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_48;
wire n_27;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_1),
.A2(n_9),
.B(n_12),
.Y(n_8)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_2),
.B(n_7),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_5),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_15),
.Y(n_13)
);

NOR5xp2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_36),
.C(n_50),
.D(n_55),
.E(n_58),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_19),
.B1(n_32),
.B2(n_35),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_17),
.A2(n_32),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_31),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_25),
.A2(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_39),
.B(n_41),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_47),
.Y(n_57)
);

OR2x4_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);


endmodule