module fake_aes_4146_n_566 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_566);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_566;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_69), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_1), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_24), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_33), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_44), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_21), .Y(n_86) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_49), .B(n_58), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_31), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_65), .Y(n_90) );
NOR2xp67_ASAP7_75t_L g91 ( .A(n_63), .B(n_57), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_20), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_46), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_45), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_52), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_61), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_43), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_51), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_64), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_50), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_54), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_66), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_32), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_67), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_75), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_18), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_76), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_12), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_19), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_34), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_25), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_60), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_15), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_35), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_28), .Y(n_115) );
NAND2xp33_ASAP7_75t_R g116 ( .A(n_90), .B(n_29), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_115), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_97), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_80), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_90), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_80), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_97), .Y(n_124) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_94), .B(n_79), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_94), .B(n_0), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_115), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_111), .B(n_2), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_97), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_81), .B(n_2), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_83), .B(n_3), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_115), .B(n_30), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_101), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_89), .B(n_3), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_135), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_124), .Y(n_143) );
INVx1_ASAP7_75t_SL g144 ( .A(n_126), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_120), .B(n_95), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_126), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_135), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_138), .B(n_96), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_138), .B(n_110), .Y(n_149) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_125), .B(n_87), .Y(n_150) );
AO22x2_ASAP7_75t_L g151 ( .A1(n_121), .A2(n_114), .B1(n_102), .B2(n_84), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_119), .B(n_98), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_125), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_134), .Y(n_154) );
BUFx10_ASAP7_75t_L g155 ( .A(n_134), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_135), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_119), .B(n_99), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_124), .Y(n_160) );
INVx1_ASAP7_75t_SL g161 ( .A(n_121), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_122), .B(n_92), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
OR2x6_ASAP7_75t_L g164 ( .A(n_132), .B(n_106), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_125), .A2(n_108), .B1(n_109), .B2(n_106), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_157), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_161), .B(n_130), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_142), .B(n_130), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_157), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
OR2x6_ASAP7_75t_L g173 ( .A(n_164), .B(n_132), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_150), .A2(n_123), .B1(n_137), .B2(n_127), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_164), .Y(n_175) );
NAND3xp33_ASAP7_75t_SL g176 ( .A(n_167), .B(n_100), .C(n_105), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_150), .A2(n_167), .B1(n_164), .B2(n_153), .Y(n_177) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_150), .A2(n_113), .B1(n_133), .B2(n_85), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_148), .B(n_122), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_164), .B(n_136), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_144), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_151), .A2(n_116), .B1(n_136), .B2(n_137), .Y(n_183) );
NOR2x2_ASAP7_75t_L g184 ( .A(n_164), .B(n_139), .Y(n_184) );
OR2x2_ASAP7_75t_SL g185 ( .A(n_146), .B(n_113), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_149), .B(n_123), .Y(n_186) );
INVxp33_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_151), .A2(n_127), .B1(n_129), .B2(n_134), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_154), .Y(n_191) );
NOR2x1_ASAP7_75t_L g192 ( .A(n_145), .B(n_129), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_152), .B(n_134), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_151), .B(n_139), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_142), .B(n_101), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_142), .A2(n_165), .B(n_163), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_142), .B(n_104), .Y(n_197) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_163), .B(n_103), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_163), .B(n_118), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_140), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_155), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_160), .B(n_118), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_179), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_179), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_179), .Y(n_206) );
AOI22x1_ASAP7_75t_L g207 ( .A1(n_198), .A2(n_165), .B1(n_163), .B2(n_151), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_182), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_175), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_181), .B(n_159), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_188), .A2(n_183), .B(n_186), .C(n_180), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_202), .Y(n_212) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_173), .B(n_165), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_173), .A2(n_166), .B1(n_165), .B2(n_131), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_202), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_196), .A2(n_154), .B(n_166), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_173), .A2(n_154), .B1(n_155), .B2(n_85), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_173), .A2(n_155), .B1(n_86), .B2(n_88), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_175), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_181), .B(n_155), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_181), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_185), .B(n_131), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_201), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_193), .A2(n_147), .B(n_141), .Y(n_224) );
INVx5_ASAP7_75t_L g225 ( .A(n_199), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_189), .Y(n_227) );
AO32x2_ASAP7_75t_L g228 ( .A1(n_178), .A2(n_117), .A3(n_128), .B1(n_135), .B2(n_91), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_184), .Y(n_229) );
CKINVDCx14_ASAP7_75t_R g230 ( .A(n_176), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_169), .B(n_86), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g233 ( .A1(n_177), .A2(n_112), .B1(n_88), .B2(n_93), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_201), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_190), .A2(n_114), .B(n_103), .C(n_93), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_174), .B(n_102), .Y(n_238) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_211), .A2(n_194), .B(n_195), .Y(n_239) );
OAI21xp33_ASAP7_75t_SL g240 ( .A1(n_238), .A2(n_212), .B(n_215), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_233), .A2(n_187), .B1(n_169), .B2(n_170), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_237), .B(n_187), .Y(n_242) );
INVx3_ASAP7_75t_SL g243 ( .A(n_208), .Y(n_243) );
OAI21x1_ASAP7_75t_SL g244 ( .A1(n_207), .A2(n_87), .B(n_192), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_224), .A2(n_198), .B(n_197), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_224), .A2(n_195), .B(n_197), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_225), .Y(n_247) );
NOR2xp67_ASAP7_75t_L g248 ( .A(n_219), .B(n_170), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_216), .A2(n_141), .B(n_140), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_229), .B(n_199), .Y(n_250) );
AO31x2_ASAP7_75t_L g251 ( .A1(n_235), .A2(n_104), .A3(n_107), .B(n_141), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_216), .A2(n_147), .B(n_140), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_214), .A2(n_147), .B(n_104), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_214), .A2(n_107), .B(n_168), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_221), .A2(n_199), .B1(n_191), .B2(n_201), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_225), .B(n_191), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_210), .B(n_201), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_210), .B(n_135), .Y(n_258) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_238), .A2(n_91), .B(n_171), .Y(n_259) );
CKINVDCx6p67_ASAP7_75t_R g260 ( .A(n_225), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_226), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_227), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_205), .A2(n_171), .B(n_168), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_209), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_236), .A2(n_218), .B1(n_219), .B2(n_232), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_206), .A2(n_200), .B(n_158), .Y(n_267) );
OR2x6_ASAP7_75t_L g268 ( .A(n_265), .B(n_209), .Y(n_268) );
OAI21xp33_ASAP7_75t_L g269 ( .A1(n_240), .A2(n_232), .B(n_222), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_261), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_265), .A2(n_225), .B1(n_231), .B2(n_209), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_261), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_267), .Y(n_273) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_244), .A2(n_228), .B(n_217), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_240), .B(n_213), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_246), .A2(n_220), .B(n_230), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_254), .A2(n_220), .B(n_128), .C(n_117), .Y(n_277) );
OAI21xp5_ASAP7_75t_SL g278 ( .A1(n_241), .A2(n_234), .B(n_223), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_254), .A2(n_128), .B(n_117), .C(n_228), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_242), .B(n_228), .Y(n_280) );
OAI21xp5_ASAP7_75t_SL g281 ( .A1(n_243), .A2(n_234), .B(n_223), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_242), .B(n_234), .Y(n_282) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_244), .A2(n_200), .B(n_128), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_262), .A2(n_243), .B1(n_258), .B2(n_250), .C(n_246), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_128), .B1(n_117), .B2(n_158), .C(n_223), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_260), .A2(n_128), .B1(n_117), .B2(n_158), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_258), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_260), .A2(n_158), .B1(n_5), .B2(n_6), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_250), .B(n_4), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_254), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_243), .A2(n_158), .B1(n_5), .B2(n_6), .C(n_7), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_270), .B(n_247), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_272), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_280), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_268), .B(n_247), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_273), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_287), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_268), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_290), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_284), .B(n_239), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_268), .B(n_259), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_273), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_283), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_279), .B(n_259), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_282), .B(n_259), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_269), .B(n_259), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
BUFx12f_ASAP7_75t_L g312 ( .A(n_278), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_274), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_297), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_294), .B(n_251), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_311), .A2(n_271), .B1(n_275), .B2(n_291), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_294), .B(n_251), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_297), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_298), .A2(n_289), .B1(n_276), .B2(n_288), .C(n_277), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_300), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_304), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_295), .B(n_251), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_312), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_304), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_295), .B(n_251), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_305), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_300), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_309), .B(n_251), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_309), .B(n_251), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_298), .B(n_274), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_308), .B(n_277), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_313), .Y(n_339) );
OR2x6_ASAP7_75t_L g340 ( .A(n_312), .B(n_253), .Y(n_340) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_313), .B(n_285), .C(n_286), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_313), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_311), .B(n_239), .Y(n_343) );
OAI33xp33_ASAP7_75t_L g344 ( .A1(n_302), .A2(n_266), .A3(n_7), .B1(n_8), .B2(n_9), .B3(n_10), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_239), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_337), .B(n_303), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_339), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_337), .B(n_345), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_345), .B(n_303), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_339), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_338), .B(n_301), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_338), .B(n_303), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_328), .B(n_302), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_336), .B(n_308), .Y(n_354) );
OAI33xp33_ASAP7_75t_L g355 ( .A1(n_327), .A2(n_301), .A3(n_296), .B1(n_305), .B2(n_306), .B3(n_266), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_336), .B(n_310), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_342), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_318), .B(n_310), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_318), .B(n_310), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_323), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_342), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_315), .B(n_296), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_319), .A2(n_322), .B(n_343), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_323), .Y(n_365) );
BUFx2_ASAP7_75t_SL g366 ( .A(n_326), .Y(n_366) );
AND2x4_ASAP7_75t_SL g367 ( .A(n_326), .B(n_299), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_334), .B(n_299), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_316), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_333), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_320), .B(n_299), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_320), .B(n_299), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_325), .B(n_307), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_333), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_317), .Y(n_375) );
AOI33xp33_ASAP7_75t_L g376 ( .A1(n_325), .A2(n_305), .A3(n_306), .B1(n_9), .B2(n_10), .B3(n_11), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_344), .A2(n_307), .B1(n_312), .B2(n_314), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_324), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_340), .A2(n_306), .B(n_314), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_324), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_329), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_334), .B(n_307), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_329), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_335), .B(n_253), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_335), .B(n_253), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_321), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_330), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_330), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_321), .B(n_249), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_332), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_391), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_348), .B(n_326), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_360), .B(n_326), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_349), .B(n_356), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_332), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_364), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_363), .B(n_331), .Y(n_399) );
NAND4xp75_ASAP7_75t_SL g400 ( .A(n_366), .B(n_340), .C(n_248), .D(n_260), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_349), .B(n_331), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_351), .B(n_340), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_340), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
INVxp33_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_367), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_351), .B(n_388), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_388), .B(n_340), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_378), .B(n_341), .C(n_248), .D(n_255), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_358), .B(n_252), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_376), .B(n_341), .C(n_158), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_366), .B(n_346), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_358), .B(n_249), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_389), .B(n_4), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_359), .B(n_249), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_389), .B(n_8), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_359), .B(n_252), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_367), .A2(n_264), .B1(n_239), .B2(n_256), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_370), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_354), .B(n_252), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_375), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_354), .B(n_11), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_391), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_368), .B(n_12), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_346), .B(n_13), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_373), .B(n_13), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_391), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_352), .B(n_14), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_352), .B(n_14), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_379), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_385), .B(n_15), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_365), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_385), .B(n_16), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_379), .Y(n_439) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_353), .B(n_16), .C(n_17), .D(n_18), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_381), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_367), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_347), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_371), .B(n_17), .Y(n_444) );
NAND4xp25_ASAP7_75t_SL g445 ( .A(n_380), .B(n_19), .C(n_20), .D(n_257), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_395), .A2(n_374), .B(n_386), .C(n_383), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_409), .B(n_394), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_405), .A2(n_372), .B(n_368), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_399), .B(n_383), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_421), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_440), .A2(n_355), .B1(n_381), .B2(n_382), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_396), .B(n_382), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_395), .A2(n_426), .B1(n_418), .B2(n_416), .Y(n_454) );
AOI322xp5_ASAP7_75t_L g455 ( .A1(n_427), .A2(n_350), .A3(n_347), .B1(n_361), .B2(n_357), .C1(n_384), .C2(n_387), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_396), .B(n_384), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_443), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_401), .B(n_386), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_424), .B(n_361), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_443), .Y(n_460) );
OAI32xp33_ASAP7_75t_L g461 ( .A1(n_405), .A2(n_357), .A3(n_350), .B1(n_390), .B2(n_264), .Y(n_461) );
OAI211xp5_ASAP7_75t_L g462 ( .A1(n_427), .A2(n_390), .B(n_264), .C(n_257), .Y(n_462) );
XOR2x2_ASAP7_75t_L g463 ( .A(n_414), .B(n_22), .Y(n_463) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_403), .A2(n_264), .B(n_245), .Y(n_464) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_400), .B(n_256), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_424), .B(n_245), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_436), .B(n_245), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_397), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_445), .A2(n_256), .B1(n_263), .B2(n_267), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_397), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_406), .B(n_256), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_428), .A2(n_263), .B1(n_26), .B2(n_27), .C(n_36), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_404), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_407), .Y(n_475) );
AOI32xp33_ASAP7_75t_L g476 ( .A1(n_432), .A2(n_267), .A3(n_37), .B1(n_38), .B2(n_39), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_411), .B(n_23), .C(n_40), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_408), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_392), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_393), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g481 ( .A1(n_432), .A2(n_42), .B1(n_47), .B2(n_48), .C1(n_53), .C2(n_55), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_406), .A2(n_442), .B1(n_426), .B2(n_402), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_401), .B(n_56), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_434), .A2(n_59), .B1(n_62), .B2(n_68), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_438), .B(n_70), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_438), .B(n_71), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g489 ( .A(n_442), .B(n_72), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_444), .B(n_418), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_434), .B(n_73), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_451), .B(n_403), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_448), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_479), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_468), .B(n_419), .Y(n_496) );
OAI21xp5_ASAP7_75t_SL g497 ( .A1(n_481), .A2(n_420), .B(n_416), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_455), .B(n_437), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_457), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_447), .B(n_410), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_477), .B(n_413), .C(n_439), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_452), .B(n_441), .Y(n_503) );
AO22x2_ASAP7_75t_SL g504 ( .A1(n_463), .A2(n_435), .B1(n_433), .B2(n_431), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_470), .B(n_415), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_471), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_446), .B(n_402), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_474), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_475), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_478), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_454), .A2(n_417), .B1(n_419), .B2(n_412), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_482), .Y(n_512) );
AO22x2_ASAP7_75t_L g513 ( .A1(n_454), .A2(n_429), .B1(n_430), .B2(n_425), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_483), .B(n_430), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_481), .A2(n_412), .B(n_417), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_450), .B(n_415), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_453), .Y(n_517) );
OAI221xp5_ASAP7_75t_SL g518 ( .A1(n_484), .A2(n_422), .B1(n_392), .B2(n_425), .C(n_77), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_458), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_456), .B(n_422), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_480), .B(n_74), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_459), .B(n_78), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_513), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_495), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_512), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g526 ( .A1(n_503), .A2(n_490), .B(n_491), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_495), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_512), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_498), .B(n_449), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_493), .B(n_466), .Y(n_530) );
AO22x2_ASAP7_75t_L g531 ( .A1(n_497), .A2(n_494), .B1(n_492), .B2(n_508), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_513), .B(n_464), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_499), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_511), .A2(n_462), .B(n_489), .Y(n_534) );
OAI31xp33_ASAP7_75t_L g535 ( .A1(n_513), .A2(n_489), .A3(n_473), .B(n_485), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_521), .Y(n_536) );
AOI221xp5_ASAP7_75t_SL g537 ( .A1(n_515), .A2(n_461), .B1(n_488), .B2(n_487), .C(n_472), .Y(n_537) );
AOI211xp5_ASAP7_75t_L g538 ( .A1(n_518), .A2(n_467), .B(n_486), .C(n_469), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g539 ( .A1(n_514), .A2(n_476), .B(n_465), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_492), .A2(n_507), .B1(n_520), .B2(n_504), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_531), .A2(n_514), .B1(n_517), .B2(n_506), .C(n_509), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_533), .Y(n_542) );
INVxp67_ASAP7_75t_L g543 ( .A(n_529), .Y(n_543) );
AOI211xp5_ASAP7_75t_L g544 ( .A1(n_540), .A2(n_502), .B(n_504), .C(n_507), .Y(n_544) );
AOI211xp5_ASAP7_75t_SL g545 ( .A1(n_539), .A2(n_521), .B(n_522), .C(n_507), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_531), .A2(n_492), .B1(n_519), .B2(n_501), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_536), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_531), .A2(n_510), .B(n_516), .Y(n_548) );
OAI21x1_ASAP7_75t_SL g549 ( .A1(n_534), .A2(n_519), .B(n_500), .Y(n_549) );
AOI211xp5_ASAP7_75t_L g550 ( .A1(n_535), .A2(n_496), .B(n_505), .C(n_500), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_544), .B(n_523), .C(n_537), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_547), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_542), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_545), .B(n_527), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_546), .A2(n_523), .B1(n_532), .B2(n_526), .C(n_527), .Y(n_555) );
AND4x1_ASAP7_75t_L g556 ( .A(n_551), .B(n_550), .C(n_541), .D(n_548), .Y(n_556) );
OAI222xp33_ASAP7_75t_L g557 ( .A1(n_554), .A2(n_543), .B1(n_523), .B2(n_532), .C1(n_536), .C2(n_549), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_552), .B(n_543), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_558), .A2(n_552), .B1(n_555), .B2(n_553), .Y(n_559) );
XOR2xp5_ASAP7_75t_L g560 ( .A(n_556), .B(n_524), .Y(n_560) );
OAI22xp33_ASAP7_75t_SL g561 ( .A1(n_559), .A2(n_557), .B1(n_524), .B2(n_528), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_560), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_562), .A2(n_538), .B1(n_530), .B2(n_525), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_563), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_564), .B(n_561), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_565), .A2(n_496), .B(n_505), .Y(n_566) );
endmodule