module fake_jpeg_13631_n_648 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_60),
.B(n_69),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_65),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_71),
.B(n_84),
.Y(n_165)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_76),
.Y(n_212)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_77),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_80),
.Y(n_224)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_82),
.Y(n_193)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_87),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_37),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_88),
.B(n_92),
.Y(n_191)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_18),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_43),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_24),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_115),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_106),
.Y(n_221)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_20),
.B(n_17),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_117),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_118),
.B(n_131),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g156 ( 
.A(n_121),
.Y(n_156)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_29),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_26),
.C(n_58),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_29),
.Y(n_126)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_28),
.Y(n_128)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

BUFx2_ASAP7_75t_SL g177 ( 
.A(n_129),
.Y(n_177)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_28),
.Y(n_130)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_38),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_57),
.B1(n_40),
.B2(n_45),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_135),
.A2(n_136),
.B1(n_52),
.B2(n_3),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_40),
.B1(n_45),
.B2(n_37),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_69),
.B(n_20),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_137),
.B(n_160),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_185),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_88),
.B(n_33),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_154),
.B(n_196),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_92),
.B(n_26),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_158),
.B(n_210),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_97),
.B(n_39),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_39),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_162),
.B(n_167),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_108),
.B(n_59),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_108),
.B(n_59),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_176),
.B(n_182),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_77),
.B(n_35),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_80),
.B(n_35),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_184),
.B(n_204),
.Y(n_262)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_121),
.B(n_38),
.CON(n_185),
.SN(n_185)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_87),
.B(n_31),
.C(n_33),
.Y(n_196)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_87),
.B(n_31),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_1),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_113),
.A2(n_58),
.B1(n_53),
.B2(n_27),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_198),
.A2(n_218),
.B1(n_52),
.B2(n_3),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_64),
.B(n_53),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_203),
.B(n_209),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_117),
.B(n_51),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_61),
.A2(n_51),
.B1(n_48),
.B2(n_34),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_110),
.B1(n_105),
.B2(n_104),
.Y(n_229)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_64),
.B(n_0),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_65),
.B(n_48),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_65),
.B(n_34),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_0),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_129),
.B(n_27),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_214),
.B(n_11),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_124),
.A2(n_38),
.B1(n_52),
.B2(n_3),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_66),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_73),
.Y(n_220)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_76),
.Y(n_222)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_78),
.Y(n_225)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_226),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_120),
.B1(n_119),
.B2(n_111),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_227),
.A2(n_229),
.B1(n_263),
.B2(n_293),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_228),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_232),
.B(n_274),
.Y(n_319)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_233),
.Y(n_334)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_234),
.Y(n_345)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_102),
.B1(n_95),
.B2(n_90),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_238),
.A2(n_250),
.B1(n_256),
.B2(n_264),
.Y(n_314)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_239),
.A2(n_281),
.B(n_283),
.Y(n_338)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_240),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_241),
.Y(n_362)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_243),
.Y(n_360)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_244),
.Y(n_353)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_209),
.A2(n_86),
.B1(n_52),
.B2(n_4),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_247),
.A2(n_174),
.B(n_194),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_248),
.B(n_272),
.Y(n_355)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_175),
.Y(n_253)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_157),
.Y(n_257)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_140),
.Y(n_258)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_185),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_165),
.B(n_4),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_260),
.B(n_273),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_207),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_218),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_179),
.Y(n_265)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_218),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_139),
.Y(n_271)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_180),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_276),
.Y(n_324)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_278),
.Y(n_327)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_178),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_279),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_148),
.B(n_11),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_280),
.B(n_282),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_192),
.B(n_149),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_148),
.B(n_12),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_191),
.B(n_13),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_285),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_287),
.Y(n_359)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_133),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_288),
.B(n_289),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_203),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_156),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_290),
.Y(n_329)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_224),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_142),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_144),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_161),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_171),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_164),
.A2(n_134),
.B1(n_189),
.B2(n_170),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_297),
.A2(n_299),
.B1(n_300),
.B2(n_302),
.Y(n_342)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_155),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_143),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_177),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_138),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_210),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_304),
.Y(n_308)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_145),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_192),
.B(n_191),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_305),
.C(n_187),
.Y(n_354)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_150),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_141),
.B(n_213),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_231),
.A2(n_165),
.B(n_134),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_306),
.B(n_354),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_307),
.A2(n_339),
.B1(n_364),
.B2(n_291),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_231),
.A2(n_132),
.B(n_188),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_318),
.A2(n_323),
.B(n_253),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_242),
.B(n_136),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_250),
.A2(n_186),
.B1(n_195),
.B2(n_211),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_343),
.B1(n_350),
.B2(n_351),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_174),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_346),
.C(n_303),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_262),
.B(n_281),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_336),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_251),
.B(n_169),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_229),
.A2(n_135),
.B1(n_153),
.B2(n_163),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_241),
.B(n_199),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_358),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_292),
.A2(n_177),
.B1(n_186),
.B2(n_151),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_261),
.B(n_231),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_305),
.A2(n_139),
.B1(n_216),
.B2(n_151),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_305),
.A2(n_159),
.B1(n_212),
.B2(n_216),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_261),
.A2(n_153),
.B1(n_159),
.B2(n_212),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_357),
.A2(n_271),
.B1(n_278),
.B2(n_252),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_261),
.B(n_146),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_303),
.B(n_246),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_363),
.B(n_296),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_247),
.A2(n_293),
.B1(n_263),
.B2(n_237),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_367),
.B(n_365),
.Y(n_423)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_270),
.C(n_288),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_372),
.C(n_391),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_266),
.C(n_265),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_314),
.A2(n_269),
.B1(n_243),
.B2(n_295),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_373),
.A2(n_377),
.B1(n_393),
.B2(n_398),
.Y(n_437)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_314),
.A2(n_274),
.B1(n_275),
.B2(n_272),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_379),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_308),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_382),
.Y(n_424)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_344),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_361),
.B(n_302),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_383),
.A2(n_316),
.B1(n_312),
.B2(n_342),
.Y(n_434)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_384),
.B(n_385),
.Y(n_432)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_335),
.A2(n_240),
.B1(n_244),
.B2(n_228),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_388),
.B(n_389),
.Y(n_444)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_310),
.A2(n_249),
.B1(n_230),
.B2(n_255),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_390),
.A2(n_395),
.B1(n_322),
.B2(n_329),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_332),
.B(n_234),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_318),
.A2(n_254),
.B(n_233),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_392),
.A2(n_375),
.B(n_401),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_394),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_310),
.A2(n_364),
.B1(n_339),
.B2(n_307),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_311),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_407),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_SL g397 ( 
.A(n_354),
.B(n_226),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_397),
.A2(n_408),
.B(n_331),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_323),
.A2(n_328),
.B1(n_336),
.B2(n_335),
.Y(n_398)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_337),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_404),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_245),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_402),
.B(n_403),
.Y(n_417)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_324),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_405),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_323),
.A2(n_285),
.B1(n_308),
.B2(n_357),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_406),
.A2(n_322),
.B1(n_329),
.B2(n_320),
.Y(n_445)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

OR2x4_ASAP7_75t_L g408 ( 
.A(n_355),
.B(n_285),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_409),
.Y(n_435)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_412),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_361),
.B(n_306),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_411),
.B(n_355),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_360),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_330),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_414),
.B(n_426),
.C(n_422),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_395),
.A2(n_358),
.B1(n_341),
.B2(n_340),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_415),
.A2(n_434),
.B1(n_439),
.B2(n_442),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_418),
.B(n_407),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_423),
.B(n_388),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_373),
.A2(n_355),
.B1(n_307),
.B2(n_316),
.Y(n_425)
);

OA22x2_ASAP7_75t_L g474 ( 
.A1(n_425),
.A2(n_445),
.B1(n_449),
.B2(n_389),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_338),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_427),
.A2(n_392),
.B(n_366),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_369),
.B(n_327),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_430),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_391),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_386),
.B(n_359),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_438),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_380),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_383),
.A2(n_312),
.B1(n_315),
.B2(n_317),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_390),
.A2(n_315),
.B1(n_317),
.B2(n_313),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_406),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_368),
.Y(n_467)
);

XOR2x2_ASAP7_75t_SL g470 ( 
.A(n_446),
.B(n_371),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_447),
.A2(n_385),
.B1(n_396),
.B2(n_384),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_377),
.A2(n_321),
.B1(n_325),
.B2(n_337),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_432),
.Y(n_452)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_453),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_450),
.B(n_353),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_454),
.B(n_462),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_421),
.A2(n_399),
.B(n_408),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_456),
.B(n_463),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_420),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_457),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_414),
.B(n_399),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_460),
.C(n_475),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_372),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_461),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_353),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_348),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_464),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_348),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_465),
.B(n_472),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_466),
.B(n_446),
.Y(n_505)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_467),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_370),
.Y(n_468)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_419),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_476),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_471),
.Y(n_490)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_419),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_473),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_474),
.Y(n_500)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_477),
.A2(n_437),
.B1(n_416),
.B2(n_433),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_419),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_480),
.Y(n_493)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_481),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_443),
.A2(n_374),
.B(n_410),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_428),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_427),
.A2(n_412),
.B(n_400),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_483),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_429),
.B(n_394),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_485),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_416),
.B(n_409),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_321),
.C(n_325),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_487),
.C(n_418),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_423),
.B(n_349),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_482),
.A2(n_437),
.B1(n_425),
.B2(n_445),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_495),
.A2(n_517),
.B1(n_464),
.B2(n_461),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_496),
.A2(n_485),
.B1(n_474),
.B2(n_484),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_460),
.B(n_426),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_504),
.B(n_511),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_459),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_506),
.B(n_455),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_467),
.A2(n_415),
.B1(n_447),
.B2(n_439),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_508),
.A2(n_473),
.B1(n_476),
.B2(n_469),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_455),
.B(n_417),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_509),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_458),
.B(n_430),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_482),
.A2(n_424),
.B1(n_448),
.B2(n_449),
.Y(n_512)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

NOR2x1_ASAP7_75t_L g513 ( 
.A(n_468),
.B(n_442),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_513),
.A2(n_440),
.B(n_435),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_475),
.B(n_486),
.C(n_487),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_515),
.B(n_516),
.C(n_518),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_471),
.B(n_424),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_477),
.A2(n_441),
.B1(n_440),
.B2(n_451),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_470),
.B(n_451),
.C(n_441),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_456),
.B(n_413),
.C(n_428),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_472),
.C(n_480),
.Y(n_540)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_519),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_525),
.A2(n_529),
.B1(n_536),
.B2(n_542),
.Y(n_556)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_526),
.Y(n_559)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_499),
.Y(n_527)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_527),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_453),
.Y(n_528)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_510),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_530),
.B(n_532),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_493),
.A2(n_483),
.B(n_466),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_531),
.A2(n_546),
.B(n_488),
.Y(n_570)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_514),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_533),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_510),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_534),
.B(n_545),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_495),
.A2(n_481),
.B1(n_452),
.B2(n_478),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g561 ( 
.A(n_537),
.B(n_505),
.Y(n_561)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_502),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_538),
.B(n_544),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_540),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_511),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_508),
.A2(n_459),
.B1(n_474),
.B2(n_479),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_501),
.B(n_474),
.C(n_413),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_543),
.B(n_547),
.C(n_550),
.Y(n_562)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_507),
.Y(n_545)
);

NAND2x1_ASAP7_75t_L g546 ( 
.A(n_491),
.B(n_404),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_501),
.B(n_435),
.C(n_349),
.Y(n_547)
);

AOI21xp33_ASAP7_75t_L g548 ( 
.A1(n_489),
.A2(n_420),
.B(n_457),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_548),
.B(n_503),
.Y(n_571)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_502),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_549),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_515),
.B(n_345),
.C(n_334),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_557),
.B(n_566),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_542),
.A2(n_500),
.B1(n_497),
.B2(n_507),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_558),
.A2(n_533),
.B1(n_539),
.B2(n_536),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_561),
.B(n_564),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_535),
.B(n_504),
.Y(n_564)
);

FAx1_ASAP7_75t_SL g565 ( 
.A(n_537),
.B(n_491),
.CI(n_518),
.CON(n_565),
.SN(n_565)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_571),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_506),
.C(n_520),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_516),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_568),
.B(n_521),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_570),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_488),
.C(n_490),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_573),
.B(n_524),
.C(n_540),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_535),
.B(n_490),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_574),
.B(n_528),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_567),
.A2(n_523),
.B1(n_500),
.B2(n_538),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_575),
.A2(n_585),
.B1(n_556),
.B2(n_572),
.Y(n_595)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_555),
.Y(n_577)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_577),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_558),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_578),
.B(n_553),
.Y(n_602)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_579),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_589),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_563),
.A2(n_531),
.B(n_543),
.Y(n_584)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_584),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_567),
.A2(n_529),
.B1(n_549),
.B2(n_524),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_562),
.B(n_546),
.C(n_544),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_586),
.B(n_592),
.C(n_573),
.Y(n_597)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_552),
.Y(n_587)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_587),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_556),
.A2(n_551),
.B1(n_563),
.B2(n_569),
.Y(n_588)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_588),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_566),
.A2(n_525),
.B(n_522),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_590),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_593),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_562),
.B(n_546),
.C(n_517),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_557),
.B(n_521),
.Y(n_593)
);

XNOR2x1_ASAP7_75t_L g611 ( 
.A(n_595),
.B(n_597),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_584),
.B(n_431),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_596),
.B(n_600),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_580),
.B(n_564),
.C(n_553),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_593),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_576),
.B(n_568),
.C(n_574),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_605),
.B(n_606),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_592),
.B(n_561),
.C(n_565),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_498),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_607),
.B(n_583),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_586),
.C(n_589),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_610),
.B(n_617),
.Y(n_627)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_612),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_582),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_613),
.B(n_615),
.Y(n_628)
);

NOR2x1_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_575),
.Y(n_614)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_614),
.Y(n_630)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_603),
.Y(n_615)
);

AO21x1_ASAP7_75t_L g616 ( 
.A1(n_608),
.A2(n_583),
.B(n_582),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_616),
.B(n_619),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_598),
.B(n_559),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_594),
.B(n_585),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_620),
.B(n_595),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_604),
.B(n_581),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_622),
.B(n_604),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_624),
.A2(n_629),
.B(n_631),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_625),
.B(n_632),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_621),
.A2(n_600),
.B(n_606),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_610),
.A2(n_609),
.B1(n_565),
.B2(n_601),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_611),
.B(n_605),
.C(n_581),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_623),
.B(n_618),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_633),
.A2(n_634),
.B(n_636),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g634 ( 
.A1(n_627),
.A2(n_614),
.B(n_612),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_623),
.A2(n_611),
.B(n_616),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_628),
.B(n_622),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_638),
.B(n_630),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_635),
.B(n_632),
.C(n_626),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_639),
.B(n_640),
.Y(n_644)
);

O2A1O1Ixp33_ASAP7_75t_SL g642 ( 
.A1(n_637),
.A2(n_631),
.B(n_554),
.C(n_560),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_513),
.C(n_420),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_643),
.B(n_641),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_644),
.C(n_376),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_345),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_647),
.B(n_334),
.Y(n_648)
);


endmodule