module fake_jpeg_7938_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_16),
.B1(n_25),
.B2(n_30),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_48),
.B1(n_51),
.B2(n_55),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g80 ( 
.A(n_46),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_16),
.B1(n_25),
.B2(n_30),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_31),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_19),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_16),
.B1(n_25),
.B2(n_27),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_17),
.B1(n_21),
.B2(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_23),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_17),
.B1(n_21),
.B2(n_15),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_20),
.B1(n_19),
.B2(n_28),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_73),
.Y(n_94)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_34),
.B1(n_18),
.B2(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_82),
.B1(n_52),
.B2(n_19),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_9),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_20),
.B1(n_19),
.B2(n_22),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_22),
.B1(n_35),
.B2(n_33),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_0),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_1),
.Y(n_117)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_1),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_98),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_78),
.B1(n_85),
.B2(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_54),
.C(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_35),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_78),
.C(n_22),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_69),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_33),
.B(n_2),
.C(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_82),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_118),
.B(n_116),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_6),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_123),
.B(n_97),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_90),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_87),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_64),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_93),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_102),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_154),
.B(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_118),
.B(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_131),
.B(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_118),
.B1(n_96),
.B2(n_100),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_127),
.B1(n_101),
.B2(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_128),
.B1(n_141),
.B2(n_137),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_117),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_140),
.C(n_132),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_146),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_157),
.A2(n_134),
.B1(n_121),
.B2(n_123),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_164),
.C(n_169),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_155),
.C(n_148),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_111),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_177),
.C(n_154),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_175),
.A2(n_179),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_148),
.C(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_98),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_6),
.Y(n_188)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_142),
.B1(n_143),
.B2(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_154),
.B1(n_168),
.B2(n_139),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_169),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_182),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_185),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_2),
.B(n_3),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_12),
.B(n_8),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_12),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_172),
.B1(n_173),
.B2(n_112),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_192),
.Y(n_198)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_195),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_181),
.C(n_172),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_191),
.C(n_194),
.Y(n_200)
);

AOI31xp67_ASAP7_75t_SL g199 ( 
.A1(n_193),
.A2(n_186),
.A3(n_185),
.B(n_4),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_4),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_201),
.B(n_4),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_198),
.A2(n_194),
.B(n_197),
.C(n_3),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_113),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_72),
.Y(n_206)
);


endmodule