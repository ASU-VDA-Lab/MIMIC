module fake_jpeg_30663_n_158 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_158);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_31),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_1),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g35 ( 
.A1(n_21),
.A2(n_1),
.B(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_2),
.C(n_3),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_30),
.C(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_4),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_15),
.B1(n_29),
.B2(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_49),
.B1(n_13),
.B2(n_58),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_15),
.B1(n_29),
.B2(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_3),
.Y(n_67)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_26),
.B1(n_23),
.B2(n_16),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_59),
.B1(n_63),
.B2(n_10),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_3),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_33),
.A2(n_17),
.B1(n_14),
.B2(n_27),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_16),
.C(n_27),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_45),
.C(n_55),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_44),
.B1(n_37),
.B2(n_15),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_7),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_6),
.B(n_8),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_57),
.B(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_10),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_84),
.B1(n_79),
.B2(n_69),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_13),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_65),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_48),
.B1(n_54),
.B2(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_87),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_62),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_85),
.C(n_86),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_54),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_79),
.B1(n_71),
.B2(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_73),
.B(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_107),
.B1(n_94),
.B2(n_95),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_89),
.B1(n_104),
.B2(n_103),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_71),
.B(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_110),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_119),
.C(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_83),
.B1(n_104),
.B2(n_96),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_102),
.B(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_116),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_103),
.B1(n_95),
.B2(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_115),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_117),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_133),
.C(n_138),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_108),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_113),
.C(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_136),
.Y(n_144)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_125),
.B1(n_116),
.B2(n_121),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_141),
.B1(n_124),
.B2(n_127),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_126),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_126),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_135),
.C(n_120),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_147),
.C(n_148),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_138),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_92),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_141),
.B(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_150),
.B(n_148),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_91),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_154),
.B(n_151),
.Y(n_155)
);

INVxp33_ASAP7_75t_SL g156 ( 
.A(n_155),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_147),
.C(n_91),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_157),
.Y(n_158)
);


endmodule