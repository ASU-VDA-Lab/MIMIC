module fake_jpeg_15722_n_18 (n_3, n_2, n_1, n_0, n_4, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_18;

wire n_13;
wire n_11;
wire n_14;
wire n_17;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

NAND2xp5_ASAP7_75t_L g5 ( 
.A(n_1),
.B(n_2),
.Y(n_5)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

HAxp5_ASAP7_75t_SL g8 ( 
.A(n_3),
.B(n_0),
.CON(n_8),
.SN(n_8)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_5),
.A2(n_0),
.B(n_2),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_7),
.C(n_10),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_6),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_10)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_11),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_6),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_6),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_8),
.C(n_7),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_15),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_14),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_11),
.C(n_7),
.Y(n_18)
);


endmodule