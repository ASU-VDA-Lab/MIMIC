module fake_jpeg_22399_n_167 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_28),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_20),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_19),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_31),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_66),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_18),
.B1(n_31),
.B2(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_59),
.B1(n_21),
.B2(n_37),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_18),
.B1(n_17),
.B2(n_29),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_25),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_19),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_18),
.B1(n_17),
.B2(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_27),
.B1(n_23),
.B2(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_24),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_1),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_44),
.B(n_21),
.C(n_30),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_42),
.B(n_32),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_89),
.B(n_51),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_77),
.B(n_87),
.C(n_67),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_35),
.B1(n_42),
.B2(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_79),
.Y(n_98)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_37),
.A3(n_36),
.B1(n_19),
.B2(n_21),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_27),
.B1(n_23),
.B2(n_30),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_84),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_88),
.Y(n_92)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_3),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_36),
.B(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_63),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_89),
.B(n_68),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_83),
.B1(n_77),
.B2(n_91),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_45),
.B(n_58),
.C(n_53),
.D(n_49),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_73),
.C(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_106),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_3),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_110),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_47),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_87),
.C(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_10),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_93),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_113),
.C(n_119),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_116),
.B(n_107),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_118),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_79),
.C(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_72),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_126),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_78),
.C(n_48),
.Y(n_124)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_103),
.B(n_105),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_8),
.B(n_13),
.C(n_7),
.D(n_6),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_8),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_137),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_105),
.B(n_94),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_129),
.C(n_123),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_101),
.B1(n_76),
.B2(n_106),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_136),
.B1(n_114),
.B2(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_101),
.B1(n_104),
.B2(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_13),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_143),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_133),
.C(n_132),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_132),
.Y(n_151)
);

AOI21x1_ASAP7_75t_SL g149 ( 
.A1(n_147),
.A2(n_138),
.B(n_133),
.Y(n_149)
);

AOI31xp33_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_140),
.A3(n_144),
.B(n_142),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_157),
.C(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_154),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_158),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_142),
.A3(n_146),
.B1(n_127),
.B2(n_55),
.C1(n_6),
.C2(n_3),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_127),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_157),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_161),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_154),
.C(n_5),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_5),
.B(n_163),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_160),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_164),
.Y(n_167)
);


endmodule