module fake_jpeg_22055_n_70 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_66;

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_36),
.B(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_39),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_48),
.B1(n_40),
.B2(n_34),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_35),
.C(n_37),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_3),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_5),
.C(n_6),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_48),
.B(n_55),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_59),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_5),
.B(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_63),
.C(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_64),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_62),
.B(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_62),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_12),
.A3(n_14),
.B1(n_19),
.B2(n_21),
.C1(n_22),
.C2(n_23),
.Y(n_69)
);

A2O1A1O1Ixp25_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_25),
.B(n_26),
.C(n_27),
.D(n_28),
.Y(n_70)
);


endmodule