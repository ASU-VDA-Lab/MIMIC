module real_aes_7099_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g515 ( .A(n_1), .Y(n_515) );
INVx1_ASAP7_75t_L g156 ( .A(n_2), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_3), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_3), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_4), .A2(n_127), .B1(n_128), .B2(n_451), .Y(n_126) );
INVx1_ASAP7_75t_L g451 ( .A(n_4), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_5), .A2(n_40), .B1(n_181), .B2(n_471), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g200 ( .A1(n_6), .A2(n_172), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_7), .B(n_170), .Y(n_526) );
AND2x6_ASAP7_75t_L g149 ( .A(n_8), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_9), .A2(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_10), .B(n_41), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_10), .B(n_41), .Y(n_125) );
INVx1_ASAP7_75t_L g206 ( .A(n_11), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_12), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g141 ( .A(n_13), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_14), .B(n_162), .Y(n_479) );
INVx1_ASAP7_75t_L g260 ( .A(n_15), .Y(n_260) );
INVx1_ASAP7_75t_L g509 ( .A(n_16), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_17), .B(n_137), .Y(n_531) );
AO32x2_ASAP7_75t_L g498 ( .A1(n_18), .A2(n_136), .A3(n_170), .B1(n_473), .B2(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_19), .B(n_181), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_20), .B(n_177), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_21), .B(n_137), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_22), .A2(n_33), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_22), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_23), .A2(n_53), .B1(n_181), .B2(n_471), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_24), .B(n_172), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_25), .A2(n_79), .B1(n_162), .B2(n_181), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_26), .B(n_181), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_27), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_28), .A2(n_258), .B(n_259), .C(n_261), .Y(n_257) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_29), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_30), .B(n_167), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_31), .B(n_160), .Y(n_159) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_32), .A2(n_457), .B1(n_739), .B2(n_745), .C1(n_748), .C2(n_749), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_33), .Y(n_449) );
INVx1_ASAP7_75t_L g195 ( .A(n_34), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_35), .B(n_167), .Y(n_496) );
INVx2_ASAP7_75t_L g147 ( .A(n_36), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_37), .B(n_181), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_38), .B(n_167), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_39), .A2(n_149), .B(n_152), .C(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g193 ( .A(n_42), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_43), .B(n_160), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_44), .A2(n_104), .B1(n_112), .B2(n_752), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_45), .B(n_181), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_46), .B(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_47), .A2(n_89), .B1(n_224), .B2(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_48), .B(n_181), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_49), .B(n_181), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_50), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_51), .B(n_514), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_52), .B(n_172), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_54), .A2(n_63), .B1(n_162), .B2(n_181), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_55), .A2(n_152), .B1(n_162), .B2(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_56), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_57), .B(n_181), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g143 ( .A(n_58), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_59), .B(n_181), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_60), .A2(n_180), .B(n_204), .C(n_205), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_61), .Y(n_251) );
INVx1_ASAP7_75t_L g202 ( .A(n_62), .Y(n_202) );
INVx1_ASAP7_75t_L g150 ( .A(n_64), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_65), .B(n_181), .Y(n_516) );
INVx1_ASAP7_75t_L g140 ( .A(n_66), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_67), .Y(n_117) );
AO32x2_ASAP7_75t_L g468 ( .A1(n_68), .A2(n_170), .A3(n_229), .B1(n_469), .B2(n_473), .Y(n_468) );
INVx1_ASAP7_75t_L g548 ( .A(n_69), .Y(n_548) );
INVx1_ASAP7_75t_L g491 ( .A(n_70), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_71), .A2(n_78), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_71), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_SL g176 ( .A1(n_72), .A2(n_177), .B(n_178), .C(n_180), .Y(n_176) );
INVxp67_ASAP7_75t_L g179 ( .A(n_73), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_74), .B(n_162), .Y(n_492) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_76), .Y(n_198) );
INVx1_ASAP7_75t_L g244 ( .A(n_77), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_78), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_80), .A2(n_149), .B(n_152), .C(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_81), .B(n_471), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_82), .B(n_162), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_83), .B(n_157), .Y(n_220) );
INVx2_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_85), .B(n_177), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_86), .B(n_162), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_87), .A2(n_149), .B(n_152), .C(n_155), .Y(n_151) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_88), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g122 ( .A(n_88), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g460 ( .A(n_88), .B(n_124), .Y(n_460) );
INVx2_ASAP7_75t_L g738 ( .A(n_88), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_90), .A2(n_102), .B1(n_162), .B2(n_163), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_91), .B(n_167), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_92), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_93), .A2(n_149), .B(n_152), .C(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_94), .Y(n_239) );
INVx1_ASAP7_75t_L g175 ( .A(n_95), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_96), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_97), .B(n_157), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_98), .B(n_162), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_99), .B(n_170), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_100), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_101), .A2(n_172), .B(n_173), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_104), .Y(n_752) );
CKINVDCx12_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x2_ASAP7_75t_L g124 ( .A(n_108), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_455), .Y(n_112) );
BUFx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_114), .B(n_452), .C(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_126), .B(n_452), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_122), .Y(n_454) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_123), .B(n_738), .Y(n_751) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g737 ( .A(n_124), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_446), .B1(n_447), .B2(n_450), .Y(n_128) );
INVx2_ASAP7_75t_L g450 ( .A(n_129), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_129), .A2(n_458), .B1(n_461), .B2(n_735), .Y(n_457) );
OR4x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_335), .C(n_395), .D(n_422), .Y(n_129) );
NAND4xp25_ASAP7_75t_SL g130 ( .A(n_131), .B(n_283), .C(n_314), .D(n_331), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_208), .B(n_210), .C(n_263), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_186), .Y(n_132) );
INVx1_ASAP7_75t_L g325 ( .A(n_133), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_133), .A2(n_366), .B1(n_414), .B2(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_168), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_134), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g276 ( .A(n_134), .B(n_188), .Y(n_276) );
AND2x2_ASAP7_75t_L g318 ( .A(n_134), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_134), .B(n_209), .Y(n_330) );
INVx1_ASAP7_75t_L g370 ( .A(n_134), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_134), .B(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g298 ( .A(n_135), .B(n_188), .Y(n_298) );
INVx3_ASAP7_75t_L g302 ( .A(n_135), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_135), .B(n_360), .Y(n_359) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_142), .B(n_164), .Y(n_135) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_136), .A2(n_189), .B(n_197), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_136), .B(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g225 ( .A(n_136), .Y(n_225) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_138), .B(n_139), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_151), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_144), .A2(n_182), .B1(n_190), .B2(n_196), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_144), .A2(n_244), .B(n_245), .Y(n_243) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
AND2x4_ASAP7_75t_L g172 ( .A(n_145), .B(n_149), .Y(n_172) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g514 ( .A(n_146), .Y(n_514) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx3_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
INVx1_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_148), .Y(n_192) );
INVx4_ASAP7_75t_SL g182 ( .A(n_149), .Y(n_182) );
BUFx3_ASAP7_75t_L g473 ( .A(n_149), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_149), .A2(n_477), .B(n_481), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_149), .A2(n_490), .B(n_493), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_149), .A2(n_508), .B(n_512), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_149), .A2(n_520), .B(n_523), .Y(n_519) );
INVx5_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
BUFx3_ASAP7_75t_L g224 ( .A(n_153), .Y(n_224) );
INVx1_ASAP7_75t_L g471 ( .A(n_153), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_159), .C(n_161), .Y(n_155) );
O2A1O1Ixp5_ASAP7_75t_SL g490 ( .A1(n_157), .A2(n_180), .B(n_491), .C(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g501 ( .A(n_157), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_157), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_157), .A2(n_545), .B(n_546), .Y(n_544) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_158), .B(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_158), .B(n_206), .Y(n_205) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_158), .A2(n_160), .B1(n_470), .B2(n_472), .Y(n_469) );
INVx2_ASAP7_75t_L g204 ( .A(n_160), .Y(n_204) );
INVx4_ASAP7_75t_L g235 ( .A(n_160), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_160), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_160), .A2(n_501), .B1(n_534), .B2(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_161), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_166), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_166), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g229 ( .A(n_167), .Y(n_229) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_167), .A2(n_253), .B(n_262), .Y(n_252) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_167), .A2(n_476), .B(n_484), .Y(n_475) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_167), .A2(n_489), .B(n_496), .Y(n_488) );
AND2x2_ASAP7_75t_L g389 ( .A(n_168), .B(n_199), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_168), .B(n_302), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_168), .B(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g209 ( .A(n_169), .B(n_188), .Y(n_209) );
INVx1_ASAP7_75t_L g271 ( .A(n_169), .Y(n_271) );
BUFx2_ASAP7_75t_L g275 ( .A(n_169), .Y(n_275) );
AND2x2_ASAP7_75t_L g319 ( .A(n_169), .B(n_187), .Y(n_319) );
OR2x2_ASAP7_75t_L g358 ( .A(n_169), .B(n_187), .Y(n_358) );
AND2x2_ASAP7_75t_L g383 ( .A(n_169), .B(n_199), .Y(n_383) );
AND2x2_ASAP7_75t_L g442 ( .A(n_169), .B(n_272), .Y(n_442) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_183), .Y(n_169) );
INVx4_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_170), .A2(n_519), .B(n_526), .Y(n_518) );
BUFx2_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_182), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_174), .A2(n_182), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_174), .A2(n_182), .B(n_256), .C(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g480 ( .A(n_177), .Y(n_480) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_181), .Y(n_236) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_184), .A2(n_200), .B(n_207), .Y(n_199) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g226 ( .A(n_185), .B(n_227), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_185), .B(n_473), .C(n_533), .Y(n_532) );
AO21x1_ASAP7_75t_L g579 ( .A1(n_185), .A2(n_533), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g417 ( .A(n_186), .Y(n_417) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_199), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_187), .B(n_199), .Y(n_303) );
AND2x2_ASAP7_75t_L g313 ( .A(n_187), .B(n_302), .Y(n_313) );
BUFx2_ASAP7_75t_L g324 ( .A(n_187), .Y(n_324) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g346 ( .A(n_188), .B(n_199), .Y(n_346) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_188), .Y(n_401) );
OAI22xp5_ASAP7_75t_SL g191 ( .A1(n_192), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_191) );
INVx2_ASAP7_75t_L g194 ( .A(n_192), .Y(n_194) );
INVx4_ASAP7_75t_L g258 ( .A(n_192), .Y(n_258) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_199), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_SL g272 ( .A(n_199), .Y(n_272) );
BUFx2_ASAP7_75t_L g297 ( .A(n_199), .Y(n_297) );
INVx2_ASAP7_75t_L g316 ( .A(n_199), .Y(n_316) );
AND2x2_ASAP7_75t_L g378 ( .A(n_199), .B(n_302), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_204), .A2(n_482), .B(n_483), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_L g547 ( .A1(n_204), .A2(n_513), .B(n_548), .C(n_549), .Y(n_547) );
AOI321xp33_ASAP7_75t_L g397 ( .A1(n_208), .A2(n_398), .A3(n_399), .B1(n_400), .B2(n_402), .C(n_403), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_209), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_209), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g391 ( .A(n_209), .B(n_370), .Y(n_391) );
AND2x2_ASAP7_75t_L g424 ( .A(n_209), .B(n_316), .Y(n_424) );
INVx1_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_240), .Y(n_211) );
OR2x2_ASAP7_75t_L g326 ( .A(n_212), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_228), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g278 ( .A(n_215), .Y(n_278) );
AND2x2_ASAP7_75t_L g288 ( .A(n_215), .B(n_242), .Y(n_288) );
AND2x2_ASAP7_75t_L g293 ( .A(n_215), .B(n_268), .Y(n_293) );
INVx1_ASAP7_75t_L g310 ( .A(n_215), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_215), .B(n_291), .Y(n_329) );
AND2x2_ASAP7_75t_L g334 ( .A(n_215), .B(n_267), .Y(n_334) );
OR2x2_ASAP7_75t_L g366 ( .A(n_215), .B(n_355), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_215), .B(n_279), .Y(n_405) );
AND2x2_ASAP7_75t_L g439 ( .A(n_215), .B(n_265), .Y(n_439) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
AOI21xp5_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_218), .B(n_225), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g261 ( .A(n_224), .Y(n_261) );
INVx1_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_225), .A2(n_507), .B(n_517), .Y(n_506) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_225), .A2(n_543), .B(n_550), .Y(n_542) );
INVx1_ASAP7_75t_L g266 ( .A(n_228), .Y(n_266) );
INVx2_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
AND2x2_ASAP7_75t_L g321 ( .A(n_228), .B(n_292), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_228), .B(n_268), .Y(n_343) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_238), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_236), .Y(n_232) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g427 ( .A(n_241), .B(n_278), .Y(n_427) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_252), .Y(n_241) );
INVx2_ASAP7_75t_L g268 ( .A(n_242), .Y(n_268) );
AND2x2_ASAP7_75t_L g421 ( .A(n_242), .B(n_281), .Y(n_421) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_249), .B(n_250), .Y(n_242) );
AND2x2_ASAP7_75t_L g267 ( .A(n_252), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g282 ( .A(n_252), .Y(n_282) );
INVx1_ASAP7_75t_L g292 ( .A(n_252), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_258), .B(n_260), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_258), .A2(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g511 ( .A(n_258), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_269), .B1(n_273), .B2(n_277), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_264), .A2(n_382), .B1(n_419), .B2(n_420), .Y(n_418) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g333 ( .A(n_266), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_267), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g328 ( .A(n_268), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_268), .B(n_281), .Y(n_355) );
INVx1_ASAP7_75t_L g371 ( .A(n_268), .Y(n_371) );
AND2x2_ASAP7_75t_L g312 ( .A(n_270), .B(n_313), .Y(n_312) );
INVx3_ASAP7_75t_SL g351 ( .A(n_270), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_270), .B(n_276), .Y(n_428) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g437 ( .A(n_273), .Y(n_437) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_274), .B(n_370), .Y(n_412) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx3_ASAP7_75t_SL g317 ( .A(n_276), .Y(n_317) );
NAND2x1_ASAP7_75t_SL g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g338 ( .A(n_278), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g345 ( .A(n_278), .B(n_282), .Y(n_345) );
AND2x2_ASAP7_75t_L g350 ( .A(n_278), .B(n_291), .Y(n_350) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_278), .Y(n_399) );
OAI311xp33_ASAP7_75t_L g422 ( .A1(n_279), .A2(n_423), .A3(n_425), .B1(n_426), .C1(n_436), .Y(n_422) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g435 ( .A(n_280), .B(n_308), .Y(n_435) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g291 ( .A(n_281), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g339 ( .A(n_281), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g394 ( .A(n_281), .Y(n_394) );
INVx1_ASAP7_75t_L g287 ( .A(n_282), .Y(n_287) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_282), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g340 ( .A(n_282), .Y(n_340) );
AOI221xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_286), .B1(n_294), .B2(n_299), .C(n_304), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_289), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx4_ASAP7_75t_L g308 ( .A(n_288), .Y(n_308) );
AND2x2_ASAP7_75t_L g402 ( .A(n_288), .B(n_321), .Y(n_402) );
AND2x2_ASAP7_75t_L g409 ( .A(n_288), .B(n_291), .Y(n_409) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_291), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g320 ( .A(n_293), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_296), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g445 ( .A(n_298), .B(n_389), .Y(n_445) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g430 ( .A(n_302), .B(n_358), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g395 ( .A1(n_303), .A2(n_396), .B(n_397), .C(n_410), .Y(n_395) );
AOI21xp33_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_309), .B(n_311), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp67_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g374 ( .A(n_308), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_309), .A2(n_404), .B1(n_405), .B2(n_406), .C(n_407), .Y(n_403) );
AND2x2_ASAP7_75t_L g380 ( .A(n_310), .B(n_321), .Y(n_380) );
AND2x2_ASAP7_75t_L g433 ( .A(n_310), .B(n_328), .Y(n_433) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_313), .B(n_351), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_320), .C(n_322), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g361 ( .A(n_316), .B(n_319), .Y(n_361) );
OR2x2_ASAP7_75t_L g404 ( .A(n_316), .B(n_358), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_317), .B(n_383), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_317), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g348 ( .A(n_318), .Y(n_348) );
INVx1_ASAP7_75t_L g414 ( .A(n_321), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B1(n_329), .B2(n_330), .Y(n_322) );
INVx1_ASAP7_75t_L g337 ( .A(n_323), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_324), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g400 ( .A(n_325), .B(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g386 ( .A(n_327), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_328), .B(n_414), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_329), .A2(n_388), .B1(n_390), .B2(n_392), .Y(n_387) );
INVx1_ASAP7_75t_L g396 ( .A(n_332), .Y(n_396) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g438 ( .A(n_333), .B(n_433), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_334), .A2(n_368), .B1(n_371), .B2(n_372), .C1(n_375), .C2(n_376), .Y(n_367) );
NAND4xp25_ASAP7_75t_SL g335 ( .A(n_336), .B(n_356), .C(n_367), .D(n_379), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_341), .B2(n_346), .C(n_347), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_339), .B(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g365 ( .A(n_340), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_341), .A2(n_411), .B1(n_413), .B2(n_415), .C(n_418), .Y(n_410) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g353 ( .A(n_345), .B(n_354), .Y(n_353) );
OAI21xp33_ASAP7_75t_L g407 ( .A1(n_346), .A2(n_408), .B(n_409), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_351), .B2(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_362), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_370), .B(n_389), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_370), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_374), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g406 ( .A(n_378), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_384), .B2(n_386), .C(n_387), .Y(n_379) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI222xp33_ASAP7_75t_L g426 ( .A1(n_389), .A2(n_427), .B1(n_428), .B2(n_429), .C1(n_431), .C2(n_434), .Y(n_426) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_393), .B(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g425 ( .A(n_399), .Y(n_425) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp33_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_439), .B2(n_440), .C(n_443), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_450), .A2(n_458), .B1(n_746), .B2(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g747 ( .A(n_461), .Y(n_747) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND3x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_655), .C(n_703), .Y(n_462) );
NOR4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_583), .C(n_628), .D(n_642), .Y(n_463) );
OAI311xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_503), .A3(n_527), .B1(n_536), .C1(n_551), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_474), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_466), .A2(n_537), .B(n_539), .Y(n_536) );
AND2x2_ASAP7_75t_L g644 ( .A(n_466), .B(n_571), .Y(n_644) );
AND2x2_ASAP7_75t_L g701 ( .A(n_466), .B(n_587), .Y(n_701) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g594 ( .A(n_467), .B(n_497), .Y(n_594) );
AND2x2_ASAP7_75t_L g651 ( .A(n_467), .B(n_599), .Y(n_651) );
INVx1_ASAP7_75t_L g692 ( .A(n_467), .Y(n_692) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_468), .Y(n_560) );
AND2x2_ASAP7_75t_L g601 ( .A(n_468), .B(n_497), .Y(n_601) );
AND2x2_ASAP7_75t_L g605 ( .A(n_468), .B(n_498), .Y(n_605) );
INVx1_ASAP7_75t_L g617 ( .A(n_468), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_473), .A2(n_544), .B(n_547), .Y(n_543) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .Y(n_474) );
AND2x2_ASAP7_75t_L g538 ( .A(n_475), .B(n_497), .Y(n_538) );
INVx2_ASAP7_75t_L g572 ( .A(n_475), .Y(n_572) );
AND2x2_ASAP7_75t_L g587 ( .A(n_475), .B(n_498), .Y(n_587) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_475), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_475), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g607 ( .A(n_475), .B(n_570), .Y(n_607) );
INVx1_ASAP7_75t_L g619 ( .A(n_475), .Y(n_619) );
INVx1_ASAP7_75t_L g660 ( .A(n_475), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_475), .B(n_560), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_480), .Y(n_477) );
NOR2xp67_ASAP7_75t_L g485 ( .A(n_486), .B(n_497), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g537 ( .A(n_487), .B(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_487), .Y(n_565) );
AND2x2_ASAP7_75t_SL g618 ( .A(n_487), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g622 ( .A(n_487), .B(n_497), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_487), .B(n_617), .Y(n_680) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g570 ( .A(n_488), .Y(n_570) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_488), .Y(n_586) );
OR2x2_ASAP7_75t_L g659 ( .A(n_488), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g566 ( .A(n_498), .Y(n_566) );
AND2x2_ASAP7_75t_L g571 ( .A(n_498), .B(n_572), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_501), .A2(n_513), .B(n_515), .C(n_516), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_501), .A2(n_524), .B(n_525), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_503), .B(n_554), .Y(n_717) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g687 ( .A(n_504), .B(n_529), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_518), .Y(n_504) );
AND2x2_ASAP7_75t_L g563 ( .A(n_505), .B(n_554), .Y(n_563) );
INVx2_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
AND2x2_ASAP7_75t_L g609 ( .A(n_505), .B(n_557), .Y(n_609) );
AND2x2_ASAP7_75t_L g676 ( .A(n_505), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_506), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g556 ( .A(n_506), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g596 ( .A(n_506), .B(n_518), .Y(n_596) );
AND2x2_ASAP7_75t_L g613 ( .A(n_506), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g539 ( .A(n_518), .B(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g557 ( .A(n_518), .Y(n_557) );
AND2x2_ASAP7_75t_L g562 ( .A(n_518), .B(n_542), .Y(n_562) );
AND2x2_ASAP7_75t_L g635 ( .A(n_518), .B(n_614), .Y(n_635) );
AND2x2_ASAP7_75t_L g700 ( .A(n_518), .B(n_690), .Y(n_700) );
OAI311xp33_ASAP7_75t_L g583 ( .A1(n_527), .A2(n_584), .A3(n_588), .B1(n_590), .C1(n_610), .Y(n_583) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g595 ( .A(n_528), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g654 ( .A(n_528), .B(n_562), .Y(n_654) );
AND2x2_ASAP7_75t_L g728 ( .A(n_528), .B(n_609), .Y(n_728) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_529), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g663 ( .A(n_529), .Y(n_663) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g554 ( .A(n_530), .Y(n_554) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_530), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g683 ( .A(n_530), .B(n_557), .Y(n_683) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g580 ( .A(n_531), .Y(n_580) );
AND2x2_ASAP7_75t_L g558 ( .A(n_538), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g611 ( .A(n_538), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g691 ( .A(n_538), .B(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_539), .A2(n_571), .B1(n_591), .B2(n_595), .C(n_597), .Y(n_590) );
INVx1_ASAP7_75t_L g715 ( .A(n_540), .Y(n_715) );
OR2x2_ASAP7_75t_L g681 ( .A(n_541), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g576 ( .A(n_542), .B(n_557), .Y(n_576) );
OR2x2_ASAP7_75t_L g578 ( .A(n_542), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g603 ( .A(n_542), .Y(n_603) );
INVx2_ASAP7_75t_L g614 ( .A(n_542), .Y(n_614) );
AND2x2_ASAP7_75t_L g641 ( .A(n_542), .B(n_579), .Y(n_641) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_542), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_558), .B1(n_561), .B2(n_564), .C(n_567), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g652 ( .A(n_554), .B(n_562), .Y(n_652) );
AND2x2_ASAP7_75t_L g702 ( .A(n_554), .B(n_556), .Y(n_702) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g589 ( .A(n_556), .B(n_560), .Y(n_589) );
AND2x2_ASAP7_75t_L g668 ( .A(n_556), .B(n_641), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_557), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g627 ( .A(n_557), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_558), .A2(n_638), .B(n_640), .Y(n_637) );
OR2x2_ASAP7_75t_L g581 ( .A(n_559), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g647 ( .A(n_559), .B(n_607), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_559), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g624 ( .A(n_560), .B(n_593), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_560), .B(n_707), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_561), .B(n_587), .Y(n_697) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g620 ( .A(n_562), .B(n_575), .Y(n_620) );
INVx1_ASAP7_75t_L g636 ( .A(n_563), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_573), .B1(n_577), .B2(n_581), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx2_ASAP7_75t_L g599 ( .A(n_570), .Y(n_599) );
INVx1_ASAP7_75t_L g612 ( .A(n_570), .Y(n_612) );
INVx1_ASAP7_75t_L g582 ( .A(n_571), .Y(n_582) );
AND2x2_ASAP7_75t_L g653 ( .A(n_571), .B(n_599), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_571), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
OR2x2_ASAP7_75t_L g577 ( .A(n_574), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_574), .B(n_690), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_574), .B(n_722), .Y(n_721) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g724 ( .A(n_576), .B(n_676), .Y(n_724) );
INVx1_ASAP7_75t_SL g690 ( .A(n_578), .Y(n_690) );
AND2x2_ASAP7_75t_L g630 ( .A(n_579), .B(n_614), .Y(n_630) );
INVx1_ASAP7_75t_L g677 ( .A(n_579), .Y(n_677) );
OAI222xp33_ASAP7_75t_L g718 ( .A1(n_584), .A2(n_674), .B1(n_719), .B2(n_720), .C1(n_723), .C2(n_725), .Y(n_718) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g639 ( .A(n_586), .Y(n_639) );
AND2x2_ASAP7_75t_L g650 ( .A(n_587), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_587), .B(n_692), .Y(n_719) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_589), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g694 ( .A(n_591), .Y(n_694) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g632 ( .A(n_594), .Y(n_632) );
AND2x2_ASAP7_75t_L g711 ( .A(n_594), .B(n_672), .Y(n_711) );
AND2x2_ASAP7_75t_L g734 ( .A(n_594), .B(n_618), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_596), .B(n_630), .Y(n_629) );
OAI32xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .A3(n_602), .B1(n_604), .B2(n_608), .Y(n_597) );
BUFx2_ASAP7_75t_L g672 ( .A(n_599), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_600), .B(n_618), .Y(n_699) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g638 ( .A(n_601), .B(n_639), .Y(n_638) );
AND2x4_ASAP7_75t_L g706 ( .A(n_601), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g695 ( .A(n_602), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AND2x2_ASAP7_75t_L g666 ( .A(n_605), .B(n_639), .Y(n_666) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_SL g628 ( .A1(n_607), .A2(n_629), .B1(n_631), .B2(n_633), .C(n_637), .Y(n_628) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g640 ( .A(n_609), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g646 ( .A(n_609), .B(n_630), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B1(n_615), .B2(n_620), .C(n_621), .Y(n_610) );
INVx1_ASAP7_75t_L g729 ( .A(n_611), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_612), .B(n_706), .Y(n_705) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_613), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_618), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g684 ( .A(n_618), .Y(n_684) );
BUFx3_ASAP7_75t_L g707 ( .A(n_619), .Y(n_707) );
INVx1_ASAP7_75t_SL g648 ( .A(n_620), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_620), .B(n_662), .Y(n_661) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_623), .B(n_625), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_622), .A2(n_723), .B1(n_727), .B2(n_729), .C(n_730), .Y(n_726) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g669 ( .A(n_627), .B(n_630), .Y(n_669) );
INVx1_ASAP7_75t_L g733 ( .A(n_627), .Y(n_733) );
INVx2_ASAP7_75t_L g722 ( .A(n_630), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_630), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g675 ( .A(n_635), .B(n_676), .Y(n_675) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_648), .C(n_649), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_653), .B2(n_654), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_651), .A2(n_713), .B1(n_714), .B2(n_716), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_654), .A2(n_731), .B(n_734), .Y(n_730) );
NOR4xp25_ASAP7_75t_SL g655 ( .A(n_656), .B(n_664), .C(n_673), .D(n_693), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_661), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B1(n_670), .B2(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g709 ( .A(n_669), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_678), .B1(n_681), .B2(n_684), .C(n_685), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g696 ( .A(n_676), .Y(n_696) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_688), .B(n_691), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_697), .C(n_698), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_698) );
CKINVDCx14_ASAP7_75t_R g708 ( .A(n_702), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_718), .C(n_726), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B1(n_709), .B2(n_710), .C(n_712), .Y(n_704) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g746 ( .A(n_736), .Y(n_746) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx16_ASAP7_75t_R g748 ( .A(n_739), .Y(n_748) );
INVx1_ASAP7_75t_L g743 ( .A(n_740), .Y(n_743) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx3_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
endmodule