module fake_jpeg_7619_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_17),
.Y(n_66)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_49),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_62),
.B1(n_17),
.B2(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_65),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_42),
.B(n_26),
.C(n_16),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_19),
.B1(n_25),
.B2(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_20),
.B1(n_30),
.B2(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_20),
.B1(n_30),
.B2(n_25),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_24),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_85),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_41),
.B1(n_43),
.B2(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_82),
.B1(n_84),
.B2(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_42),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_88),
.B1(n_91),
.B2(n_69),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_39),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_62),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_46),
.B1(n_41),
.B2(n_43),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_41),
.B1(n_42),
.B2(n_39),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_93),
.B(n_42),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_45),
.A2(n_34),
.B1(n_28),
.B2(n_20),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_28),
.B1(n_24),
.B2(n_32),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_36),
.B1(n_35),
.B2(n_27),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_66),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_99),
.C(n_108),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_97),
.B(n_107),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_56),
.B1(n_57),
.B2(n_36),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_105),
.B1(n_111),
.B2(n_27),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_48),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_68),
.B1(n_22),
.B2(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_76),
.B(n_86),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_110),
.B(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_68),
.B1(n_22),
.B2(n_23),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_121),
.B1(n_92),
.B2(n_27),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_48),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_119),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_76),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_77),
.B(n_23),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_77),
.B1(n_94),
.B2(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

OA22x2_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_83),
.B1(n_68),
.B2(n_44),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_128),
.B(n_150),
.Y(n_160)
);

AO21x2_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_83),
.B(n_48),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_103),
.B(n_119),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_90),
.B1(n_78),
.B2(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_139),
.B1(n_144),
.B2(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_98),
.B1(n_123),
.B2(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_149),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_145),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_44),
.B1(n_67),
.B2(n_54),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_55),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_44),
.B1(n_67),
.B2(n_52),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_55),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_118),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_107),
.C(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_26),
.B(n_16),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_162),
.C(n_148),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_159),
.B(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_164),
.B1(n_177),
.B2(n_128),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_158),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_116),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_163),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_10),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_166),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_10),
.Y(n_166)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_173),
.B(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_98),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_26),
.B(n_16),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_0),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_0),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_26),
.B(n_2),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_190),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_145),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_130),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_150),
.C(n_147),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_162),
.C(n_151),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_158),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_133),
.B1(n_125),
.B2(n_139),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_197),
.B1(n_202),
.B2(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_125),
.B1(n_128),
.B2(n_132),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_177),
.B(n_178),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_200),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_128),
.B1(n_127),
.B2(n_144),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_131),
.C(n_128),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_129),
.B1(n_124),
.B2(n_126),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_126),
.B1(n_137),
.B2(n_136),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_162),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_215),
.C(n_216),
.Y(n_232)
);

BUFx4f_ASAP7_75t_SL g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_204),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_213),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_160),
.B(n_174),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_210),
.B1(n_196),
.B2(n_185),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_174),
.B(n_160),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_157),
.B1(n_154),
.B2(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_170),
.B1(n_153),
.B2(n_155),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_212),
.A2(n_219),
.B1(n_167),
.B2(n_26),
.Y(n_247)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_160),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_227),
.B1(n_196),
.B2(n_185),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_157),
.B1(n_197),
.B2(n_193),
.Y(n_219)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_189),
.B(n_174),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_165),
.Y(n_244)
);

XOR2x1_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_173),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_229),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_181),
.A2(n_199),
.B1(n_180),
.B2(n_200),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_173),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_164),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_180),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_241),
.B(n_217),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_179),
.C(n_159),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_243),
.C(n_249),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_207),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_248),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_176),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_239),
.B(n_220),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_136),
.C(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_167),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_218),
.B1(n_210),
.B2(n_221),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_26),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_54),
.C(n_52),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_52),
.B1(n_8),
.B2(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_14),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_229),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_252),
.B(n_261),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_267),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_220),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_268),
.B(n_248),
.Y(n_283)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_207),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_245),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_249),
.C(n_232),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_278),
.C(n_266),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_240),
.B1(n_245),
.B2(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_276),
.B1(n_14),
.B2(n_13),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_209),
.B(n_212),
.C(n_210),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_280),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_232),
.C(n_243),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_262),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_264),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_258),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_265),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_285),
.B(n_287),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_267),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_290),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_289),
.B(n_296),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_262),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_269),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_274),
.B(n_12),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_293),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_257),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_297),
.B(n_1),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_295),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_13),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_284),
.C(n_276),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_2),
.B(n_3),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_301),
.C(n_307),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_11),
.A3(n_8),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_6),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_305),
.Y(n_314)
);

BUFx4f_ASAP7_75t_SL g305 ( 
.A(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_2),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_3),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_312),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_304),
.A2(n_294),
.B1(n_287),
.B2(n_4),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_2),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_5),
.B(n_7),
.C(n_314),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_305),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_301),
.C(n_6),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_320),
.A2(n_318),
.B(n_319),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_321),
.C(n_7),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_7),
.Y(n_325)
);


endmodule