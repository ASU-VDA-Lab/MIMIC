module fake_jpeg_14482_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx12f_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_39),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_0),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_39),
.C(n_31),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_14),
.Y(n_90)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_1),
.Y(n_70)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_69),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_16),
.B(n_39),
.C(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_66),
.B(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_28),
.B1(n_33),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_81),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_43),
.B(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_71),
.B(n_73),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_27),
.B1(n_28),
.B2(n_23),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_93),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_27),
.B1(n_28),
.B2(n_23),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_39),
.B1(n_17),
.B2(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_35),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_90),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_86),
.B(n_88),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_17),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_55),
.B1(n_44),
.B2(n_59),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_41),
.B(n_29),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_38),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_61),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_30),
.B1(n_25),
.B2(n_18),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_62),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_45),
.B(n_34),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_10),
.Y(n_111)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_31),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_111),
.B(n_117),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_116),
.A2(n_132),
.B1(n_110),
.B2(n_12),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_30),
.C(n_18),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_30),
.B1(n_18),
.B2(n_5),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_131),
.B1(n_92),
.B2(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_3),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_139),
.Y(n_161)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_65),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_65),
.B(n_6),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_9),
.C(n_10),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_105),
.B1(n_92),
.B2(n_63),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_149),
.A2(n_171),
.B1(n_129),
.B2(n_140),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_67),
.B1(n_91),
.B2(n_108),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_153),
.B1(n_160),
.B2(n_173),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_79),
.B1(n_98),
.B2(n_75),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_80),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_83),
.B1(n_80),
.B2(n_110),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_168),
.B1(n_124),
.B2(n_119),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_98),
.B1(n_75),
.B2(n_79),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_130),
.B(n_126),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_163),
.A2(n_172),
.B(n_175),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_96),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_165),
.B(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_101),
.B1(n_87),
.B2(n_83),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_87),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_172),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_72),
.B1(n_96),
.B2(n_99),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_99),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_101),
.B1(n_110),
.B2(n_72),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_11),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_161),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_120),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_183),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_151),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_214),
.C(n_194),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_145),
.B1(n_131),
.B2(n_125),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_199),
.B1(n_158),
.B2(n_174),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_203),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_137),
.B(n_112),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_206),
.B(n_211),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_112),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_212),
.Y(n_219)
);

XOR2x1_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_117),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_160),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_114),
.B1(n_138),
.B2(n_141),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_215),
.Y(n_240)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_114),
.B1(n_138),
.B2(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_209),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_148),
.B(n_111),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_210),
.B(n_213),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_173),
.A2(n_13),
.B1(n_134),
.B2(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_206),
.B(n_205),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_159),
.A2(n_175),
.B1(n_161),
.B2(n_176),
.Y(n_215)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_167),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_207),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_220),
.B(n_222),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_230),
.B1(n_233),
.B2(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_191),
.C(n_184),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_158),
.C(n_178),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_164),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_182),
.B1(n_164),
.B2(n_169),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_185),
.A2(n_211),
.B1(n_199),
.B2(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_213),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_185),
.A2(n_205),
.B1(n_196),
.B2(n_206),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_190),
.B(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_235),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_202),
.B1(n_190),
.B2(n_209),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_223),
.B1(n_243),
.B2(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_240),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_200),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_220),
.C(n_234),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_187),
.B1(n_197),
.B2(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_187),
.B1(n_219),
.B2(n_228),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_219),
.A2(n_241),
.B(n_231),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_227),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_238),
.Y(n_264)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_266),
.B(n_230),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_249),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_245),
.A2(n_234),
.B1(n_233),
.B2(n_231),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_222),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_277),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_279),
.C(n_283),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_249),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_229),
.C(n_225),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_267),
.B(n_237),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_284),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_237),
.C(n_257),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_237),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_252),
.C(n_260),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_276),
.C(n_281),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_254),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_273),
.A2(n_261),
.B(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

INVx11_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_301),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_271),
.C(n_283),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_250),
.B(n_272),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_279),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_308),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_278),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_290),
.B(n_292),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_311),
.Y(n_320)
);

OAI322xp33_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_259),
.A3(n_296),
.B1(n_286),
.B2(n_258),
.C1(n_295),
.C2(n_288),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_291),
.C(n_247),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_308),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_309),
.B1(n_305),
.B2(n_285),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.C(n_315),
.Y(n_323)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_319),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_305),
.B1(n_303),
.B2(n_302),
.Y(n_319)
);

AOI222xp33_ASAP7_75t_SL g321 ( 
.A1(n_318),
.A2(n_302),
.B1(n_315),
.B2(n_299),
.C1(n_304),
.C2(n_306),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_319),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_312),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_323),
.B(n_317),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_324),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_329),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_324),
.Y(n_331)
);


endmodule