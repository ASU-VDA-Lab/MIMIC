module fake_ariane_2479_n_2073 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2073);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2073;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_2016;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_40),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_95),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_25),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_127),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_34),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_58),
.Y(n_207)
);

BUFx8_ASAP7_75t_SL g208 ( 
.A(n_152),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_27),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_40),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_137),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_117),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_89),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_80),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_75),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_20),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_76),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_52),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_38),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_94),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_38),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_56),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_105),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_109),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_23),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_47),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_196),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_193),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_59),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_159),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_125),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_53),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_3),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_44),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_122),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_56),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_134),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_192),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_79),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_108),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_171),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_36),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_65),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_37),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_138),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_92),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_33),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_99),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_115),
.Y(n_261)
);

INVx4_ASAP7_75t_R g262 ( 
.A(n_42),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_67),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_79),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_124),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_87),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_145),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_150),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_161),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_176),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_163),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_151),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_67),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_103),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_155),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_184),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_48),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_133),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_147),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_36),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_188),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_1),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_114),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_119),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_154),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_91),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_123),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_169),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_189),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_166),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_198),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_5),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_5),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_45),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_14),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_160),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_106),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_149),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_4),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_86),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_112),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_165),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_46),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_187),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_31),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_81),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_46),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_59),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_10),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_22),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_42),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_98),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_11),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_44),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_62),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_186),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_74),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_14),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_61),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_27),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_175),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_164),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_34),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_31),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_70),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_174),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_3),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_43),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_173),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_13),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_25),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_179),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_185),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_83),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_32),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_35),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_191),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_52),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_70),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_178),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_97),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_121),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_82),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_9),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_172),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_180),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_77),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_162),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_85),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_22),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_139),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_116),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_39),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_100),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_167),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_43),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_148),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_181),
.Y(n_365)
);

BUFx8_ASAP7_75t_SL g366 ( 
.A(n_18),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_93),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_41),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_4),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_51),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_63),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_51),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_19),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_41),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_156),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_21),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_53),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_157),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_68),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_1),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_101),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_78),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_35),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_48),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_60),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_68),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_9),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_50),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_19),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_135),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_72),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_55),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_263),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_366),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_250),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_263),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_208),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_237),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_263),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_263),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_253),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_268),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_274),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_302),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_2),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_263),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_263),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_263),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_263),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_2),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_263),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_204),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_204),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_212),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_307),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_212),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_215),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_215),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_219),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_223),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_223),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_207),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_380),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_380),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_239),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_243),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_217),
.B(n_6),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_256),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_298),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_223),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_203),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_297),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_201),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_332),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_219),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_225),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_225),
.A2(n_199),
.B(n_195),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_283),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_203),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_228),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_228),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_214),
.B(n_224),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_283),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_231),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_231),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_269),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_269),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_282),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_209),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_323),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_217),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_226),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_226),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_378),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_206),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_209),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_282),
.Y(n_464)
);

INVxp33_ASAP7_75t_SL g465 ( 
.A(n_210),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_285),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_285),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_218),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_221),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_292),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_222),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_223),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_378),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_235),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_292),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_209),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_223),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_272),
.B(n_6),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_378),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g480 ( 
.A(n_229),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_223),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_294),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_272),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_272),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_235),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_294),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_312),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_251),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_230),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_312),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_289),
.B(n_7),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_348),
.B(n_7),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_272),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_348),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_353),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_278),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_353),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_375),
.B(n_8),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_415),
.B(n_289),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_415),
.B(n_277),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_416),
.B(n_277),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_375),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_435),
.B(n_477),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_416),
.B(n_227),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_472),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_472),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_417),
.B(n_370),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_412),
.B(n_278),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_417),
.B(n_370),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_472),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_472),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_414),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_401),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_420),
.B(n_278),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_442),
.A2(n_352),
.B(n_273),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_408),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_408),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_409),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_409),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_420),
.B(n_421),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_424),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

XNOR2x2_ASAP7_75t_R g534 ( 
.A(n_427),
.B(n_262),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_410),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_442),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_428),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_411),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_411),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_481),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_481),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_422),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_422),
.B(n_423),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_440),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_440),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_441),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_446),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_451),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_452),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_453),
.B(n_278),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_453),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_454),
.B(n_290),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_454),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_455),
.B(n_205),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_464),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

AND2x2_ASAP7_75t_SL g566 ( 
.A(n_407),
.B(n_352),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_466),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_466),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_448),
.B(n_252),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_470),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_470),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_475),
.B(n_482),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_475),
.B(n_482),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_486),
.B(n_266),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_487),
.Y(n_578)
);

NOR2x1_ASAP7_75t_L g579 ( 
.A(n_487),
.B(n_303),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_490),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_490),
.B(n_310),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_457),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_494),
.B(n_279),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_494),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_520),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_513),
.B(n_465),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_522),
.B(n_478),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_582),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_571),
.B(n_438),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_555),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_555),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_565),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_582),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_507),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_537),
.B(n_456),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_561),
.A2(n_463),
.B1(n_476),
.B2(n_491),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_565),
.B(n_480),
.Y(n_598)
);

BUFx4f_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_499),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_522),
.B(n_491),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_555),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_520),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_557),
.B(n_485),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_565),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_565),
.B(n_462),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_458),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_519),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_557),
.B(n_581),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_581),
.B(n_432),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_519),
.B(n_397),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_520),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_555),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_555),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_519),
.B(n_399),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_520),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_566),
.A2(n_498),
.B1(n_492),
.B2(n_450),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_563),
.B(n_434),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_563),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_563),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_563),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_528),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_574),
.B(n_495),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_561),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_563),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_574),
.B(n_581),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_565),
.B(n_468),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_528),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_563),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_563),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_566),
.A2(n_372),
.B1(n_373),
.B2(n_363),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_565),
.B(n_469),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_528),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_572),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_576),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_528),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_572),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_572),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_565),
.B(n_471),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_566),
.A2(n_450),
.B1(n_399),
.B2(n_413),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_499),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_572),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_572),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_565),
.B(n_495),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_576),
.B(n_489),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_499),
.Y(n_650)
);

AND2x2_ASAP7_75t_SL g651 ( 
.A(n_559),
.B(n_251),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_503),
.A2(n_425),
.B1(n_402),
.B2(n_444),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_583),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_583),
.B(n_443),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_560),
.B(n_497),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_501),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_503),
.A2(n_461),
.B1(n_473),
.B2(n_449),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_501),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_502),
.B(n_497),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_501),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_560),
.B(n_479),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_572),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_504),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_503),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_504),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_506),
.B(n_460),
.C(n_459),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_503),
.A2(n_484),
.B1(n_493),
.B2(n_483),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_504),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_503),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_503),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_572),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_577),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_560),
.B(n_436),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_510),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_549),
.B(n_395),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_577),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_560),
.B(n_398),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_510),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_510),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_536),
.B(n_303),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_577),
.Y(n_682)
);

INVxp33_ASAP7_75t_L g683 ( 
.A(n_502),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_445),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_549),
.B(n_496),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_505),
.B(n_488),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_506),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_577),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_577),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_577),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_577),
.B(n_202),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_577),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_543),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_564),
.B(n_474),
.Y(n_694)
);

INVxp33_ASAP7_75t_L g695 ( 
.A(n_502),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_512),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_559),
.B(n_236),
.C(n_234),
.Y(n_697)
);

BUFx6f_ASAP7_75t_SL g698 ( 
.A(n_505),
.Y(n_698)
);

AND3x2_ASAP7_75t_L g699 ( 
.A(n_534),
.B(n_300),
.C(n_281),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_543),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_512),
.B(n_209),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_545),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_530),
.B(n_300),
.C(n_281),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_543),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_545),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_548),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_508),
.A2(n_244),
.B1(n_246),
.B2(n_242),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_548),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_517),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_517),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_564),
.B(n_350),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_545),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_548),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_564),
.B(n_403),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_551),
.B(n_404),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_552),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_512),
.B(n_377),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_545),
.B(n_211),
.Y(n_718)
);

BUFx6f_ASAP7_75t_SL g719 ( 
.A(n_505),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_521),
.Y(n_720)
);

INVxp33_ASAP7_75t_SL g721 ( 
.A(n_530),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_545),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_552),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_569),
.B(n_213),
.Y(n_724)
);

NOR2x1p5_ASAP7_75t_L g725 ( 
.A(n_544),
.B(n_394),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_505),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_569),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_505),
.A2(n_311),
.B1(n_314),
.B2(n_301),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_521),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_544),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_552),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_505),
.B(n_405),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_687),
.B(n_569),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_585),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_662),
.A2(n_301),
.B1(n_314),
.B2(n_311),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_693),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_588),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_698),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_585),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_585),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_698),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_651),
.A2(n_514),
.B1(n_546),
.B2(n_542),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_693),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_721),
.B(n_569),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_613),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_613),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_613),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_651),
.A2(n_514),
.B1(n_546),
.B2(n_542),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_639),
.B(n_569),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_651),
.A2(n_514),
.B1(n_546),
.B2(n_542),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_610),
.B(n_578),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_617),
.B(n_406),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_730),
.B(n_578),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_702),
.B(n_536),
.Y(n_754)
);

OAI221xp5_ASAP7_75t_L g755 ( 
.A1(n_619),
.A2(n_345),
.B1(n_316),
.B2(n_317),
.C(n_325),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_594),
.B(n_578),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_700),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_653),
.B(n_578),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_653),
.B(n_578),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_600),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_628),
.B(n_515),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_612),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_610),
.B(n_575),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_610),
.B(n_554),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_702),
.B(n_536),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_654),
.B(n_515),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_610),
.B(n_554),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_618),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_593),
.B(n_418),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_630),
.B(n_558),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_704),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_635),
.A2(n_514),
.B1(n_546),
.B2(n_542),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_685),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_605),
.B(n_419),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_630),
.B(n_558),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_618),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_617),
.B(n_575),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_704),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_604),
.B(n_558),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_605),
.B(n_430),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_586),
.A2(n_553),
.B1(n_570),
.B2(n_567),
.Y(n_782)
);

OAI221xp5_ASAP7_75t_L g783 ( 
.A1(n_635),
.A2(n_345),
.B1(n_316),
.B2(n_317),
.C(n_325),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_609),
.B(n_431),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_702),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_618),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_596),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_650),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_701),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_604),
.B(n_567),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_600),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_604),
.B(n_570),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_604),
.B(n_573),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_706),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_701),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_706),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_587),
.A2(n_644),
.B1(n_728),
.B2(n_717),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_650),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_708),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_649),
.B(n_573),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_589),
.B(n_573),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_627),
.B(n_580),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_665),
.A2(n_580),
.B(n_521),
.C(n_525),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_715),
.B(n_580),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_600),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_627),
.B(n_524),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_717),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_708),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_670),
.B(n_547),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_713),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_675),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_702),
.B(n_536),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_665),
.B(n_524),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_698),
.Y(n_814)
);

BUFx8_ASAP7_75t_L g815 ( 
.A(n_698),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_670),
.B(n_536),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_675),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_671),
.B(n_524),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_SL g819 ( 
.A1(n_671),
.A2(n_523),
.B(n_547),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_675),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_670),
.B(n_536),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_696),
.B(n_433),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_683),
.B(n_695),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_608),
.B(n_676),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_726),
.B(n_525),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_601),
.B(n_525),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_726),
.B(n_526),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_608),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_719),
.A2(n_579),
.B1(n_514),
.B2(n_550),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_597),
.B(n_334),
.C(n_329),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_670),
.B(n_547),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_667),
.B(n_527),
.C(n_526),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_L g833 ( 
.A(n_652),
.B(n_527),
.C(n_526),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_659),
.B(n_527),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_713),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_705),
.B(n_536),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_601),
.B(n_529),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_659),
.B(n_529),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_680),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_601),
.B(n_529),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_716),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_716),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_601),
.B(n_531),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_657),
.B(n_514),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_705),
.B(n_536),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_655),
.A2(n_535),
.B(n_538),
.C(n_531),
.Y(n_846)
);

AND2x2_ASAP7_75t_SL g847 ( 
.A(n_598),
.B(n_547),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_723),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_680),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_705),
.B(n_531),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_601),
.B(n_535),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_707),
.B(n_550),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_705),
.B(n_535),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_719),
.A2(n_579),
.B1(n_556),
.B2(n_562),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_611),
.B(n_538),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_712),
.B(n_538),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_611),
.B(n_539),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_SL g858 ( 
.A(n_719),
.B(n_437),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_681),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_719),
.A2(n_550),
.B1(n_562),
.B2(n_556),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_587),
.A2(n_556),
.B1(n_562),
.B2(n_550),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_587),
.A2(n_556),
.B1(n_568),
.B2(n_562),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_686),
.B(n_439),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_686),
.A2(n_584),
.B1(n_568),
.B2(n_338),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_709),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_686),
.B(n_568),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_731),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_709),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_709),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_645),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_SL g871 ( 
.A(n_699),
.B(n_310),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_592),
.B(n_539),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_731),
.Y(n_873)
);

BUFx5_ASAP7_75t_L g874 ( 
.A(n_681),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_611),
.B(n_539),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_611),
.B(n_568),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_SL g877 ( 
.A(n_587),
.B(n_310),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_712),
.B(n_722),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_686),
.A2(n_584),
.B1(n_254),
.B2(n_255),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_645),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_712),
.B(n_584),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_611),
.B(n_584),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_712),
.B(n_540),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_587),
.B(n_678),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_722),
.B(n_540),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_722),
.B(n_540),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_722),
.B(n_540),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_714),
.B(n_259),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_727),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_727),
.Y(n_890)
);

OAI22xp33_ASAP7_75t_L g891 ( 
.A1(n_686),
.A2(n_334),
.B1(n_335),
.B2(n_329),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_697),
.B(n_711),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_727),
.B(n_540),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_732),
.B(n_264),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_822),
.Y(n_895)
);

O2A1O1Ixp5_ASAP7_75t_L g896 ( 
.A1(n_852),
.A2(n_631),
.B(n_643),
.C(n_636),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_767),
.B(n_727),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_760),
.B(n_645),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_767),
.B(n_679),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_754),
.A2(n_599),
.B(n_710),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_736),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_826),
.A2(n_710),
.B(n_729),
.C(n_656),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_758),
.B(n_679),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_760),
.B(n_679),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_824),
.B(n_668),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_734),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_758),
.B(n_607),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_826),
.A2(n_729),
.B1(n_710),
.B2(n_658),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_761),
.B(n_674),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_738),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_837),
.A2(n_729),
.B(n_656),
.C(n_661),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_766),
.A2(n_599),
.B(n_658),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_774),
.A2(n_877),
.B1(n_837),
.B2(n_884),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_761),
.B(n_684),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_775),
.B(n_725),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_739),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_763),
.A2(n_621),
.B(n_694),
.C(n_703),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_797),
.A2(n_661),
.B1(n_666),
.B2(n_664),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_760),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_797),
.A2(n_666),
.B1(n_720),
.B2(n_669),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_743),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_828),
.B(n_718),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_757),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_765),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_766),
.A2(n_812),
.B(n_845),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_749),
.B(n_669),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_733),
.B(n_720),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_772),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_762),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_789),
.B(n_725),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_845),
.A2(n_599),
.B(n_591),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_823),
.B(n_377),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_759),
.B(n_637),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_801),
.B(n_637),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_755),
.A2(n_523),
.B(n_337),
.C(n_342),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_801),
.B(n_640),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_781),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_812),
.A2(n_724),
.B(n_606),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_878),
.A2(n_606),
.B(n_592),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_816),
.A2(n_616),
.B(n_590),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_795),
.B(n_640),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_819),
.A2(n_622),
.B(n_616),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_807),
.B(n_620),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_805),
.A2(n_647),
.B1(n_595),
.B2(n_615),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_760),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_821),
.A2(n_624),
.B(n_622),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_840),
.A2(n_647),
.B1(n_595),
.B2(n_615),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_823),
.B(n_595),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_780),
.B(n_620),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_790),
.B(n_620),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_821),
.A2(n_625),
.B(n_624),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_756),
.A2(n_633),
.B(n_625),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_753),
.A2(n_634),
.B(n_633),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_791),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_738),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_791),
.B(n_595),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_792),
.B(n_626),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_784),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_741),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_741),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_881),
.A2(n_638),
.B(n_634),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_800),
.B(n_626),
.Y(n_962)
);

BUFx12f_ASAP7_75t_L g963 ( 
.A(n_815),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_853),
.A2(n_856),
.B(n_872),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_843),
.A2(n_851),
.B1(n_870),
.B2(n_806),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_870),
.A2(n_647),
.B1(n_614),
.B2(n_623),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_850),
.A2(n_831),
.B(n_809),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_800),
.B(n_626),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_885),
.A2(n_642),
.B(n_638),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_884),
.A2(n_681),
.B1(n_648),
.B2(n_647),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_886),
.A2(n_893),
.B(n_887),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_815),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_787),
.B(n_377),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_778),
.B(n_632),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_850),
.A2(n_646),
.B(n_642),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_793),
.B(n_632),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_744),
.A2(n_632),
.B(n_335),
.C(n_342),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_883),
.A2(n_660),
.B(n_646),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_804),
.B(n_614),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_844),
.B(n_614),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_830),
.A2(n_681),
.B1(n_614),
.B2(n_623),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_779),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_752),
.B(n_377),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_771),
.B(n_603),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_883),
.A2(n_663),
.B(n_660),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_814),
.B(n_681),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_858),
.B(n_310),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_776),
.B(n_603),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_802),
.B(n_681),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_794),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_740),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_813),
.A2(n_673),
.B(n_663),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_818),
.A2(n_677),
.B(n_673),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_847),
.A2(n_682),
.B(n_677),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_834),
.A2(n_838),
.B1(n_796),
.B2(n_808),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_825),
.A2(n_688),
.B(n_682),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_827),
.A2(n_689),
.B(n_688),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_814),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_788),
.A2(n_690),
.B(n_689),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_788),
.A2(n_690),
.B(n_623),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_863),
.B(n_737),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_782),
.B(n_681),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_751),
.B(n_894),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_SL g1004 ( 
.A1(n_803),
.A2(n_692),
.B(n_672),
.C(n_641),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_866),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_791),
.B(n_602),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_894),
.B(n_615),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_798),
.A2(n_623),
.B(n_615),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_791),
.B(n_785),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_798),
.A2(n_641),
.B(n_629),
.Y(n_1010)
);

O2A1O1Ixp5_ASAP7_75t_L g1011 ( 
.A1(n_764),
.A2(n_692),
.B(n_672),
.C(n_641),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_735),
.A2(n_783),
.B1(n_861),
.B2(n_876),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_745),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_785),
.B(n_602),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_768),
.B(n_629),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_773),
.B(n_672),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_773),
.B(n_672),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_891),
.A2(n_369),
.B(n_337),
.C(n_360),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_745),
.Y(n_1019)
);

AOI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_888),
.A2(n_692),
.B(n_691),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_799),
.A2(n_692),
.B1(n_602),
.B2(n_321),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_861),
.B(n_602),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_876),
.B(n_602),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_855),
.A2(n_330),
.B1(n_389),
.B2(n_387),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_880),
.B(n_602),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_746),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_889),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_890),
.A2(n_523),
.B(n_511),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_888),
.B(n_284),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_770),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_880),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_882),
.B(n_540),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_735),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_855),
.A2(n_369),
.B(n_360),
.C(n_374),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_811),
.A2(n_511),
.B(n_500),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_892),
.A2(n_511),
.B(n_500),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_817),
.A2(n_516),
.B(n_500),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_820),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_882),
.B(n_374),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_857),
.B(n_286),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_746),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_810),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_857),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_835),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_833),
.B(n_386),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_820),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_859),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_841),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_874),
.B(n_290),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_874),
.B(n_290),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_839),
.A2(n_518),
.B(n_532),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_879),
.B(n_388),
.C(n_386),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_735),
.B(n_384),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_742),
.B(n_388),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_849),
.A2(n_220),
.B(n_216),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_871),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_842),
.A2(n_392),
.B(n_391),
.C(n_533),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_848),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_875),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_874),
.B(n_290),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_742),
.B(n_748),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_875),
.B(n_390),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_867),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_747),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_748),
.B(n_391),
.Y(n_1065)
);

CKINVDCx10_ASAP7_75t_R g1066 ( 
.A(n_832),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_873),
.B(n_864),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_750),
.B(n_392),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_899),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1059),
.B(n_750),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_895),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_L g1072 ( 
.A(n_1029),
.B(n_305),
.C(n_299),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_937),
.Y(n_1073)
);

AO21x2_ASAP7_75t_L g1074 ( 
.A1(n_942),
.A2(n_862),
.B(n_854),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1061),
.A2(n_869),
.B1(n_868),
.B2(n_865),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_913),
.B(n_860),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_919),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_901),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_SL g1079 ( 
.A1(n_922),
.A2(n_846),
.B(n_869),
.C(n_868),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_963),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1067),
.A2(n_865),
.B1(n_859),
.B2(n_829),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_1029),
.A2(n_1003),
.B(n_1040),
.C(n_922),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1040),
.B(n_747),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1067),
.A2(n_859),
.B1(n_769),
.B2(n_777),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_995),
.A2(n_859),
.B1(n_769),
.B2(n_777),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_1003),
.A2(n_786),
.B(n_533),
.C(n_390),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1001),
.A2(n_1043),
.B1(n_905),
.B2(n_958),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_929),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_974),
.B(n_786),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1012),
.A2(n_354),
.B1(n_313),
.B2(n_315),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_983),
.B(n_874),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_1005),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_921),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_923),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1012),
.A2(n_376),
.B1(n_319),
.B2(n_320),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_909),
.A2(n_533),
.B(n_262),
.C(n_541),
.Y(n_1096)
);

AOI221xp5_ASAP7_75t_L g1097 ( 
.A1(n_1018),
.A2(n_326),
.B1(n_309),
.B2(n_351),
.C(n_331),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_919),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_915),
.A2(n_836),
.B1(n_874),
.B2(n_385),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_972),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_974),
.B(n_836),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_907),
.A2(n_836),
.B(n_874),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_972),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_914),
.B(n_836),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_R g1105 ( 
.A(n_1056),
.B(n_836),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_932),
.B(n_973),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_897),
.B(n_532),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_1020),
.A2(n_533),
.B(n_541),
.C(n_532),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1007),
.A2(n_533),
.B(n_383),
.C(n_346),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_948),
.A2(n_371),
.B1(n_379),
.B2(n_382),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_924),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_955),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_948),
.A2(n_384),
.B1(n_232),
.B2(n_296),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1052),
.A2(n_532),
.B(n_541),
.C(n_384),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_980),
.B(n_541),
.Y(n_1115)
);

NAND2x1p5_ASAP7_75t_L g1116 ( 
.A(n_955),
.B(n_384),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_L g1117 ( 
.A(n_1007),
.B(n_361),
.C(n_291),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1024),
.B(n_233),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1036),
.A2(n_509),
.B(n_290),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1053),
.A2(n_304),
.B1(n_367),
.B2(n_365),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_964),
.A2(n_261),
.B(n_364),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_930),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_928),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_1056),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_930),
.B(n_8),
.Y(n_1125)
);

INVx5_ASAP7_75t_L g1126 ( 
.A(n_986),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_982),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_903),
.A2(n_260),
.B(n_362),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_987),
.B(n_1030),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_990),
.B(n_10),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1066),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_971),
.A2(n_258),
.B(n_359),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_919),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_919),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_984),
.A2(n_257),
.B(n_358),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1042),
.B(n_12),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_965),
.B(n_238),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1034),
.A2(n_12),
.B(n_13),
.C(n_16),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1044),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1048),
.B(n_16),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1058),
.B(n_17),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_945),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_906),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_959),
.B(n_17),
.Y(n_1144)
);

INVxp67_ASAP7_75t_SL g1145 ( 
.A(n_980),
.Y(n_1145)
);

NOR2x1_ASAP7_75t_L g1146 ( 
.A(n_959),
.B(n_240),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_945),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_988),
.A2(n_265),
.B(n_356),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1034),
.A2(n_902),
.B(n_911),
.C(n_1057),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_902),
.A2(n_911),
.B(n_1063),
.C(n_977),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_941),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_925),
.A2(n_295),
.B(n_355),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_918),
.B(n_290),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_945),
.B(n_241),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1054),
.A2(n_306),
.B1(n_349),
.B2(n_347),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_927),
.A2(n_247),
.B(n_341),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1033),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_943),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_986),
.B(n_910),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_R g1160 ( 
.A(n_910),
.B(n_245),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_R g1161 ( 
.A(n_960),
.B(n_248),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_945),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1031),
.B(n_249),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1065),
.A2(n_308),
.B1(n_340),
.B2(n_339),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_917),
.A2(n_267),
.B(n_270),
.C(n_271),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_918),
.B(n_290),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_954),
.B(n_275),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_920),
.A2(n_1068),
.B1(n_908),
.B2(n_935),
.Y(n_1168)
);

AND3x1_ASAP7_75t_SL g1169 ( 
.A(n_1027),
.B(n_24),
.C(n_26),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1027),
.B(n_276),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_960),
.B(n_280),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_SL g1172 ( 
.A(n_935),
.B(n_1045),
.C(n_1039),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_989),
.A2(n_287),
.B(n_336),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_954),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1004),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_920),
.B(n_28),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_954),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_954),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_979),
.B(n_288),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1004),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_926),
.B(n_30),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_934),
.B(n_33),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_936),
.B(n_37),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_998),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_998),
.B(n_1023),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_916),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_979),
.B(n_293),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1047),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_938),
.A2(n_318),
.B(n_333),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_898),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1047),
.B(n_90),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1002),
.A2(n_322),
.B(n_327),
.C(n_328),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1032),
.B(n_290),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_962),
.B(n_45),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_900),
.A2(n_88),
.B(n_102),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_1016),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1038),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1062),
.B(n_49),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_912),
.A2(n_104),
.B(n_107),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1038),
.B(n_49),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1046),
.B(n_50),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1055),
.B(n_54),
.C(n_55),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1046),
.B(n_290),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_968),
.A2(n_1000),
.B(n_999),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1028),
.A2(n_509),
.B(n_110),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_991),
.Y(n_1206)
);

BUFx5_ASAP7_75t_L g1207 ( 
.A(n_1049),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_991),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_969),
.A2(n_140),
.B(n_190),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_SL g1210 ( 
.A1(n_1015),
.A2(n_54),
.B(n_57),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_961),
.A2(n_132),
.B(n_177),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1013),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_994),
.B(n_63),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1009),
.B(n_509),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_898),
.B(n_509),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_904),
.B(n_64),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_904),
.B(n_65),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1017),
.B(n_976),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1022),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1082),
.A2(n_957),
.B1(n_950),
.B2(n_949),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1105),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_1103),
.B(n_1006),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1078),
.Y(n_1223)
);

OAI22x1_ASAP7_75t_L g1224 ( 
.A1(n_1087),
.A2(n_970),
.B1(n_981),
.B2(n_956),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1093),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1106),
.B(n_1019),
.Y(n_1226)
);

BUFx8_ASAP7_75t_L g1227 ( 
.A(n_1131),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1102),
.A2(n_931),
.B(n_1014),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1150),
.A2(n_1011),
.B(n_896),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1094),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1124),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1145),
.B(n_1070),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1092),
.B(n_1019),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1088),
.Y(n_1234)
);

AOI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1152),
.A2(n_951),
.B1(n_946),
.B2(n_940),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1090),
.A2(n_1021),
.B1(n_947),
.B2(n_933),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1205),
.A2(n_997),
.B(n_996),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1168),
.A2(n_944),
.B1(n_966),
.B2(n_967),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1104),
.A2(n_993),
.B(n_992),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_1088),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1204),
.A2(n_952),
.B(n_953),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1195),
.A2(n_1060),
.B(n_1050),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1149),
.A2(n_1008),
.B(n_1010),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1083),
.A2(n_978),
.B(n_985),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1080),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1101),
.A2(n_939),
.B(n_975),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1118),
.B(n_956),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1092),
.B(n_1064),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_L g1249 ( 
.A(n_1100),
.B(n_1006),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1152),
.A2(n_1037),
.B(n_1035),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1199),
.A2(n_1050),
.B(n_1049),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1085),
.A2(n_1064),
.A3(n_1026),
.B(n_1041),
.Y(n_1252)
);

AOI31xp67_ASAP7_75t_L g1253 ( 
.A1(n_1193),
.A2(n_1014),
.A3(n_1025),
.B(n_1041),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1085),
.A2(n_1025),
.B(n_1026),
.Y(n_1254)
);

INVx3_ASAP7_75t_SL g1255 ( 
.A(n_1144),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1073),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1069),
.A2(n_1051),
.B(n_120),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1071),
.B(n_66),
.Y(n_1258)
);

NOR2xp67_ASAP7_75t_L g1259 ( 
.A(n_1129),
.B(n_1170),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1151),
.B(n_66),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1144),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1084),
.A2(n_1107),
.B(n_1081),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1116),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1122),
.B(n_69),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1125),
.B(n_71),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_1079),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_1266)
);

AOI221x1_ASAP7_75t_L g1267 ( 
.A1(n_1090),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.C(n_76),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1111),
.B(n_77),
.Y(n_1268)
);

INVx3_ASAP7_75t_SL g1269 ( 
.A(n_1216),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1077),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1160),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1084),
.A2(n_131),
.B(n_111),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1107),
.A2(n_1081),
.B(n_1089),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1110),
.A2(n_78),
.B(n_118),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1126),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1076),
.A2(n_126),
.B(n_128),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1158),
.B(n_509),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1120),
.B(n_509),
.C(n_141),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1126),
.B(n_129),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_SL g1280 ( 
.A1(n_1165),
.A2(n_142),
.B(n_144),
.C(n_146),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1168),
.A2(n_158),
.B(n_509),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1075),
.A2(n_1108),
.B(n_1209),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1123),
.B(n_1127),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1075),
.A2(n_1211),
.B(n_1096),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1210),
.A2(n_1086),
.B(n_1185),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1137),
.A2(n_1115),
.B(n_1074),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1179),
.B(n_1187),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1196),
.A2(n_1172),
.B(n_1166),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1077),
.Y(n_1289)
);

O2A1O1Ixp5_ASAP7_75t_L g1290 ( 
.A1(n_1213),
.A2(n_1091),
.B(n_1154),
.C(n_1167),
.Y(n_1290)
);

AOI221x1_ASAP7_75t_L g1291 ( 
.A1(n_1095),
.A2(n_1176),
.B1(n_1202),
.B2(n_1198),
.C(n_1194),
.Y(n_1291)
);

AO22x1_ASAP7_75t_L g1292 ( 
.A1(n_1095),
.A2(n_1216),
.B1(n_1217),
.B2(n_1146),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1171),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1139),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1217),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1157),
.B(n_1208),
.Y(n_1296)
);

OAI21xp33_ASAP7_75t_L g1297 ( 
.A1(n_1113),
.A2(n_1183),
.B(n_1182),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1130),
.A2(n_1141),
.B1(n_1136),
.B2(n_1140),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1214),
.A2(n_1153),
.B(n_1191),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1115),
.A2(n_1074),
.B(n_1181),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1097),
.B(n_1197),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1109),
.A2(n_1175),
.B(n_1180),
.C(n_1138),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1116),
.B(n_1190),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1161),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1077),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1173),
.A2(n_1117),
.B(n_1132),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1098),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1192),
.A2(n_1201),
.B(n_1200),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1099),
.A2(n_1218),
.B(n_1114),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1143),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1186),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1203),
.A2(n_1163),
.B(n_1219),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1212),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1169),
.A2(n_1219),
.B1(n_1159),
.B2(n_1164),
.Y(n_1314)
);

AOI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1155),
.A2(n_1121),
.B1(n_1189),
.B2(n_1156),
.C(n_1128),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1135),
.A2(n_1148),
.B(n_1184),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1126),
.A2(n_1191),
.B1(n_1112),
.B2(n_1215),
.Y(n_1317)
);

AO32x2_ASAP7_75t_L g1318 ( 
.A1(n_1162),
.A2(n_1177),
.A3(n_1207),
.B1(n_1206),
.B2(n_1178),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1133),
.A2(n_1134),
.A3(n_1177),
.B(n_1162),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1174),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1207),
.A2(n_1206),
.A3(n_1215),
.B(n_1142),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1098),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1112),
.B(n_1206),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1188),
.A2(n_1098),
.B(n_1142),
.C(n_1147),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1142),
.B(n_1147),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1188),
.A2(n_1215),
.B(n_1147),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1207),
.A2(n_1082),
.B(n_899),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1207),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1082),
.B(n_1145),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1078),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1082),
.B(n_913),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1119),
.A2(n_1205),
.B(n_1204),
.Y(n_1332)
);

CKINVDCx6p67_ASAP7_75t_R g1333 ( 
.A(n_1080),
.Y(n_1333)
);

BUFx10_ASAP7_75t_L g1334 ( 
.A(n_1144),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1092),
.B(n_824),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1082),
.A2(n_774),
.B(n_1029),
.C(n_1072),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_SL g1337 ( 
.A(n_1080),
.B(n_752),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1077),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1082),
.B(n_1145),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1082),
.A2(n_899),
.B1(n_1067),
.B2(n_1061),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1085),
.A2(n_1075),
.A3(n_1084),
.B(n_1168),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1085),
.A2(n_1075),
.A3(n_1084),
.B(n_1168),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1124),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1088),
.Y(n_1344)
);

AO32x2_ASAP7_75t_L g1345 ( 
.A1(n_1090),
.A2(n_1033),
.A3(n_1095),
.B1(n_1168),
.B2(n_1075),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1078),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_SL g1347 ( 
.A1(n_1082),
.A2(n_1150),
.B(n_1149),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1082),
.B(n_824),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1082),
.B(n_824),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1124),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_SL g1351 ( 
.A1(n_1082),
.A2(n_899),
.B(n_1079),
.C(n_897),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1082),
.A2(n_911),
.B(n_902),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1078),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1082),
.B(n_774),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1078),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1082),
.B(n_824),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1078),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1092),
.B(n_824),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1085),
.A2(n_1075),
.A3(n_1084),
.B(n_1168),
.Y(n_1359)
);

AND2x6_ASAP7_75t_L g1360 ( 
.A(n_1159),
.B(n_986),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1082),
.A2(n_899),
.B(n_907),
.Y(n_1361)
);

AOI221x1_ASAP7_75t_L g1362 ( 
.A1(n_1090),
.A2(n_1095),
.B1(n_1029),
.B2(n_1168),
.C(n_1152),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1082),
.A2(n_899),
.B(n_907),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1119),
.A2(n_1205),
.B(n_1204),
.Y(n_1364)
);

CKINVDCx8_ASAP7_75t_R g1365 ( 
.A(n_1073),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1105),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1082),
.A2(n_899),
.B(n_907),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1090),
.A2(n_654),
.B1(n_657),
.B2(n_822),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1196),
.A2(n_1096),
.B(n_1172),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_SL g1370 ( 
.A1(n_1082),
.A2(n_899),
.B(n_1079),
.C(n_897),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1082),
.B(n_824),
.Y(n_1371)
);

AOI21xp33_ASAP7_75t_L g1372 ( 
.A1(n_1082),
.A2(n_1029),
.B(n_1168),
.Y(n_1372)
);

NOR2xp67_ASAP7_75t_SL g1373 ( 
.A(n_1080),
.B(n_752),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1082),
.A2(n_899),
.B(n_907),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1350),
.Y(n_1375)
);

BUFx4f_ASAP7_75t_SL g1376 ( 
.A(n_1227),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1283),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1372),
.B2(n_1331),
.Y(n_1378)
);

BUFx4_ASAP7_75t_SL g1379 ( 
.A(n_1245),
.Y(n_1379)
);

NAND2x1p5_ASAP7_75t_L g1380 ( 
.A(n_1275),
.B(n_1279),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1354),
.B(n_1335),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1223),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1225),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1293),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1230),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1240),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1294),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1358),
.B(n_1232),
.Y(n_1388)
);

INVx6_ASAP7_75t_L g1389 ( 
.A(n_1334),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1330),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1227),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1297),
.A2(n_1298),
.B1(n_1348),
.B2(n_1371),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1233),
.B(n_1232),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1297),
.A2(n_1298),
.B1(n_1356),
.B2(n_1349),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1307),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1336),
.A2(n_1340),
.B1(n_1329),
.B2(n_1339),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1333),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1256),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1346),
.Y(n_1399)
);

INVx6_ASAP7_75t_L g1400 ( 
.A(n_1334),
.Y(n_1400)
);

BUFx4f_ASAP7_75t_SL g1401 ( 
.A(n_1263),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1340),
.A2(n_1347),
.B1(n_1308),
.B2(n_1329),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1353),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1355),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1240),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1305),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1339),
.A2(n_1247),
.B1(n_1314),
.B2(n_1274),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1357),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1310),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1343),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1274),
.A2(n_1373),
.B1(n_1337),
.B2(n_1314),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1308),
.A2(n_1259),
.B1(n_1269),
.B2(n_1295),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1304),
.A2(n_1362),
.B1(n_1309),
.B2(n_1352),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1301),
.A2(n_1309),
.B1(n_1352),
.B2(n_1265),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1311),
.Y(n_1415)
);

OAI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1267),
.A2(n_1255),
.B1(n_1268),
.B2(n_1291),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1226),
.A2(n_1248),
.B1(n_1278),
.B2(n_1313),
.Y(n_1417)
);

BUFx4f_ASAP7_75t_SL g1418 ( 
.A(n_1234),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1292),
.A2(n_1271),
.B1(n_1303),
.B2(n_1231),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1221),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1270),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1302),
.A2(n_1236),
.B1(n_1367),
.B2(n_1363),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1365),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1366),
.Y(n_1424)
);

OAI22x1_ASAP7_75t_L g1425 ( 
.A1(n_1261),
.A2(n_1320),
.B1(n_1264),
.B2(n_1296),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1236),
.A2(n_1374),
.B1(n_1361),
.B2(n_1281),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1260),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1262),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1344),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1258),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1220),
.A2(n_1238),
.B1(n_1327),
.B2(n_1222),
.Y(n_1431)
);

INVx8_ASAP7_75t_L g1432 ( 
.A(n_1360),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1222),
.A2(n_1277),
.B1(n_1279),
.B2(n_1345),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1318),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1220),
.A2(n_1238),
.B1(n_1222),
.B2(n_1315),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1270),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1270),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1345),
.A2(n_1288),
.B1(n_1369),
.B2(n_1273),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1345),
.A2(n_1288),
.B1(n_1369),
.B2(n_1229),
.Y(n_1439)
);

BUFx8_ASAP7_75t_L g1440 ( 
.A(n_1289),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1249),
.B(n_1360),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1319),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1252),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1289),
.Y(n_1444)
);

BUFx4f_ASAP7_75t_SL g1445 ( 
.A(n_1289),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1338),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1360),
.B(n_1322),
.Y(n_1447)
);

BUFx4f_ASAP7_75t_SL g1448 ( 
.A(n_1338),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1229),
.A2(n_1300),
.B1(n_1286),
.B2(n_1272),
.Y(n_1449)
);

BUFx4_ASAP7_75t_R g1450 ( 
.A(n_1328),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1360),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1325),
.Y(n_1452)
);

AO22x1_ASAP7_75t_L g1453 ( 
.A1(n_1275),
.A2(n_1323),
.B1(n_1322),
.B2(n_1338),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_SL g1454 ( 
.A(n_1224),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1326),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1317),
.A2(n_1257),
.B1(n_1312),
.B2(n_1276),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1299),
.Y(n_1457)
);

INVx6_ASAP7_75t_L g1458 ( 
.A(n_1324),
.Y(n_1458)
);

BUFx2_ASAP7_75t_SL g1459 ( 
.A(n_1316),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1321),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1290),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1266),
.Y(n_1462)
);

BUFx4f_ASAP7_75t_SL g1463 ( 
.A(n_1253),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1243),
.A2(n_1254),
.B1(n_1244),
.B2(n_1235),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1306),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1341),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1285),
.Y(n_1467)
);

BUFx2_ASAP7_75t_R g1468 ( 
.A(n_1351),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1341),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1243),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1342),
.B(n_1359),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1342),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1359),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1239),
.B2(n_1359),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1241),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1251),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1284),
.A2(n_1250),
.B1(n_1282),
.B2(n_1239),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1370),
.B(n_1246),
.Y(n_1478)
);

BUFx10_ASAP7_75t_L g1479 ( 
.A(n_1280),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1250),
.A2(n_1228),
.B(n_1242),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1237),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1237),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1332),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1364),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1350),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1287),
.A2(n_1029),
.B1(n_774),
.B2(n_877),
.Y(n_1486)
);

OAI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1362),
.A2(n_1287),
.B1(n_877),
.B2(n_1274),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1256),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1307),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1287),
.A2(n_1053),
.B1(n_735),
.B2(n_877),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1307),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1287),
.A2(n_1082),
.B1(n_1354),
.B2(n_1029),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1256),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1335),
.B(n_1358),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1287),
.A2(n_1053),
.B1(n_735),
.B2(n_877),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1256),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1283),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1283),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1240),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1307),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1287),
.A2(n_1082),
.B1(n_1354),
.B2(n_1029),
.Y(n_1506)
);

CKINVDCx6p67_ASAP7_75t_R g1507 ( 
.A(n_1350),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1362),
.A2(n_1287),
.B1(n_877),
.B2(n_1274),
.Y(n_1508)
);

AO22x1_ASAP7_75t_L g1509 ( 
.A1(n_1287),
.A2(n_1053),
.B1(n_1304),
.B2(n_830),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1305),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1334),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1283),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1287),
.A2(n_1053),
.B1(n_735),
.B2(n_877),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1227),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1283),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1287),
.A2(n_1368),
.B1(n_1053),
.B2(n_735),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1256),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1256),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1283),
.Y(n_1522)
);

OAI22x1_ASAP7_75t_L g1523 ( 
.A1(n_1287),
.A2(n_1314),
.B1(n_1269),
.B2(n_1087),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1483),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1443),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1443),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1470),
.Y(n_1528)
);

AO21x1_ASAP7_75t_SL g1529 ( 
.A1(n_1402),
.A2(n_1478),
.B(n_1394),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1452),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1388),
.B(n_1377),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_L g1532 ( 
.A(n_1493),
.B(n_1506),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1472),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1471),
.B(n_1466),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1472),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1396),
.B(n_1422),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1384),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1442),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1426),
.A2(n_1482),
.B(n_1481),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1469),
.B(n_1382),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1463),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1428),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1428),
.Y(n_1543)
);

CKINVDCx14_ASAP7_75t_R g1544 ( 
.A(n_1375),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1463),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1393),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1409),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1383),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1415),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1385),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1387),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1501),
.B(n_1502),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1390),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1469),
.B(n_1457),
.Y(n_1554)
);

INVx4_ASAP7_75t_R g1555 ( 
.A(n_1454),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1399),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1403),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1404),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1408),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1485),
.B(n_1423),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1434),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1487),
.A2(n_1508),
.B(n_1474),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1457),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1467),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1474),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1484),
.A2(n_1480),
.B(n_1456),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1402),
.B(n_1439),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1438),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1496),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1486),
.A2(n_1407),
.B1(n_1508),
.B2(n_1487),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1438),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1439),
.B(n_1414),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1378),
.A2(n_1414),
.B1(n_1497),
.B2(n_1498),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1431),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1451),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1513),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1440),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_SL g1578 ( 
.A(n_1516),
.Y(n_1578)
);

INVxp33_ASAP7_75t_L g1579 ( 
.A(n_1419),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1440),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1476),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1507),
.B(n_1420),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1420),
.B(n_1424),
.Y(n_1583)
);

BUFx2_ASAP7_75t_SL g1584 ( 
.A(n_1386),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1435),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1517),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1381),
.B(n_1413),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1522),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1392),
.B(n_1394),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1379),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1405),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1465),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1424),
.B(n_1410),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1405),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1376),
.B(n_1418),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1413),
.B(n_1392),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1477),
.B(n_1427),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1378),
.A2(n_1417),
.B(n_1411),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1460),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1445),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1456),
.A2(n_1417),
.B(n_1462),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1464),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1475),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1475),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1433),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1458),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1459),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1458),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1430),
.B(n_1425),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1432),
.B(n_1380),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1491),
.A2(n_1515),
.B1(n_1499),
.B2(n_1511),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1477),
.B(n_1412),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1450),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1412),
.B(n_1509),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1449),
.A2(n_1380),
.B(n_1416),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1461),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1461),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1491),
.A2(n_1515),
.B1(n_1499),
.B2(n_1511),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1461),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1458),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1455),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1416),
.B(n_1523),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1450),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1449),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1447),
.A2(n_1441),
.B(n_1479),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1453),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1489),
.A2(n_1498),
.B1(n_1497),
.B2(n_1495),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1479),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1489),
.A2(n_1514),
.B1(n_1503),
.B2(n_1495),
.C(n_1519),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1444),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1468),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1503),
.A2(n_1518),
.B1(n_1519),
.B2(n_1514),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1421),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1437),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1432),
.B(n_1504),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1446),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_L g1637 ( 
.A(n_1518),
.B(n_1406),
.C(n_1510),
.D(n_1490),
.Y(n_1637)
);

INVx5_ASAP7_75t_SL g1638 ( 
.A(n_1610),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1597),
.B(n_1510),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1597),
.B(n_1406),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1524),
.B(n_1436),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1532),
.A2(n_1492),
.B(n_1505),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1546),
.B(n_1398),
.Y(n_1643)
);

AOI21xp33_ASAP7_75t_L g1644 ( 
.A1(n_1596),
.A2(n_1395),
.B(n_1520),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1598),
.A2(n_1536),
.B(n_1589),
.C(n_1624),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1540),
.B(n_1554),
.Y(n_1646)
);

A2O1A1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1536),
.A2(n_1521),
.B(n_1488),
.C(n_1500),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1565),
.B(n_1494),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1570),
.A2(n_1379),
.B(n_1448),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1550),
.B(n_1376),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1540),
.B(n_1448),
.Y(n_1651)
);

A2O1A1Ixp33_ASAP7_75t_L g1652 ( 
.A1(n_1573),
.A2(n_1445),
.B(n_1512),
.C(n_1400),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1567),
.B(n_1389),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1573),
.A2(n_1389),
.B(n_1512),
.C(n_1400),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1565),
.B(n_1429),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1524),
.B(n_1389),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1558),
.B(n_1418),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1625),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1576),
.B(n_1397),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1628),
.B(n_1400),
.Y(n_1660)
);

AO32x2_ASAP7_75t_L g1661 ( 
.A1(n_1591),
.A2(n_1391),
.A3(n_1401),
.B1(n_1594),
.B2(n_1572),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1534),
.B(n_1401),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1615),
.A2(n_1596),
.B(n_1601),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1625),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1567),
.A2(n_1614),
.B(n_1622),
.C(n_1632),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1585),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1586),
.B(n_1530),
.Y(n_1668)
);

NOR2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1577),
.B(n_1580),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1585),
.B(n_1588),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1554),
.B(n_1607),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1588),
.B(n_1587),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1556),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1556),
.B(n_1557),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1592),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1569),
.B(n_1583),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1601),
.A2(n_1614),
.B(n_1622),
.Y(n_1678)
);

AND2x4_ASAP7_75t_SL g1679 ( 
.A(n_1613),
.B(n_1623),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1630),
.B(n_1621),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1611),
.A2(n_1618),
.B1(n_1627),
.B2(n_1629),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1630),
.B(n_1621),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1562),
.B(n_1574),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1592),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1612),
.B(n_1636),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1587),
.B(n_1531),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1557),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1566),
.A2(n_1539),
.B(n_1602),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1574),
.A2(n_1619),
.B(n_1617),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_SL g1691 ( 
.A1(n_1590),
.A2(n_1595),
.B(n_1593),
.C(n_1616),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_SL g1692 ( 
.A1(n_1619),
.A2(n_1545),
.B(n_1541),
.C(n_1560),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1554),
.B(n_1541),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1572),
.A2(n_1600),
.B1(n_1620),
.B2(n_1631),
.Y(n_1694)
);

AND2x2_ASAP7_75t_SL g1695 ( 
.A(n_1568),
.B(n_1571),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1562),
.A2(n_1637),
.B1(n_1620),
.B2(n_1608),
.Y(n_1696)
);

INVx11_ASAP7_75t_L g1697 ( 
.A(n_1544),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1579),
.A2(n_1568),
.B(n_1571),
.C(n_1605),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1559),
.B(n_1542),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1561),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1566),
.A2(n_1542),
.B(n_1543),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1543),
.B(n_1561),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1553),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1552),
.B(n_1547),
.Y(n_1704)
);

OAI21xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1635),
.A2(n_1610),
.B(n_1528),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1547),
.B(n_1549),
.Y(n_1706)
);

O2A1O1Ixp33_ASAP7_75t_SL g1707 ( 
.A1(n_1545),
.A2(n_1631),
.B(n_1528),
.C(n_1555),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1563),
.B(n_1529),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1634),
.B(n_1633),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1538),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1609),
.A2(n_1605),
.B(n_1606),
.C(n_1608),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1533),
.A2(n_1535),
.B1(n_1609),
.B2(n_1526),
.C(n_1527),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1700),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1681),
.A2(n_1606),
.B1(n_1610),
.B2(n_1626),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1710),
.Y(n_1715)
);

AND2x2_ASAP7_75t_SL g1716 ( 
.A(n_1695),
.B(n_1575),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1676),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1688),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1702),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1699),
.B(n_1535),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1708),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1604),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1689),
.B(n_1603),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1658),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1705),
.B(n_1594),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1699),
.B(n_1533),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1674),
.Y(n_1727)
);

BUFx12f_ASAP7_75t_L g1728 ( 
.A(n_1669),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1665),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1684),
.B(n_1526),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1638),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1646),
.B(n_1672),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1673),
.B(n_1527),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1668),
.B(n_1564),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1646),
.B(n_1564),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1667),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1670),
.B(n_1525),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1663),
.A2(n_1599),
.B1(n_1626),
.B2(n_1525),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1667),
.B(n_1584),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1672),
.B(n_1581),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1701),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1679),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1675),
.B(n_1581),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1697),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1693),
.B(n_1671),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1639),
.B(n_1584),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1712),
.B(n_1686),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1658),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1658),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1664),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1657),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1706),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1664),
.Y(n_1754)
);

INVxp67_ASAP7_75t_SL g1755 ( 
.A(n_1717),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1716),
.A2(n_1683),
.B1(n_1666),
.B2(n_1695),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1738),
.A2(n_1666),
.B1(n_1645),
.B2(n_1683),
.C(n_1698),
.Y(n_1757)
);

INVx4_ASAP7_75t_L g1758 ( 
.A(n_1728),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1722),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1715),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1715),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1732),
.B(n_1639),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1733),
.B(n_1687),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1736),
.B(n_1640),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1745),
.B(n_1640),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1741),
.A2(n_1647),
.B(n_1696),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1715),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1730),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1732),
.B(n_1721),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1736),
.B(n_1680),
.Y(n_1771)
);

OAI211xp5_ASAP7_75t_L g1772 ( 
.A1(n_1741),
.A2(n_1642),
.B(n_1691),
.C(n_1649),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1728),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1730),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1713),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1721),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1728),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1747),
.B(n_1682),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1721),
.B(n_1677),
.Y(n_1779)
);

INVx4_ASAP7_75t_L g1780 ( 
.A(n_1744),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1721),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1734),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1747),
.B(n_1648),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1722),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1733),
.B(n_1643),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1713),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1734),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1745),
.B(n_1651),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1733),
.B(n_1720),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1722),
.Y(n_1790)
);

NAND2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1716),
.B(n_1731),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1718),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1745),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1718),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1727),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1740),
.B(n_1648),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1720),
.B(n_1709),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1723),
.Y(n_1798)
);

AOI222xp33_ASAP7_75t_L g1799 ( 
.A1(n_1738),
.A2(n_1678),
.B1(n_1711),
.B2(n_1694),
.C1(n_1654),
.C2(n_1655),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1726),
.B(n_1704),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1727),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1753),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1744),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1716),
.A2(n_1655),
.B1(n_1644),
.B2(n_1653),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1745),
.B(n_1651),
.Y(n_1805)
);

NAND4xp25_ASAP7_75t_L g1806 ( 
.A(n_1752),
.B(n_1650),
.C(n_1659),
.D(n_1647),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1725),
.B(n_1651),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1753),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1743),
.B(n_1690),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1749),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1752),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1749),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1731),
.Y(n_1813)
);

INVxp67_ASAP7_75t_SL g1814 ( 
.A(n_1748),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1807),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1798),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1781),
.B(n_1724),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1769),
.B(n_1737),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1810),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_1737),
.Y(n_1820)
);

INVx4_ASAP7_75t_L g1821 ( 
.A(n_1758),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1781),
.B(n_1724),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1793),
.B(n_1770),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1761),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1807),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1793),
.B(n_1724),
.Y(n_1826)
);

NOR2x1_ASAP7_75t_L g1827 ( 
.A(n_1758),
.B(n_1641),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1789),
.B(n_1764),
.Y(n_1828)
);

INVxp67_ASAP7_75t_SL g1829 ( 
.A(n_1767),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1812),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_L g1831 ( 
.A(n_1772),
.B(n_1754),
.C(n_1751),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1795),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1755),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1802),
.B(n_1726),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1801),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1789),
.B(n_1734),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1775),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1808),
.B(n_1743),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1798),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1786),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1792),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1770),
.B(n_1750),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1757),
.A2(n_1716),
.B(n_1725),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1759),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1759),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1794),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1776),
.B(n_1750),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1764),
.B(n_1729),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1784),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1760),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1803),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1762),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1782),
.B(n_1743),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_R g1854 ( 
.A(n_1803),
.B(n_1578),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1780),
.B(n_1773),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1787),
.B(n_1719),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1768),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1776),
.B(n_1750),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1776),
.B(n_1735),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1797),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1785),
.B(n_1729),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1816),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1824),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1837),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1851),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_SL g1866 ( 
.A(n_1843),
.B(n_1825),
.C(n_1815),
.Y(n_1866)
);

INVxp33_ASAP7_75t_L g1867 ( 
.A(n_1854),
.Y(n_1867)
);

OR2x6_ASAP7_75t_L g1868 ( 
.A(n_1843),
.B(n_1758),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1829),
.A2(n_1756),
.B1(n_1799),
.B2(n_1714),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1815),
.B(n_1766),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1816),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1825),
.B(n_1766),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1829),
.B(n_1783),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1823),
.B(n_1766),
.Y(n_1874)
);

CKINVDCx16_ASAP7_75t_R g1875 ( 
.A(n_1851),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1828),
.B(n_1785),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1819),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1823),
.B(n_1788),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1837),
.Y(n_1879)
);

NAND2x1_ASAP7_75t_SL g1880 ( 
.A(n_1827),
.B(n_1807),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1819),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1830),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1823),
.B(n_1788),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1816),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1827),
.B(n_1788),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1830),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1828),
.B(n_1800),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_L g1888 ( 
.A(n_1821),
.B(n_1806),
.C(n_1777),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1832),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1842),
.B(n_1805),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1860),
.B(n_1811),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1839),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1839),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1842),
.B(n_1805),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1836),
.B(n_1800),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1836),
.B(n_1797),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1832),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1839),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1860),
.B(n_1809),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1851),
.B(n_1773),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1835),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1835),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1840),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1818),
.B(n_1778),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1818),
.B(n_1765),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1844),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1820),
.B(n_1771),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1844),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1876),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1873),
.B(n_1833),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1864),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1873),
.B(n_1833),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1863),
.B(n_1820),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1887),
.B(n_1876),
.Y(n_1914)
);

INVx2_ASAP7_75t_SL g1915 ( 
.A(n_1880),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_SL g1916 ( 
.A(n_1875),
.B(n_1780),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1875),
.B(n_1831),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1887),
.B(n_1834),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1865),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1895),
.B(n_1834),
.Y(n_1920)
);

AND2x2_ASAP7_75t_SL g1921 ( 
.A(n_1888),
.B(n_1821),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1865),
.B(n_1904),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1879),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1877),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1891),
.B(n_1840),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1895),
.B(n_1841),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1867),
.B(n_1780),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1877),
.Y(n_1928)
);

NOR2xp67_ASAP7_75t_L g1929 ( 
.A(n_1866),
.B(n_1831),
.Y(n_1929)
);

INVx1_ASAP7_75t_SL g1930 ( 
.A(n_1880),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1874),
.B(n_1878),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1896),
.B(n_1861),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1874),
.B(n_1821),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1881),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1885),
.B(n_1878),
.Y(n_1935)
);

NAND2xp33_ASAP7_75t_R g1936 ( 
.A(n_1868),
.B(n_1777),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1883),
.B(n_1821),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1883),
.B(n_1842),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1885),
.B(n_1855),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1896),
.B(n_1841),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1881),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1905),
.B(n_1899),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1869),
.B(n_1846),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1882),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1885),
.B(n_1859),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1905),
.B(n_1861),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1885),
.B(n_1859),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1919),
.B(n_1900),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1914),
.Y(n_1949)
);

AOI32xp33_ASAP7_75t_L g1950 ( 
.A1(n_1943),
.A2(n_1868),
.A3(n_1870),
.B1(n_1872),
.B2(n_1869),
.Y(n_1950)
);

NAND3xp33_ASAP7_75t_L g1951 ( 
.A(n_1929),
.B(n_1868),
.C(n_1882),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1916),
.B(n_1868),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1914),
.B(n_1942),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1909),
.B(n_1907),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1915),
.B(n_1930),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1917),
.A2(n_1868),
.B1(n_1915),
.B2(n_1935),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1909),
.A2(n_1908),
.B1(n_1862),
.B2(n_1906),
.Y(n_1957)
);

A2O1A1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1921),
.A2(n_1910),
.B(n_1912),
.C(n_1942),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1924),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1931),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1939),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1921),
.A2(n_1889),
.B(n_1886),
.Y(n_1962)
);

AOI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1922),
.A2(n_1886),
.B1(n_1889),
.B2(n_1897),
.C(n_1903),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1911),
.B(n_1907),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1923),
.B(n_1899),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1936),
.A2(n_1908),
.B1(n_1906),
.B2(n_1893),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1939),
.A2(n_1872),
.B(n_1870),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1931),
.B(n_1937),
.Y(n_1968)
);

AOI222xp33_ASAP7_75t_L g1969 ( 
.A1(n_1923),
.A2(n_1908),
.B1(n_1906),
.B2(n_1862),
.C1(n_1871),
.C2(n_1884),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1924),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1935),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1935),
.A2(n_1890),
.B1(n_1894),
.B2(n_1791),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1927),
.B(n_1890),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1941),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1913),
.A2(n_1925),
.B(n_1945),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1926),
.A2(n_1862),
.B1(n_1898),
.B2(n_1893),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1953),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1949),
.B(n_1932),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1959),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1970),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1968),
.B(n_1937),
.Y(n_1981)
);

CKINVDCx16_ASAP7_75t_R g1982 ( 
.A(n_1961),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_SL g1983 ( 
.A1(n_1951),
.A2(n_1580),
.B1(n_1577),
.B2(n_1941),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1958),
.A2(n_1933),
.B(n_1928),
.C(n_1934),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1974),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1971),
.B(n_1933),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1960),
.B(n_1938),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1973),
.B(n_1938),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1950),
.A2(n_1962),
.B(n_1966),
.C(n_1948),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1954),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1965),
.Y(n_1991)
);

AOI211xp5_ASAP7_75t_L g1992 ( 
.A1(n_1956),
.A2(n_1944),
.B(n_1932),
.C(n_1946),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1964),
.Y(n_1993)
);

NOR2x1_ASAP7_75t_L g1994 ( 
.A(n_1955),
.B(n_1945),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1967),
.A2(n_1946),
.B1(n_1918),
.B2(n_1920),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1975),
.B(n_1940),
.Y(n_1996)
);

NOR2x1p5_ASAP7_75t_SL g1997 ( 
.A(n_1962),
.B(n_1871),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1963),
.B(n_1969),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1969),
.B(n_1918),
.Y(n_1999)
);

OAI21xp33_ASAP7_75t_SL g2000 ( 
.A1(n_1994),
.A2(n_1952),
.B(n_1947),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1982),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1988),
.B(n_1894),
.Y(n_2002)
);

AOI21xp33_ASAP7_75t_L g2003 ( 
.A1(n_1998),
.A2(n_1957),
.B(n_1976),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1990),
.B(n_1920),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1977),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1999),
.A2(n_1871),
.B1(n_1884),
.B2(n_1892),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1990),
.B(n_1947),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_SL g2008 ( 
.A(n_1989),
.B(n_1600),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1978),
.Y(n_2009)
);

AOI211x1_ASAP7_75t_SL g2010 ( 
.A1(n_1989),
.A2(n_1995),
.B(n_1996),
.C(n_1992),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1990),
.B(n_1897),
.Y(n_2011)
);

AOI211xp5_ASAP7_75t_L g2012 ( 
.A1(n_1983),
.A2(n_1972),
.B(n_1707),
.C(n_1691),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1988),
.B(n_1987),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1987),
.B(n_1903),
.Y(n_2014)
);

OAI21xp33_ASAP7_75t_L g2015 ( 
.A1(n_2008),
.A2(n_1997),
.B(n_1986),
.Y(n_2015)
);

NOR3x1_ASAP7_75t_L g2016 ( 
.A(n_2013),
.B(n_1991),
.C(n_1984),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_2001),
.Y(n_2017)
);

OAI211xp5_ASAP7_75t_L g2018 ( 
.A1(n_2000),
.A2(n_1993),
.B(n_1986),
.C(n_1979),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2014),
.Y(n_2019)
);

O2A1O1Ixp5_ASAP7_75t_L g2020 ( 
.A1(n_2003),
.A2(n_1985),
.B(n_1980),
.C(n_1981),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2011),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2004),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_2008),
.B(n_2002),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2007),
.Y(n_2024)
);

OAI211xp5_ASAP7_75t_L g2025 ( 
.A1(n_2010),
.A2(n_1981),
.B(n_1902),
.C(n_1901),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_2009),
.A2(n_1902),
.B1(n_1901),
.B2(n_1846),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_2006),
.A2(n_1892),
.B(n_1884),
.Y(n_2027)
);

OAI21xp33_ASAP7_75t_L g2028 ( 
.A1(n_2005),
.A2(n_1822),
.B(n_1817),
.Y(n_2028)
);

OAI211xp5_ASAP7_75t_SL g2029 ( 
.A1(n_2012),
.A2(n_1853),
.B(n_1838),
.C(n_1739),
.Y(n_2029)
);

AOI221xp5_ASAP7_75t_L g2030 ( 
.A1(n_2015),
.A2(n_1898),
.B1(n_1893),
.B2(n_1892),
.C(n_1857),
.Y(n_2030)
);

OAI211xp5_ASAP7_75t_L g2031 ( 
.A1(n_2018),
.A2(n_1817),
.B(n_1822),
.C(n_1826),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2017),
.Y(n_2032)
);

NAND4xp25_ASAP7_75t_L g2033 ( 
.A(n_2016),
.B(n_1739),
.C(n_1826),
.D(n_1817),
.Y(n_2033)
);

OAI311xp33_ASAP7_75t_L g2034 ( 
.A1(n_2028),
.A2(n_1804),
.A3(n_1714),
.B1(n_1826),
.C1(n_1856),
.Y(n_2034)
);

O2A1O1Ixp33_ASAP7_75t_L g2035 ( 
.A1(n_2020),
.A2(n_2025),
.B(n_2022),
.C(n_2021),
.Y(n_2035)
);

NAND4xp75_ASAP7_75t_L g2036 ( 
.A(n_2023),
.B(n_1898),
.C(n_1662),
.D(n_1822),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2019),
.Y(n_2037)
);

OAI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_2024),
.A2(n_1857),
.B1(n_1838),
.B2(n_1856),
.Y(n_2038)
);

OAI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_2027),
.A2(n_1858),
.B(n_1847),
.Y(n_2039)
);

AOI211x1_ASAP7_75t_L g2040 ( 
.A1(n_2031),
.A2(n_2026),
.B(n_2029),
.C(n_1685),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2035),
.A2(n_2029),
.B1(n_1850),
.B2(n_1852),
.C(n_1849),
.Y(n_2041)
);

OAI211xp5_ASAP7_75t_L g2042 ( 
.A1(n_2032),
.A2(n_2037),
.B(n_2033),
.C(n_2030),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2036),
.B(n_1847),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2034),
.A2(n_1850),
.B1(n_1852),
.B2(n_1845),
.C(n_1849),
.Y(n_2044)
);

OAI211xp5_ASAP7_75t_L g2045 ( 
.A1(n_2039),
.A2(n_1858),
.B(n_1847),
.C(n_1814),
.Y(n_2045)
);

AOI211xp5_ASAP7_75t_L g2046 ( 
.A1(n_2038),
.A2(n_1707),
.B(n_1662),
.C(n_1692),
.Y(n_2046)
);

NAND3xp33_ASAP7_75t_L g2047 ( 
.A(n_2035),
.B(n_1858),
.C(n_1754),
.Y(n_2047)
);

NOR2xp67_ASAP7_75t_L g2048 ( 
.A(n_2033),
.B(n_1859),
.Y(n_2048)
);

OAI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_2035),
.A2(n_1849),
.B(n_1845),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_2048),
.B(n_2043),
.Y(n_2050)
);

OR2x6_ASAP7_75t_L g2051 ( 
.A(n_2042),
.B(n_1844),
.Y(n_2051)
);

NOR2x1_ASAP7_75t_L g2052 ( 
.A(n_2047),
.B(n_1779),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_2049),
.B(n_1779),
.Y(n_2053)
);

NAND4xp75_ASAP7_75t_L g2054 ( 
.A(n_2040),
.B(n_1660),
.C(n_1656),
.D(n_1746),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2045),
.Y(n_2055)
);

AOI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_2050),
.A2(n_2041),
.B1(n_2044),
.B2(n_2046),
.C(n_1845),
.Y(n_2056)
);

NAND3x1_ASAP7_75t_L g2057 ( 
.A(n_2055),
.B(n_1853),
.C(n_1763),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_2051),
.B(n_1748),
.C(n_1751),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_2052),
.B(n_1805),
.Y(n_2059)
);

AO22x2_ASAP7_75t_L g2060 ( 
.A1(n_2059),
.A2(n_2054),
.B1(n_2053),
.B2(n_2051),
.Y(n_2060)
);

XNOR2xp5_ASAP7_75t_L g2061 ( 
.A(n_2057),
.B(n_1804),
.Y(n_2061)
);

OAI22x1_ASAP7_75t_L g2062 ( 
.A1(n_2061),
.A2(n_2058),
.B1(n_2060),
.B2(n_2056),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_2062),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2062),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2063),
.B(n_1784),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2064),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2066),
.Y(n_2067)
);

OAI21x1_ASAP7_75t_L g2068 ( 
.A1(n_2065),
.A2(n_1848),
.B(n_1791),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2067),
.Y(n_2069)
);

OAI222xp33_ASAP7_75t_L g2070 ( 
.A1(n_2069),
.A2(n_2068),
.B1(n_1848),
.B2(n_1790),
.C1(n_1796),
.C2(n_1660),
.Y(n_2070)
);

XNOR2xp5_ASAP7_75t_L g2071 ( 
.A(n_2070),
.B(n_1599),
.Y(n_2071)
);

OAI221xp5_ASAP7_75t_R g2072 ( 
.A1(n_2071),
.A2(n_1555),
.B1(n_1692),
.B2(n_1742),
.C(n_1661),
.Y(n_2072)
);

AOI211xp5_ASAP7_75t_L g2073 ( 
.A1(n_2072),
.A2(n_1813),
.B(n_1746),
.C(n_1652),
.Y(n_2073)
);


endmodule