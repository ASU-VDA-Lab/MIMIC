module fake_jpeg_3340_n_360 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_51),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_48),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_20),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_19),
.A2(n_28),
.B1(n_26),
.B2(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_79),
.B1(n_80),
.B2(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_68),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_67),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_32),
.B(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_23),
.B(n_7),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_74),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_19),
.B1(n_29),
.B2(n_26),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_88),
.B1(n_104),
.B2(n_111),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_45),
.A2(n_44),
.B1(n_41),
.B2(n_40),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_44),
.B1(n_31),
.B2(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_31),
.B1(n_25),
.B2(n_39),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_41),
.B(n_40),
.C(n_39),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_111),
.B(n_96),
.C(n_85),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_59),
.A2(n_17),
.B1(n_31),
.B2(n_38),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_38),
.B1(n_30),
.B2(n_24),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_64),
.B1(n_69),
.B2(n_60),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_24),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_117),
.B(n_126),
.Y(n_180)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_118),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_146),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_121),
.Y(n_171)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_140),
.Y(n_161)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_30),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_127),
.B(n_129),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_134),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_144),
.B(n_145),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_137),
.B(n_138),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_49),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_63),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_149),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_48),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_150),
.Y(n_166)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_158),
.B1(n_89),
.B2(n_56),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_17),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_58),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_154),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_79),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_156),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_82),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_64),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_22),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_100),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_54),
.C(n_90),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_179),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_107),
.C(n_97),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_107),
.B1(n_76),
.B2(n_72),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_181),
.B1(n_189),
.B2(n_144),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_98),
.C(n_78),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_119),
.A2(n_66),
.B1(n_62),
.B2(n_95),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_120),
.A2(n_95),
.B1(n_89),
.B2(n_22),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_137),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_203),
.Y(n_231)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_127),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_199),
.Y(n_222)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_155),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_191),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_205),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_116),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_161),
.B(n_146),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_131),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_182),
.B(n_160),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_160),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_208),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_130),
.B1(n_145),
.B2(n_149),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_214),
.B1(n_215),
.B2(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_118),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_166),
.B(n_158),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_168),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_130),
.B1(n_125),
.B2(n_128),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_171),
.B(n_175),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_236),
.B(n_192),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_181),
.B1(n_176),
.B2(n_167),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_224),
.B1(n_229),
.B2(n_215),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_167),
.B1(n_171),
.B2(n_163),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_235),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_167),
.B1(n_189),
.B2(n_162),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_230),
.A2(n_209),
.B1(n_204),
.B2(n_207),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_179),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_210),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_184),
.B(n_192),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_202),
.C(n_198),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_240),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_232),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_224),
.B(n_233),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_253),
.B(n_216),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_213),
.B1(n_214),
.B2(n_196),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_223),
.B1(n_219),
.B2(n_228),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_193),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_249),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_252),
.B1(n_256),
.B2(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_234),
.C(n_235),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_208),
.Y(n_252)
);

XOR2x1_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_173),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_188),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_206),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_172),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_220),
.A2(n_197),
.B1(n_194),
.B2(n_178),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_237),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_265),
.Y(n_280)
);

AO22x2_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_221),
.B1(n_229),
.B2(n_227),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_272),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_270),
.B1(n_172),
.B2(n_170),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_249),
.B1(n_223),
.B2(n_257),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_225),
.B(n_183),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_148),
.B(n_135),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_225),
.C(n_121),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_121),
.C(n_173),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_278),
.C(n_246),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_239),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_250),
.C(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_238),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_286),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_284),
.C(n_296),
.Y(n_298)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_238),
.C(n_240),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_266),
.B1(n_259),
.B2(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_291),
.B1(n_292),
.B2(n_275),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_244),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_289),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_170),
.B1(n_186),
.B2(n_143),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_186),
.B1(n_164),
.B2(n_151),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_164),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_293),
.B(n_295),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_271),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_122),
.B1(n_134),
.B2(n_133),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_134),
.C(n_133),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_303),
.B1(n_10),
.B2(n_12),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_280),
.C(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_262),
.B1(n_261),
.B2(n_269),
.Y(n_303)
);

OA21x2_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_272),
.B(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_268),
.Y(n_305)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_280),
.B(n_262),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_313),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_262),
.B(n_139),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_37),
.B(n_1),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_132),
.C(n_22),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_292),
.C(n_291),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_298),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_300),
.A2(n_295),
.B(n_12),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_321),
.B(n_305),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_319),
.B1(n_306),
.B2(n_311),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_22),
.B1(n_10),
.B2(n_16),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_7),
.C(n_16),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_5),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_37),
.B1(n_33),
.B2(n_7),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_324),
.A2(n_322),
.B1(n_325),
.B2(n_320),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_325),
.Y(n_330)
);

INVx11_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_298),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_328),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_332),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_307),
.C(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_334),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_335),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_319),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_314),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_326),
.A2(n_308),
.B(n_324),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_4),
.B(n_12),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_332),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_345),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_330),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_346),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_330),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_348),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_309),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_349),
.A2(n_342),
.B1(n_343),
.B2(n_336),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_4),
.Y(n_355)
);

O2A1O1Ixp33_ASAP7_75t_SL g354 ( 
.A1(n_351),
.A2(n_4),
.B(n_15),
.C(n_2),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_354),
.A2(n_355),
.B(n_356),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_352),
.A2(n_0),
.B(n_1),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_352),
.C(n_350),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_0),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_359),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_360)
);


endmodule