module real_jpeg_6797_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_323;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_0),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_0),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_0),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_0),
.B(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_0),
.B(n_482),
.Y(n_481)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_2),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_2),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_2),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_2),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_2),
.B(n_262),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_2),
.B(n_405),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_3),
.B(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_3),
.A2(n_254),
.B(n_256),
.Y(n_253)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_3),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_3),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_3),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_3),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_3),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_3),
.B(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_4),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_5),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_5),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_5),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_5),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_5),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_5),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_5),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_5),
.B(n_428),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_6),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_6),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_6),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_6),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_6),
.B(n_277),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_6),
.B(n_262),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_6),
.B(n_410),
.Y(n_409)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_8),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_10),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_10),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_10),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_10),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_203),
.Y(n_202)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_12),
.Y(n_93)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_12),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_12),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_12),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_13),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_13),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_13),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_13),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_13),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_13),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_13),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_13),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_14),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_14),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_14),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_14),
.B(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_15),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_464),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_221),
.B(n_461),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_177),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_SL g461 ( 
.A1(n_19),
.A2(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_136),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_20),
.B(n_136),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_21),
.B(n_102),
.C(n_116),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.C(n_82),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_22),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_48),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_23),
.B(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_26),
.B(n_33),
.C(n_37),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_28),
.A2(n_33),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_28),
.B(n_202),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_28),
.A2(n_33),
.B1(n_201),
.B2(n_202),
.Y(n_429)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_39),
.C(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_34),
.A2(n_37),
.B1(n_110),
.B2(n_113),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_34),
.B(n_276),
.C(n_280),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_34),
.A2(n_37),
.B1(n_280),
.B2(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_37),
.B(n_105),
.C(n_110),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_38),
.B(n_48),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_39),
.A2(n_120),
.B1(n_121),
.B2(n_125),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_39),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_39),
.A2(n_44),
.B1(n_125),
.B2(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_43),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_43),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_43),
.Y(n_343)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_44),
.Y(n_147)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_47),
.Y(n_212)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_47),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_47),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_55),
.Y(n_246)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_56),
.Y(n_374)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_58),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_61),
.C(n_64),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_58),
.B(n_191),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_62),
.B(n_190),
.C(n_194),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_63),
.A2(n_64),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_65),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_66),
.A2(n_82),
.B1(n_83),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_76),
.C(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_71),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_73),
.B(n_86),
.C(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_73),
.A2(n_80),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.C(n_98),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_84),
.A2(n_85),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.C(n_92),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_86),
.A2(n_92),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_86),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_86),
.A2(n_160),
.B1(n_166),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_86),
.A2(n_160),
.B1(n_386),
.B2(n_388),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_86),
.B(n_388),
.Y(n_430)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_87),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_88),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_88),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_88),
.B(n_243),
.C(n_247),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_88),
.A2(n_162),
.B1(n_243),
.B2(n_313),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_92),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_94),
.A2(n_98),
.B1(n_99),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_98),
.A2(n_99),
.B1(n_169),
.B2(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_99),
.B(n_165),
.C(n_169),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.C(n_115),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_105),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_104),
.B(n_231),
.C(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_104),
.A2(n_105),
.B1(n_231),
.B2(n_232),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_105),
.B(n_122),
.C(n_125),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_110),
.Y(n_113)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_112),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_115),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_118),
.B(n_119),
.C(n_126),
.Y(n_468)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_122),
.A2(n_123),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_122),
.A2(n_123),
.B1(n_149),
.B2(n_475),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_123),
.B(n_201),
.C(n_207),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_127),
.B(n_131),
.C(n_134),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_129),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_137),
.B(n_140),
.CI(n_142),
.CON(n_220),
.SN(n_220)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_164),
.C(n_173),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_158),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_144),
.B(n_148),
.Y(n_297)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_156),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_149),
.Y(n_475)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_156),
.Y(n_198)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_155),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_158),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_173),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_166),
.B(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_166),
.A2(n_188),
.B1(n_284),
.B2(n_285),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_167),
.Y(n_379)
);

INVx8_ASAP7_75t_L g403 ( 
.A(n_167),
.Y(n_403)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_168),
.Y(n_412)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_220),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_178),
.B(n_220),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_179),
.B(n_181),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_183),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_199),
.C(n_217),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_184),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.C(n_197),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_189),
.B(n_197),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_199),
.B(n_217),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_209),
.C(n_213),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_200),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_201),
.A2(n_202),
.B1(n_207),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_206),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_206),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_207),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_212),
.Y(n_346)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_220),
.Y(n_487)
);

AOI221xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_358),
.B1(n_454),
.B2(n_459),
.C(n_460),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_301),
.C(n_305),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_223),
.A2(n_455),
.B(n_458),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_294),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_224),
.B(n_294),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_268),
.C(n_271),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_225),
.B(n_268),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_251),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_226),
.B(n_252),
.C(n_265),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_241),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_228),
.B(n_242),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_230),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_235),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_236),
.B(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g387 ( 
.A(n_240),
.Y(n_387)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_247),
.B(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_265),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_261),
.C(n_263),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_253),
.A2(n_256),
.B(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_263),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_288),
.C(n_292),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.C(n_282),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_273),
.B(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_275),
.A2(n_282),
.B1(n_283),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_275),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_276),
.B(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_292),
.Y(n_309)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_298),
.C(n_300),
.Y(n_302)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_301),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_302),
.B(n_303),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_331),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_306),
.A2(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_329),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_307),
.B(n_329),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.C(n_327),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_327),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.C(n_318),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_314),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_316),
.B(n_392),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.C(n_324),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_319),
.A2(n_320),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_356),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_332),
.B(n_356),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.C(n_353),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_333),
.B(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_335),
.B(n_353),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.C(n_351),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_336),
.B(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_339),
.A2(n_351),
.B1(n_352),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_339),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_344),
.C(n_347),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_340),
.A2(n_341),
.B1(n_347),
.B2(n_348),
.Y(n_434)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_344),
.B(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_449),
.B(n_453),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_436),
.B(n_448),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_423),
.B(n_435),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_397),
.B(n_422),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_389),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_389),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_375),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_364),
.B(n_376),
.C(n_385),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_370),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_371),
.C(n_372),
.Y(n_432)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_385),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_380),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_380),
.Y(n_390)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_386),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.C(n_395),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_390),
.B(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_395),
.B1(n_396),
.B2(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_391),
.Y(n_420)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_416),
.B(n_421),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_408),
.B(n_415),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_407),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_407),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_404),
.Y(n_417)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_413),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_418),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_425),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_431),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_426),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_432),
.C(n_433),
.Y(n_447)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_429),
.CI(n_430),
.CON(n_426),
.SN(n_426)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_447),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_447),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_444),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_441),
.C(n_444),
.Y(n_450)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_442),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_450),
.B(n_451),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_484),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_467),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_476),
.B1(n_477),
.B2(n_483),
.Y(n_471)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_472),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_479),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_481),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);


endmodule