module fake_ariane_593_n_466 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_466);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_466;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_373;
wire n_299;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_261;
wire n_220;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_387;
wire n_406;
wire n_139;
wire n_349;
wire n_391;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_143;
wire n_152;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_331;
wire n_401;
wire n_267;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_465;
wire n_247;
wire n_240;
wire n_369;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_390;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_464;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_182;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_460;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_351;
wire n_393;
wire n_359;
wire n_155;

INVx2_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_8),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_11),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_74),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_46),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_19),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_39),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_45),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_89),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_34),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_51),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_78),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_61),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_42),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_65),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_69),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_33),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_37),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_83),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_11),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_86),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_59),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_85),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_60),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_70),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_7),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_77),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_90),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_30),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_41),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_64),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_55),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_134),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_63),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_112),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_72),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_81),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_48),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_10),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_53),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_82),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_43),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_110),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_14),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_1),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_123),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_3),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_54),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_22),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_67),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_126),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_84),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_13),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_52),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_88),
.Y(n_213)
);

INVxp33_ASAP7_75t_SL g214 ( 
.A(n_66),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_47),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_49),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_93),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_76),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_125),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_79),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_50),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_9),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_105),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_98),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_102),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_56),
.Y(n_231)
);

BUFx8_ASAP7_75t_SL g232 ( 
.A(n_116),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_71),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_27),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_99),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_113),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_0),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_145),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_1),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_2),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_3),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_151),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_4),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_5),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_159),
.B(n_6),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_164),
.B(n_7),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_167),
.B(n_8),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_141),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_166),
.B(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_169),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_135),
.B(n_10),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_12),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_170),
.B(n_12),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_31),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_185),
.B(n_15),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_172),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_195),
.B(n_16),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_232),
.Y(n_269)
);

BUFx8_ASAP7_75t_SL g270 ( 
.A(n_138),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_139),
.B(n_17),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_147),
.B(n_18),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_153),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_210),
.B(n_18),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_174),
.B(n_20),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_144),
.Y(n_284)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_155),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_171),
.B(n_21),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_136),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_226),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_190),
.Y(n_290)
);

AO22x2_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_180),
.B1(n_199),
.B2(n_143),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_213),
.B1(n_227),
.B2(n_156),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_270),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_238),
.A2(n_214),
.B1(n_140),
.B2(n_142),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_256),
.B(n_233),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_R g296 ( 
.A1(n_240),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_R g298 ( 
.A1(n_245),
.A2(n_261),
.B1(n_248),
.B2(n_244),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_247),
.A2(n_149),
.B1(n_150),
.B2(n_148),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_152),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_253),
.A2(n_231),
.B1(n_229),
.B2(n_228),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_281),
.A2(n_221),
.B1(n_220),
.B2(n_219),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g306 ( 
.A1(n_277),
.A2(n_217),
.B1(n_216),
.B2(n_215),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_254),
.A2(n_212),
.B1(n_208),
.B2(n_207),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

AO22x2_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

AO22x2_ASAP7_75t_L g316 ( 
.A1(n_275),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_316)
);

AO22x2_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_241),
.B1(n_242),
.B2(n_255),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g318 ( 
.A1(n_241),
.A2(n_28),
.B1(n_29),
.B2(n_157),
.Y(n_318)
);

AO22x2_ASAP7_75t_L g319 ( 
.A1(n_242),
.A2(n_28),
.B1(n_29),
.B2(n_157),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_R g320 ( 
.A1(n_255),
.A2(n_157),
.B1(n_197),
.B2(n_194),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_246),
.B(n_154),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_249),
.A2(n_198),
.B1(n_191),
.B2(n_189),
.Y(n_322)
);

AO22x2_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_157),
.B1(n_187),
.B2(n_186),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_251),
.A2(n_188),
.B1(n_184),
.B2(n_182),
.Y(n_324)
);

OR2x6_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_272),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_278),
.A2(n_179),
.B1(n_178),
.B2(n_177),
.Y(n_326)
);

AO22x2_ASAP7_75t_L g327 ( 
.A1(n_260),
.A2(n_157),
.B1(n_176),
.B2(n_175),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g328 ( 
.A1(n_258),
.A2(n_173),
.B1(n_168),
.B2(n_165),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_162),
.B1(n_161),
.B2(n_158),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_297),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_276),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_292),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_252),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_267),
.Y(n_339)
);

OR2x6_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_266),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_295),
.B(n_259),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_302),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_280),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_273),
.Y(n_349)
);

NAND2x1p5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_323),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_291),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_289),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_306),
.B(n_289),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_239),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_320),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_279),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_R g363 ( 
.A(n_298),
.B(n_32),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_285),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_334),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_328),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_332),
.B(n_300),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_294),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_336),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_343),
.B(n_322),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_346),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_324),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_290),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_338),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_362),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_363),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_296),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_263),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_352),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_359),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_35),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_36),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_348),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_361),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_384),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_353),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_374),
.B(n_335),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_367),
.B(n_355),
.Y(n_399)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_383),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_365),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_371),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_38),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_400),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_402),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_404),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_387),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_410),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_399),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_369),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_395),
.A2(n_394),
.B1(n_385),
.B2(n_382),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_420),
.A2(n_368),
.B1(n_419),
.B2(n_375),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_419),
.A2(n_408),
.B1(n_373),
.B2(n_390),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_416),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_417),
.A2(n_373),
.B1(n_390),
.B2(n_391),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_398),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_421),
.A2(n_390),
.B1(n_391),
.B2(n_378),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_427),
.A2(n_423),
.B1(n_425),
.B2(n_422),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_401),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_429),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_412),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_418),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_431),
.A2(n_413),
.B1(n_414),
.B2(n_389),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_434),
.A2(n_393),
.B1(n_392),
.B2(n_379),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_433),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_430),
.A2(n_377),
.B1(n_409),
.B2(n_407),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_438),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_265),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_436),
.C(n_437),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_440),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_442),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_444),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_443),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_443),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_445),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_446),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_447),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_449),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_451),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_452),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_453),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_454),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_455),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_456),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

AO22x2_ASAP7_75t_L g459 ( 
.A1(n_458),
.A2(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_459),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_460),
.A2(n_133),
.B1(n_96),
.B2(n_97),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_461),
.Y(n_462)
);

OA22x2_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_463),
.Y(n_464)
);

AOI221xp5_ASAP7_75t_L g465 ( 
.A1(n_464),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.C(n_118),
.Y(n_465)
);

AOI211xp5_ASAP7_75t_L g466 ( 
.A1(n_465),
.A2(n_119),
.B(n_120),
.C(n_122),
.Y(n_466)
);


endmodule