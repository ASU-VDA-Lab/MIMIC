module fake_jpeg_7609_n_209 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_1),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_1),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_17),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_3),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_4),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_23),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_11),
.C(n_14),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_13),
.B(n_14),
.C(n_12),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_16),
.B1(n_26),
.B2(n_30),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_65),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_66),
.B(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_59),
.B1(n_16),
.B2(n_15),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_5),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_16),
.B1(n_22),
.B2(n_28),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_75),
.B1(n_81),
.B2(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_22),
.B1(n_27),
.B2(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_17),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_68),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_27),
.B1(n_25),
.B2(n_20),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_92),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_20),
.B1(n_25),
.B2(n_38),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_95),
.B1(n_60),
.B2(n_63),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_46),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_38),
.B1(n_39),
.B2(n_31),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_48),
.C(n_38),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_103),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_70),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_116),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_52),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_117),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_31),
.C(n_20),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_79),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_131),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_76),
.B1(n_66),
.B2(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_140),
.B1(n_114),
.B2(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_80),
.B(n_78),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_112),
.B(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_92),
.B1(n_83),
.B2(n_89),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_105),
.B1(n_111),
.B2(n_99),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_6),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_139),
.A2(n_106),
.B(n_117),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_83),
.B1(n_78),
.B2(n_88),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_6),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_126),
.B(n_132),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_136),
.B1(n_126),
.B2(n_124),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_116),
.C(n_100),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_110),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_107),
.C(n_106),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_135),
.B(n_140),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_156),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_134),
.B(n_128),
.C(n_125),
.D(n_139),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_157),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_69),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_128),
.B(n_122),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_101),
.B1(n_79),
.B2(n_98),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_127),
.B1(n_137),
.B2(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_172),
.B(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_149),
.C(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_177),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_151),
.C(n_147),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_133),
.B1(n_156),
.B2(n_128),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_169),
.B1(n_172),
.B2(n_165),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_122),
.C(n_152),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_163),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_139),
.C(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_185),
.A2(n_186),
.B(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_166),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_170),
.B(n_164),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_184),
.B(n_31),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_190),
.B1(n_179),
.B2(n_178),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_163),
.B1(n_166),
.B2(n_12),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_188),
.B(n_190),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_192),
.A2(n_10),
.B1(n_13),
.B2(n_31),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_198),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_10),
.C(n_8),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_198),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_193),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_205),
.B(n_7),
.CI(n_8),
.CON(n_206),
.SN(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_206),
.A2(n_9),
.B1(n_203),
.B2(n_207),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_206),
.Y(n_209)
);


endmodule