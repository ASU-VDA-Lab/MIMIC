module fake_jpeg_13364_n_537 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_537);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_21),
.B(n_0),
.CON(n_56),
.SN(n_56)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_56),
.B(n_0),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_57),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_31),
.B(n_8),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_71),
.Y(n_107)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_31),
.A2(n_7),
.B(n_16),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_31),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_99),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_101),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_39),
.B(n_44),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_20),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_62),
.A2(n_44),
.B1(n_48),
.B2(n_43),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_151),
.B1(n_20),
.B2(n_25),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_67),
.A2(n_43),
.B1(n_44),
.B2(n_35),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_26),
.B(n_40),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_65),
.A2(n_85),
.B1(n_100),
.B2(n_99),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_135),
.A2(n_139),
.B1(n_55),
.B2(n_53),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_51),
.B1(n_41),
.B2(n_35),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_158),
.B1(n_25),
.B2(n_50),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_66),
.A2(n_51),
.B1(n_35),
.B2(n_27),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_57),
.B(n_46),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_154),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_40),
.B(n_26),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_56),
.A2(n_44),
.B1(n_20),
.B2(n_41),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_86),
.B(n_20),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_20),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_70),
.B(n_46),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_73),
.A2(n_51),
.B1(n_41),
.B2(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_75),
.B(n_46),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_159),
.B(n_20),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_96),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_162),
.B(n_163),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_161),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_164),
.A2(n_189),
.B1(n_166),
.B2(n_173),
.Y(n_231)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_25),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_166),
.B(n_196),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_194),
.B1(n_215),
.B2(n_120),
.Y(n_218)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_169),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_173),
.Y(n_227)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_174),
.B(n_181),
.Y(n_241)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_19),
.B1(n_52),
.B2(n_38),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_96),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_184),
.Y(n_265)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_130),
.A2(n_38),
.B1(n_24),
.B2(n_23),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_139),
.A2(n_103),
.B1(n_97),
.B2(n_94),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_50),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_20),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_208),
.C(n_134),
.Y(n_250)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_143),
.B(n_86),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_201),
.B(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_207),
.Y(n_247)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_203),
.Y(n_223)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_205),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_136),
.A2(n_92),
.B1(n_90),
.B2(n_78),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_158),
.B1(n_58),
.B2(n_60),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_113),
.B(n_50),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_127),
.B(n_89),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_212),
.Y(n_251)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_151),
.A2(n_19),
.B1(n_52),
.B2(n_23),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_49),
.B1(n_37),
.B2(n_28),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_146),
.Y(n_255)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_216),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_218),
.A2(n_257),
.B1(n_263),
.B2(n_264),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_112),
.B1(n_116),
.B2(n_141),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_225),
.A2(n_243),
.B1(n_249),
.B2(n_258),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_231),
.B(n_232),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_160),
.B1(n_141),
.B2(n_116),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_170),
.A2(n_160),
.B1(n_104),
.B2(n_119),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_227),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_215),
.A2(n_93),
.B1(n_79),
.B2(n_61),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_209),
.A2(n_206),
.B1(n_173),
.B2(n_198),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_196),
.A2(n_134),
.B(n_80),
.C(n_77),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_260),
.A2(n_244),
.B(n_182),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_206),
.A2(n_126),
.B1(n_115),
.B2(n_122),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_179),
.A2(n_122),
.B1(n_119),
.B2(n_108),
.Y(n_264)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_209),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_289),
.C(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_242),
.B(n_198),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_184),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_206),
.B1(n_197),
.B2(n_191),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_273),
.A2(n_226),
.B1(n_246),
.B2(n_261),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_248),
.A2(n_199),
.B1(n_172),
.B2(n_211),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_274),
.A2(n_304),
.B(n_269),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx11_ASAP7_75t_L g326 ( 
.A(n_275),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_204),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_276),
.B(n_284),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_165),
.B1(n_180),
.B2(n_175),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_277),
.A2(n_287),
.B1(n_293),
.B2(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_171),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_281),
.Y(n_318)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_252),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_185),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_202),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_195),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_292),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_249),
.A2(n_186),
.B1(n_214),
.B2(n_207),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_224),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_227),
.B(n_200),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_243),
.A2(n_106),
.B1(n_212),
.B2(n_41),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_227),
.B(n_183),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_309),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_221),
.B(n_205),
.C(n_216),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_248),
.A2(n_51),
.B1(n_27),
.B2(n_168),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_221),
.B(n_26),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_128),
.B1(n_49),
.B2(n_37),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_305),
.B1(n_34),
.B2(n_24),
.Y(n_325)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_260),
.A2(n_263),
.B1(n_232),
.B2(n_238),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_302),
.A2(n_220),
.B1(n_254),
.B2(n_230),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_238),
.A2(n_40),
.B(n_23),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_251),
.B(n_36),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_264),
.A2(n_203),
.B1(n_188),
.B2(n_128),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_232),
.A2(n_28),
.B1(n_49),
.B2(n_37),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_306),
.Y(n_341)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_229),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_307),
.B(n_245),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_232),
.A2(n_52),
.B1(n_38),
.B2(n_36),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_19),
.B1(n_24),
.B2(n_34),
.Y(n_342)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_222),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_228),
.B(n_28),
.C(n_34),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_0),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_349),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_323),
.B1(n_325),
.B2(n_332),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_283),
.A2(n_254),
.B1(n_234),
.B2(n_228),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_322),
.A2(n_327),
.B1(n_335),
.B2(n_342),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_295),
.A2(n_234),
.B1(n_233),
.B2(n_237),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_324),
.A2(n_329),
.B(n_303),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_283),
.A2(n_233),
.B1(n_237),
.B2(n_229),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_285),
.A2(n_262),
.B(n_256),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_281),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_1),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_271),
.A2(n_256),
.B(n_226),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_331),
.A2(n_345),
.B(n_292),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_236),
.B1(n_259),
.B2(n_222),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_279),
.A2(n_261),
.B1(n_259),
.B2(n_236),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_300),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_337),
.A2(n_344),
.B1(n_348),
.B2(n_274),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_240),
.B1(n_223),
.B2(n_246),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_343),
.A2(n_322),
.B1(n_327),
.B2(n_293),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_282),
.A2(n_246),
.B1(n_226),
.B2(n_239),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_294),
.A2(n_239),
.B(n_262),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_284),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_346),
.B(n_267),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_298),
.A2(n_245),
.B1(n_36),
.B2(n_12),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_310),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_334),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_354),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_349),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_328),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_355),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_315),
.A2(n_270),
.B1(n_286),
.B2(n_308),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_356),
.A2(n_360),
.B1(n_368),
.B2(n_384),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_268),
.C(n_289),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_367),
.C(n_369),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_330),
.A2(n_278),
.B1(n_282),
.B2(n_304),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_361),
.A2(n_343),
.B1(n_312),
.B2(n_336),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_288),
.Y(n_363)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_366),
.Y(n_401)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_314),
.B(n_272),
.C(n_276),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_317),
.A2(n_306),
.B1(n_301),
.B2(n_290),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_296),
.C(n_277),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_291),
.C(n_307),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_373),
.C(n_381),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_375),
.B(n_377),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_305),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_376),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_317),
.B(n_287),
.C(n_309),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_324),
.Y(n_408)
);

NAND2x1_ASAP7_75t_SL g375 ( 
.A(n_329),
.B(n_266),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_297),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_378),
.A2(n_321),
.B1(n_323),
.B2(n_344),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_313),
.B(n_12),
.C(n_17),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_379),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_383),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_275),
.C(n_2),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_351),
.A2(n_11),
.B(n_16),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_321),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_319),
.B(n_12),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_387),
.C(n_350),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_1),
.C(n_2),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_392),
.B1(n_402),
.B2(n_405),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_389),
.A2(n_13),
.B1(n_16),
.B2(n_6),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_347),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_397),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_357),
.A2(n_378),
.B1(n_372),
.B2(n_363),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_347),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_387),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_337),
.B1(n_329),
.B2(n_331),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_328),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_408),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_369),
.A2(n_332),
.B1(n_313),
.B2(n_325),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_364),
.C(n_376),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_411),
.C(n_417),
.Y(n_424)
);

XNOR2x1_ASAP7_75t_SL g407 ( 
.A(n_377),
.B(n_335),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_407),
.B(n_419),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_345),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_360),
.A2(n_356),
.B1(n_377),
.B2(n_352),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_414),
.A2(n_375),
.B1(n_381),
.B2(n_371),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_359),
.A2(n_338),
.B1(n_341),
.B2(n_340),
.Y(n_416)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_416),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_373),
.B(n_341),
.C(n_340),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_365),
.A2(n_338),
.B1(n_348),
.B2(n_339),
.Y(n_418)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_385),
.B(n_339),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_422),
.A2(n_436),
.B1(n_444),
.B2(n_415),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_368),
.Y(n_428)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_366),
.Y(n_429)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_430),
.B(n_431),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_405),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_396),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_375),
.C(n_333),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_446),
.C(n_400),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_414),
.A2(n_384),
.B1(n_382),
.B2(n_386),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_333),
.Y(n_437)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_437),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_410),
.A2(n_326),
.B(n_342),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_439),
.B(n_389),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_410),
.A2(n_326),
.B(n_13),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_390),
.B(n_326),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_404),
.Y(n_458)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_392),
.B(n_1),
.Y(n_442)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_402),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_443)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_415),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_399),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_391),
.B(n_5),
.C(n_11),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_440),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_448),
.B(n_458),
.Y(n_479)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_453),
.A2(n_466),
.B1(n_468),
.B2(n_425),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_406),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_459),
.B(n_446),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_424),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_467),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_463),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_397),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_398),
.C(n_408),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_464),
.B(n_423),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_422),
.A2(n_415),
.B1(n_407),
.B2(n_398),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_411),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_469),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_447),
.A2(n_420),
.B(n_429),
.C(n_428),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_470),
.A2(n_480),
.B(n_483),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_435),
.C(n_425),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_477),
.C(n_448),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_427),
.Y(n_472)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_472),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_451),
.A2(n_436),
.B1(n_432),
.B2(n_442),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_473),
.A2(n_481),
.B1(n_457),
.B2(n_456),
.Y(n_498)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_453),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_423),
.C(n_438),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_484),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_450),
.B(n_413),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_465),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_437),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_450),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_487),
.B(n_458),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_493),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_473),
.A2(n_468),
.B1(n_466),
.B2(n_395),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_496),
.Y(n_507)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_485),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_490),
.B(n_482),
.Y(n_508)
);

AOI21x1_ASAP7_75t_SL g493 ( 
.A1(n_483),
.A2(n_409),
.B(n_439),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_462),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_476),
.A2(n_409),
.B(n_455),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_497),
.A2(n_501),
.B(n_470),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_500),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_467),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_419),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_475),
.A2(n_395),
.B1(n_456),
.B2(n_457),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_481),
.A2(n_413),
.B(n_464),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_475),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_502),
.B(n_508),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_503),
.B(n_504),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_486),
.A2(n_477),
.B1(n_443),
.B2(n_445),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_494),
.B(n_485),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_505),
.A2(n_506),
.B(n_509),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_482),
.C(n_479),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_399),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_512),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_513),
.B(n_499),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_5),
.C(n_17),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_514),
.A2(n_492),
.B(n_495),
.Y(n_517)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_517),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_497),
.B(n_489),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_518),
.A2(n_511),
.B(n_504),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_513),
.C(n_510),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_488),
.C(n_500),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_522),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_493),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_524),
.A2(n_526),
.B(n_14),
.Y(n_531)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_516),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_519),
.B1(n_515),
.B2(n_523),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_530),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_525),
.A2(n_523),
.B(n_510),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_531),
.A2(n_527),
.B(n_15),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_532),
.B(n_16),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_533),
.B(n_14),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_14),
.B1(n_15),
.B2(n_393),
.Y(n_536)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_536),
.Y(n_537)
);


endmodule