module fake_ariane_1432_n_2485 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2485);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2485;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2271;
wire n_2116;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_2075;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1865;
wire n_1710;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_39),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_43),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_417),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_508),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_479),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_194),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_324),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_444),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_312),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_112),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_122),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_474),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_341),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_127),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_90),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_316),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_174),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_495),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_9),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_247),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_116),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_46),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_183),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_307),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_290),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_258),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_178),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_199),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_155),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_111),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_461),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_176),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_438),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_288),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_320),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_228),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_416),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_509),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_229),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_132),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_108),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_317),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_294),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_498),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_139),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_128),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_415),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_328),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_230),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_51),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_366),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_477),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_66),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_216),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_291),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_0),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_344),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_302),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_56),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_132),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_401),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_75),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_504),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_323),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_197),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_28),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_484),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_378),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_11),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_281),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_515),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_88),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_166),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_71),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_17),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_81),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_150),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_376),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_493),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_109),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_246),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_17),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_131),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_28),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_204),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_77),
.Y(n_612)
);

BUFx2_ASAP7_75t_SL g613 ( 
.A(n_507),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_471),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_482),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_492),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_384),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_516),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_177),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_221),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_68),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_150),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_56),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_196),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_501),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_276),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_86),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_145),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_411),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_514),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_500),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_505),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_18),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_98),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_129),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_244),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_20),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_177),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_437),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_502),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_267),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_126),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_214),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_226),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_261),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_284),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_442),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_496),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_395),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_4),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_480),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_248),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_176),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_237),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_262),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_510),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_334),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_347),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_72),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_85),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_467),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_240),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_193),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_82),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_494),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_104),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_2),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_122),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_459),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_308),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_160),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_358),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_511),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_306),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_208),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_275),
.Y(n_678)
);

CKINVDCx14_ASAP7_75t_R g679 ( 
.A(n_40),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_121),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_456),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_185),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_435),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_491),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_419),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_145),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_22),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_483),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_490),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_430),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_298),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_260),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_133),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_280),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_15),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_227),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_421),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_191),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_175),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_367),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_473),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_167),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_321),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_59),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_481),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_455),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_488),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_325),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_30),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_319),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_29),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_136),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_497),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_374),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_454),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_25),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_71),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_101),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_441),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_209),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_406),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_287),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_422),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_499),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_485),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_32),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_362),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_114),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_396),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_402),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_111),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_436),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_243),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_475),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_427),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_106),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_7),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_338),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_30),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_80),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_57),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_239),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_174),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_135),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_155),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_365),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_329),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_478),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_556),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_556),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_745),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_745),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_527),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_535),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_535),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_534),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_567),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_595),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_543),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_547),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_553),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_573),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_558),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_571),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_585),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_585),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_611),
.Y(n_767)
);

INVxp33_ASAP7_75t_SL g768 ( 
.A(n_548),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_695),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_535),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_611),
.Y(n_771)
);

CKINVDCx16_ASAP7_75t_R g772 ( 
.A(n_679),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_580),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_564),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_535),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_574),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_588),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_522),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_679),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_592),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_599),
.Y(n_781)
);

INVxp33_ASAP7_75t_L g782 ( 
.A(n_554),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_523),
.Y(n_783)
);

INVxp33_ASAP7_75t_SL g784 ( 
.A(n_538),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_610),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_662),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_622),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_677),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_624),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_677),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_539),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_629),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_635),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_677),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_680),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_682),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_541),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_702),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_545),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_552),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_718),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_566),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_720),
.Y(n_803)
);

CKINVDCx14_ASAP7_75t_R g804 ( 
.A(n_526),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_572),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_576),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_726),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_728),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_537),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_582),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_744),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_586),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_554),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_591),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_598),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_623),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_623),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_637),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_637),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_689),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_630),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_579),
.Y(n_823)
);

BUFx2_ASAP7_75t_SL g824 ( 
.A(n_526),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_640),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_644),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_731),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_600),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_630),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_639),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_564),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_684),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_581),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_628),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_601),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_723),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_602),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_526),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_684),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_546),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_546),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_603),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_639),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_546),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_606),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_703),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_704),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_608),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_703),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_762),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_765),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_757),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_824),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_758),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_765),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_776),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_766),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_770),
.Y(n_858)
);

CKINVDCx16_ASAP7_75t_R g859 ( 
.A(n_772),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_794),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_809),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_766),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_753),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_838),
.B(n_722),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_756),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_786),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_759),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_767),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_760),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_778),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_767),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_761),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_763),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_764),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_783),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_791),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_771),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_797),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_840),
.B(n_605),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_773),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_771),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_777),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_799),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_780),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_800),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_829),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_802),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_809),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_781),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_785),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_829),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_805),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_787),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_830),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_769),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_774),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_806),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_779),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_830),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_774),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_789),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_792),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_793),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_810),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_812),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_849),
.B(n_529),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_795),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_831),
.Y(n_908)
);

INVxp33_ASAP7_75t_SL g909 ( 
.A(n_814),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_796),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_841),
.B(n_530),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_822),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_815),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_798),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_864),
.A2(n_768),
.B1(n_784),
.B2(n_828),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_SL g916 ( 
.A1(n_851),
.A2(n_704),
.B1(n_847),
.B2(n_843),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_861),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_861),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_870),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_888),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_911),
.B(n_528),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_888),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_858),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_863),
.B(n_846),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_865),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_860),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_867),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_869),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_866),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_872),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_873),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_896),
.B(n_844),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_R g933 ( 
.A(n_875),
.B(n_804),
.Y(n_933)
);

OA21x2_ASAP7_75t_L g934 ( 
.A1(n_906),
.A2(n_532),
.B(n_528),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_874),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_854),
.B(n_912),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_880),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_908),
.B(n_831),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_876),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_882),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_884),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_889),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_900),
.B(n_832),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_890),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_893),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_901),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_898),
.B(n_804),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_902),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_903),
.B(n_832),
.Y(n_949)
);

XNOR2x2_ASAP7_75t_R g950 ( 
.A(n_851),
.B(n_843),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_878),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_883),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_895),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_907),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_859),
.B(n_782),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_857),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_910),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_914),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_885),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_887),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_879),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_853),
.Y(n_962)
);

AND3x2_ASAP7_75t_L g963 ( 
.A(n_852),
.B(n_834),
.C(n_833),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_892),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_897),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_904),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_905),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_913),
.B(n_782),
.Y(n_968)
);

CKINVDCx16_ASAP7_75t_R g969 ( 
.A(n_862),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_850),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_856),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_909),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_899),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_877),
.Y(n_974)
);

AND2x6_ASAP7_75t_L g975 ( 
.A(n_894),
.B(n_532),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_855),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_855),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_891),
.Y(n_978)
);

INVxp67_ASAP7_75t_SL g979 ( 
.A(n_868),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_868),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_871),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_871),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_881),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_881),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_886),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_886),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_891),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_864),
.A2(n_768),
.B1(n_661),
.B2(n_670),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_870),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_896),
.B(n_821),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_908),
.B(n_839),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_863),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_863),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_908),
.B(n_839),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_908),
.B(n_846),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_863),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_861),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_861),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_863),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_896),
.B(n_835),
.Y(n_1000)
);

CKINVDCx11_ASAP7_75t_R g1001 ( 
.A(n_857),
.Y(n_1001)
);

CKINVDCx8_ASAP7_75t_R g1002 ( 
.A(n_859),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_863),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_895),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_923),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_968),
.Y(n_1006)
);

INVxp33_ASAP7_75t_SL g1007 ( 
.A(n_972),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_965),
.B(n_837),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_917),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_926),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_936),
.B(n_836),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_918),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_SL g1013 ( 
.A(n_1002),
.B(n_672),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_920),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_925),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_998),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_927),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_922),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_921),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_961),
.B(n_842),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_965),
.B(n_845),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_922),
.Y(n_1022)
);

INVxp33_ASAP7_75t_SL g1023 ( 
.A(n_919),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_955),
.B(n_848),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_997),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_997),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_918),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_918),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_965),
.B(n_989),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_918),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_930),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_927),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_953),
.B(n_749),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_927),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_927),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_954),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_935),
.B(n_593),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_931),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_954),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_954),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_937),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_953),
.B(n_750),
.Y(n_1042)
);

AND3x2_ASAP7_75t_L g1043 ( 
.A(n_970),
.B(n_847),
.C(n_803),
.Y(n_1043)
);

AO21x2_ASAP7_75t_L g1044 ( 
.A1(n_949),
.A2(n_536),
.B(n_531),
.Y(n_1044)
);

AO22x2_ASAP7_75t_L g1045 ( 
.A1(n_988),
.A2(n_698),
.B1(n_621),
.B2(n_801),
.Y(n_1045)
);

INVx5_ASAP7_75t_L g1046 ( 
.A(n_921),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_959),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_954),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_941),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1004),
.B(n_751),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_965),
.B(n_807),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_935),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_944),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_928),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_1000),
.B(n_672),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_940),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_956),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_921),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_942),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_945),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_948),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_957),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_924),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_988),
.B(n_915),
.C(n_1000),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_924),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_946),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_1004),
.B(n_710),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_947),
.B(n_752),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_934),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_934),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_929),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_958),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_939),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_964),
.B(n_540),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_992),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_SL g1076 ( 
.A(n_951),
.B(n_710),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_993),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_996),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_943),
.B(n_659),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_999),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1003),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_921),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_969),
.B(n_808),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_990),
.B(n_811),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_L g1085 ( 
.A(n_932),
.B(n_612),
.C(n_609),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_949),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_938),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_962),
.B(n_557),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_938),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_991),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_990),
.B(n_813),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_932),
.B(n_816),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_991),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_978),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_952),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_994),
.Y(n_1096)
);

AND3x2_ASAP7_75t_L g1097 ( 
.A(n_979),
.B(n_818),
.C(n_817),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_994),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_960),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_995),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_971),
.B(n_625),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_995),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_943),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_921),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_963),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_963),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_975),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_975),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_975),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_966),
.B(n_626),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_967),
.B(n_568),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_975),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_984),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_983),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_933),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_984),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_984),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_933),
.B(n_746),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_979),
.B(n_636),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_974),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_976),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_984),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_987),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_987),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_973),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_982),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_987),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_987),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_973),
.Y(n_1130)
);

NAND2xp33_ASAP7_75t_SL g1131 ( 
.A(n_973),
.B(n_645),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_985),
.B(n_577),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_973),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1001),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_977),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_985),
.B(n_584),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_986),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_980),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_981),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_950),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_916),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_SL g1142 ( 
.A(n_916),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_917),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1082),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1072),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1055),
.B(n_666),
.C(n_655),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1072),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_R g1148 ( 
.A(n_1099),
.B(n_652),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1047),
.Y(n_1149)
);

AND2x6_ASAP7_75t_L g1150 ( 
.A(n_1082),
.B(n_667),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1017),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1006),
.B(n_665),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1029),
.B(n_819),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1011),
.B(n_823),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1092),
.B(n_668),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1052),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1067),
.B(n_669),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1064),
.B(n_709),
.C(n_687),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1017),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_1029),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1077),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1017),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1006),
.B(n_673),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1116),
.B(n_686),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1047),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1052),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_1029),
.B(n_825),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1023),
.B(n_693),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1077),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1078),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1018),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1078),
.Y(n_1172)
);

XOR2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1076),
.B(n_826),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1015),
.Y(n_1174)
);

CKINVDCx16_ASAP7_75t_R g1175 ( 
.A(n_1073),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_1029),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1092),
.B(n_699),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1057),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1018),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_L g1180 ( 
.A(n_1082),
.B(n_711),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1022),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1017),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_R g1183 ( 
.A(n_1099),
.B(n_1116),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_1082),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1031),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1011),
.B(n_827),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1038),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1071),
.Y(n_1188)
);

OAI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1073),
.A2(n_716),
.B1(n_736),
.B2(n_712),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1083),
.B(n_717),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1019),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1103),
.B(n_737),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1084),
.B(n_739),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1051),
.B(n_754),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1022),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_1095),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1041),
.Y(n_1197)
);

CKINVDCx16_ASAP7_75t_R g1198 ( 
.A(n_1095),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1023),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1095),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1025),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1090),
.B(n_740),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1020),
.B(n_741),
.Y(n_1203)
);

NAND3x1_ASAP7_75t_L g1204 ( 
.A(n_1140),
.B(n_594),
.C(n_587),
.Y(n_1204)
);

INVx4_ASAP7_75t_L g1205 ( 
.A(n_1046),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1134),
.Y(n_1206)
);

AND2x4_ASAP7_75t_SL g1207 ( 
.A(n_1127),
.B(n_657),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1134),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1049),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1134),
.B(n_613),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1093),
.B(n_743),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1051),
.B(n_754),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1025),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1094),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1051),
.B(n_755),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1100),
.B(n_590),
.Y(n_1216)
);

AND2x6_ASAP7_75t_L g1217 ( 
.A(n_1104),
.B(n_667),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1026),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1053),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1026),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1066),
.Y(n_1221)
);

INVxp33_ASAP7_75t_SL g1222 ( 
.A(n_1111),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1087),
.B(n_732),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1114),
.B(n_755),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1009),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1020),
.B(n_657),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1007),
.B(n_657),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1009),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1024),
.B(n_524),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1101),
.A2(n_615),
.B1(n_616),
.B2(n_597),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1007),
.B(n_633),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1134),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1087),
.B(n_748),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_1046),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1014),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1014),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1126),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1046),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1075),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1024),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1076),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1089),
.B(n_638),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1080),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1084),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1046),
.B(n_525),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1126),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1046),
.B(n_533),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1081),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1037),
.B(n_542),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1042),
.B(n_775),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1089),
.B(n_643),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1016),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1096),
.B(n_1098),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1114),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1032),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1013),
.B(n_649),
.Y(n_1256)
);

AND3x4_ASAP7_75t_L g1257 ( 
.A(n_1135),
.B(n_788),
.C(n_775),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1005),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1010),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1054),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1033),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1042),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1112),
.B(n_664),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1114),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1112),
.B(n_675),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1016),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1019),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1043),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1032),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1008),
.A2(n_685),
.B1(n_692),
.B2(n_678),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1019),
.B(n_544),
.Y(n_1271)
);

AND2x6_ASAP7_75t_L g1272 ( 
.A(n_1104),
.B(n_688),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1085),
.B(n_1120),
.C(n_1121),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1050),
.B(n_788),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1054),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1130),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1058),
.B(n_549),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1058),
.Y(n_1278)
);

INVxp33_ASAP7_75t_L g1279 ( 
.A(n_1050),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1091),
.B(n_790),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1130),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1056),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1056),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1034),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1119),
.B(n_697),
.Y(n_1285)
);

OAI221xp5_ASAP7_75t_L g1286 ( 
.A1(n_1122),
.A2(n_708),
.B1(n_724),
.B2(n_714),
.C(n_701),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1059),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1096),
.B(n_729),
.Y(n_1288)
);

BUFx10_ASAP7_75t_L g1289 ( 
.A(n_1097),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1059),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1142),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1034),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1117),
.B(n_730),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1060),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

NOR3xp33_ASAP7_75t_L g1296 ( 
.A(n_1008),
.B(n_735),
.C(n_734),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1133),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1143),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1117),
.B(n_1118),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1098),
.B(n_738),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1060),
.Y(n_1301)
);

NOR2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1137),
.B(n_742),
.Y(n_1302)
);

BUFx10_ASAP7_75t_L g1303 ( 
.A(n_1138),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1061),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1061),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1118),
.B(n_747),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1062),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1062),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1123),
.B(n_790),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1035),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1115),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1131),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1035),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_1131),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1102),
.B(n_820),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1058),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1063),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1115),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1133),
.Y(n_1320)
);

INVx5_ASAP7_75t_L g1321 ( 
.A(n_1113),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_1063),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1086),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1142),
.A2(n_688),
.B1(n_550),
.B2(n_559),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1137),
.B(n_551),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1063),
.Y(n_1326)
);

BUFx4f_ASAP7_75t_L g1327 ( 
.A(n_1106),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1142),
.Y(n_1328)
);

NAND2xp33_ASAP7_75t_L g1329 ( 
.A(n_1021),
.B(n_560),
.Y(n_1329)
);

AND2x6_ASAP7_75t_L g1330 ( 
.A(n_1107),
.B(n_537),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1086),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1036),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1102),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1036),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1141),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1091),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1039),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1039),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1137),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1068),
.B(n_0),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1040),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1065),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1124),
.B(n_561),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1135),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1139),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1021),
.B(n_563),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1222),
.B(n_1106),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1262),
.B(n_1079),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1157),
.A2(n_1045),
.B1(n_1139),
.B2(n_1136),
.C(n_1132),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1183),
.B(n_1105),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1336),
.B(n_1261),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1151),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1244),
.B(n_1125),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1155),
.B(n_1125),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1174),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1185),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1145),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1187),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1175),
.B(n_1105),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1177),
.B(n_1128),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1196),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1256),
.A2(n_1045),
.B1(n_1074),
.B2(n_1132),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1285),
.B(n_1128),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1279),
.B(n_1129),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1197),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1250),
.B(n_1129),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1145),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1209),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1219),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1274),
.B(n_1074),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1221),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1160),
.B(n_1176),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1170),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1240),
.B(n_1141),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1323),
.B(n_1141),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1196),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1231),
.B(n_1136),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1331),
.B(n_1045),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1170),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1165),
.B(n_1065),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1160),
.B(n_1176),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1304),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1227),
.B(n_1088),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1280),
.B(n_1065),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1200),
.B(n_1113),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1253),
.B(n_1088),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1193),
.B(n_1044),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1333),
.B(n_1040),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1154),
.B(n_1186),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1239),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1340),
.B(n_1327),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1327),
.B(n_1344),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1206),
.Y(n_1393)
);

OAI22x1_ASAP7_75t_SL g1394 ( 
.A1(n_1199),
.A2(n_569),
.B1(n_570),
.B2(n_565),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1307),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1345),
.B(n_1048),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1335),
.B(n_1048),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1196),
.B(n_1107),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1168),
.A2(n_1108),
.B(n_1110),
.C(n_1109),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1315),
.B(n_1109),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1243),
.B(n_1248),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1241),
.B(n_1027),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1263),
.A2(n_1044),
.B1(n_1012),
.B2(n_1028),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1149),
.B(n_1188),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1208),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1214),
.B(n_1012),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1178),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1147),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1265),
.B(n_1044),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1161),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1169),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1313),
.B(n_1012),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1172),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1302),
.B(n_1027),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1312),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1192),
.B(n_1028),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1202),
.B(n_1030),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1211),
.B(n_1030),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1319),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1339),
.A2(n_1070),
.B1(n_1069),
.B2(n_578),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1153),
.B(n_1069),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1225),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1230),
.A2(n_1070),
.B(n_583),
.C(n_589),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_SL g1424 ( 
.A(n_1232),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1153),
.B(n_1),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1258),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1198),
.B(n_1303),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1194),
.B(n_1),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1194),
.B(n_2),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1303),
.B(n_575),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1273),
.A2(n_604),
.B(n_607),
.C(n_596),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1257),
.A2(n_555),
.B1(n_562),
.B2(n_537),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1200),
.B(n_1167),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1190),
.B(n_3),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1146),
.B(n_1203),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1228),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1259),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1212),
.B(n_3),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1229),
.B(n_614),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1167),
.B(n_537),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1212),
.B(n_4),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1235),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1260),
.Y(n_1443)
);

AND2x4_ASAP7_75t_SL g1444 ( 
.A(n_1210),
.B(n_555),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1226),
.B(n_617),
.Y(n_1445)
);

BUFx5_ASAP7_75t_L g1446 ( 
.A(n_1150),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1189),
.B(n_618),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1148),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1215),
.B(n_5),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1207),
.B(n_1215),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1236),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1237),
.B(n_619),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1246),
.B(n_1318),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1216),
.B(n_5),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1329),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1324),
.B(n_6),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1249),
.A2(n_1277),
.B(n_1271),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1254),
.A2(n_1264),
.B1(n_1158),
.B2(n_1191),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1210),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1318),
.B(n_620),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1291),
.B(n_8),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1328),
.B(n_9),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1322),
.B(n_1254),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1322),
.B(n_627),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1252),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1152),
.B(n_631),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1224),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1286),
.A2(n_634),
.B1(n_641),
.B2(n_632),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1223),
.B(n_10),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1264),
.B(n_642),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1289),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1266),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1295),
.Y(n_1473)
);

NOR2xp67_ASAP7_75t_L g1474 ( 
.A(n_1182),
.B(n_225),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1275),
.A2(n_562),
.B1(n_555),
.B2(n_646),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1233),
.B(n_10),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1242),
.B(n_11),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1156),
.A2(n_648),
.B(n_647),
.Y(n_1478)
);

NOR3xp33_ASAP7_75t_L g1479 ( 
.A(n_1346),
.B(n_651),
.C(n_650),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1296),
.B(n_653),
.Y(n_1480)
);

NOR3xp33_ASAP7_75t_L g1481 ( 
.A(n_1164),
.B(n_656),
.C(n_654),
.Y(n_1481)
);

NAND2x1_ASAP7_75t_L g1482 ( 
.A(n_1205),
.B(n_555),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1163),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1268),
.B(n_12),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1282),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1298),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1251),
.B(n_12),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1283),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1288),
.B(n_13),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1300),
.B(n_13),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1287),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1326),
.B(n_658),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1290),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1294),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1301),
.A2(n_562),
.B1(n_663),
.B2(n_660),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1326),
.B(n_671),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1305),
.A2(n_562),
.B1(n_676),
.B2(n_674),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1166),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1151),
.B(n_681),
.Y(n_1499)
);

NOR2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1342),
.B(n_683),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1224),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1308),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1276),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1171),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1299),
.B(n_14),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1151),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1316),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1159),
.B(n_690),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1179),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1309),
.B(n_14),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1181),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1281),
.B(n_15),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1270),
.A2(n_694),
.B(n_696),
.C(n_691),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1297),
.A2(n_705),
.B1(n_706),
.B2(n_700),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1342),
.B(n_707),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1320),
.B(n_713),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1325),
.B(n_719),
.C(n_715),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1343),
.B(n_16),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1293),
.A2(n_725),
.B1(n_727),
.B2(n_721),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1306),
.B(n_16),
.Y(n_1520)
);

NAND2xp33_ASAP7_75t_L g1521 ( 
.A(n_1159),
.B(n_733),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1159),
.Y(n_1522)
);

O2A1O1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1180),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1523)
);

AND2x6_ASAP7_75t_SL g1524 ( 
.A(n_1310),
.B(n_19),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1191),
.A2(n_809),
.B(n_232),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1195),
.B(n_21),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1201),
.B(n_21),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1213),
.B(n_22),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1218),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1220),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_SL g1531 ( 
.A(n_1289),
.B(n_809),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1310),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1255),
.B(n_23),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1162),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1255),
.B(n_23),
.Y(n_1535)
);

NOR2x1p5_ASAP7_75t_L g1536 ( 
.A(n_1182),
.B(n_24),
.Y(n_1536)
);

AOI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1245),
.A2(n_233),
.B(n_231),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1255),
.B(n_24),
.Y(n_1538)
);

BUFx8_ASAP7_75t_L g1539 ( 
.A(n_1150),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1334),
.B(n_25),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1144),
.B(n_26),
.Y(n_1541)
);

OAI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1173),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.C(n_31),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1267),
.A2(n_235),
.B(n_234),
.Y(n_1543)
);

O2A1O1Ixp5_ASAP7_75t_L g1544 ( 
.A1(n_1247),
.A2(n_32),
.B(n_27),
.C(n_31),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1341),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1311),
.Y(n_1546)
);

NOR3xp33_ASAP7_75t_L g1547 ( 
.A(n_1314),
.B(n_33),
.C(n_34),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1184),
.B(n_33),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1269),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1332),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1337),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1338),
.B(n_34),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1162),
.B(n_35),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1269),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1162),
.B(n_35),
.Y(n_1555)
);

AND2x6_ASAP7_75t_L g1556 ( 
.A(n_1267),
.B(n_236),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1269),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1411),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1377),
.B(n_1389),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_R g1560 ( 
.A(n_1448),
.B(n_1150),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1393),
.Y(n_1561)
);

INVx5_ASAP7_75t_L g1562 ( 
.A(n_1556),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1355),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1356),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1383),
.B(n_1284),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1348),
.B(n_1284),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1407),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1391),
.B(n_1284),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1357),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1397),
.B(n_1374),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1367),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1450),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1461),
.B(n_1292),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1381),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1381),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1358),
.Y(n_1576)
);

INVx5_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1447),
.A2(n_1204),
.B1(n_1150),
.B2(n_1278),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1468),
.A2(n_1317),
.B1(n_1278),
.B2(n_1217),
.Y(n_1579)
);

INVx5_ASAP7_75t_L g1580 ( 
.A(n_1556),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1501),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1541),
.B(n_1292),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1373),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1434),
.B(n_1292),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1467),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1365),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1349),
.B(n_1217),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1351),
.B(n_1217),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1433),
.B(n_1321),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1440),
.B(n_1205),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1405),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1379),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1433),
.B(n_1321),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1503),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1471),
.B(n_1321),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1468),
.A2(n_1317),
.B1(n_1272),
.B2(n_1217),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1401),
.B(n_1272),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1387),
.B(n_1272),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1362),
.A2(n_1272),
.B1(n_1330),
.B2(n_1238),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1368),
.B(n_1330),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1601)
);

BUFx2_ASAP7_75t_SL g1602 ( 
.A(n_1424),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1361),
.B(n_1234),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1518),
.A2(n_1238),
.B(n_1234),
.C(n_1330),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1459),
.Y(n_1605)
);

INVx5_ASAP7_75t_L g1606 ( 
.A(n_1556),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1390),
.B(n_1330),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1424),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1376),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1382),
.Y(n_1610)
);

INVx4_ASAP7_75t_L g1611 ( 
.A(n_1352),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1375),
.B(n_36),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1541),
.B(n_36),
.Y(n_1613)
);

BUFx4f_ASAP7_75t_L g1614 ( 
.A(n_1444),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1352),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1426),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1395),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1353),
.B(n_1404),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1440),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1507),
.B(n_37),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1392),
.B(n_37),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1402),
.B(n_38),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1359),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1362),
.B(n_38),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1370),
.B(n_39),
.Y(n_1625)
);

BUFx8_ASAP7_75t_L g1626 ( 
.A(n_1484),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1500),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1350),
.B(n_521),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1428),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1422),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1427),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1437),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1456),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1364),
.B(n_41),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1436),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1352),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1522),
.Y(n_1637)
);

AND2x2_ASAP7_75t_SL g1638 ( 
.A(n_1432),
.B(n_42),
.Y(n_1638)
);

OR2x2_ASAP7_75t_SL g1639 ( 
.A(n_1462),
.B(n_43),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1386),
.B(n_44),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1363),
.B(n_44),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1408),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1347),
.B(n_45),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1440),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1516),
.B(n_1454),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1522),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1435),
.B(n_45),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1536),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1442),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1534),
.B(n_238),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1412),
.B(n_46),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1398),
.B(n_1549),
.Y(n_1652)
);

O2A1O1Ixp5_ASAP7_75t_L g1653 ( 
.A1(n_1520),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1653)
);

AND2x6_ASAP7_75t_SL g1654 ( 
.A(n_1439),
.B(n_47),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1410),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1413),
.B(n_48),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1425),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1415),
.Y(n_1658)
);

A2O1A1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1455),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1451),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1519),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1483),
.B(n_52),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1419),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1545),
.B(n_53),
.Y(n_1664)
);

OR2x6_ASAP7_75t_L g1665 ( 
.A(n_1372),
.B(n_54),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1443),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1398),
.B(n_520),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1522),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_L g1669 ( 
.A(n_1517),
.B(n_54),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1546),
.B(n_55),
.Y(n_1670)
);

INVx5_ASAP7_75t_L g1671 ( 
.A(n_1534),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1539),
.B(n_1531),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1384),
.B(n_55),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1539),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1485),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1414),
.B(n_57),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1458),
.B(n_1519),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1488),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_R g1679 ( 
.A(n_1521),
.B(n_241),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1469),
.B(n_58),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1491),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1409),
.B(n_58),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1429),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1406),
.B(n_59),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1685)
);

INVx5_ASAP7_75t_L g1686 ( 
.A(n_1506),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1506),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1493),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1378),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_L g1690 ( 
.A(n_1554),
.B(n_242),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1465),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1494),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1438),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1502),
.Y(n_1694)
);

AND2x6_ASAP7_75t_SL g1695 ( 
.A(n_1445),
.B(n_63),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1354),
.B(n_1360),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1529),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1487),
.B(n_63),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1557),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1489),
.B(n_1490),
.Y(n_1700)
);

O2A1O1Ixp5_ASAP7_75t_L g1701 ( 
.A1(n_1457),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1498),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1472),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1441),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1533),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1400),
.B(n_64),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1530),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1473),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1449),
.B(n_65),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1504),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1535),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1486),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1512),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1394),
.Y(n_1714)
);

AOI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1399),
.A2(n_67),
.B(n_68),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1509),
.Y(n_1716)
);

OAI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1542),
.A2(n_1547),
.B1(n_1523),
.B2(n_1466),
.C(n_1423),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1511),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1532),
.B(n_519),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1430),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1550),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1421),
.B(n_67),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1538),
.A2(n_72),
.B1(n_69),
.B2(n_70),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1480),
.A2(n_1496),
.B1(n_1515),
.B2(n_1492),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1524),
.B(n_69),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1524),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1478),
.A2(n_74),
.B1(n_70),
.B2(n_73),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1551),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1416),
.B(n_73),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1526),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1396),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1527),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1540),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1528),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1417),
.B(n_74),
.Y(n_1735)
);

BUFx8_ASAP7_75t_L g1736 ( 
.A(n_1446),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1552),
.Y(n_1737)
);

BUFx4f_ASAP7_75t_L g1738 ( 
.A(n_1452),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1388),
.Y(n_1739)
);

AO22x1_ASAP7_75t_L g1740 ( 
.A1(n_1481),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1366),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1418),
.B(n_76),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1548),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_SL g1744 ( 
.A(n_1479),
.B(n_78),
.C(n_79),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1380),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1505),
.B(n_78),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1510),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1446),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1544),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_SL g1750 ( 
.A(n_1446),
.B(n_245),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1403),
.B(n_79),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1537),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1553),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1453),
.Y(n_1754)
);

INVx11_ASAP7_75t_L g1755 ( 
.A(n_1626),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1724),
.A2(n_1513),
.B(n_1431),
.C(n_1403),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1559),
.A2(n_1555),
.B1(n_1508),
.B2(n_1499),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1638),
.A2(n_1514),
.B1(n_1385),
.B2(n_1464),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1562),
.B(n_1577),
.Y(n_1759)
);

AOI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1677),
.A2(n_1420),
.B(n_1482),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1561),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1645),
.B(n_1470),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1594),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1574),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1558),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1591),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1562),
.A2(n_1463),
.B(n_1543),
.Y(n_1767)
);

AOI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1685),
.A2(n_1525),
.B(n_1474),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1567),
.B(n_1460),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1741),
.B(n_1495),
.Y(n_1770)
);

CKINVDCx10_ASAP7_75t_R g1771 ( 
.A(n_1665),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1608),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1566),
.B(n_1497),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1647),
.A2(n_1475),
.B1(n_1474),
.B2(n_1446),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1747),
.B(n_1446),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1565),
.B(n_80),
.Y(n_1776)
);

AOI21x1_ASAP7_75t_L g1777 ( 
.A1(n_1751),
.A2(n_250),
.B(n_249),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1601),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1562),
.A2(n_81),
.B(n_82),
.Y(n_1779)
);

BUFx4f_ASAP7_75t_L g1780 ( 
.A(n_1574),
.Y(n_1780)
);

NAND2x1p5_ASAP7_75t_L g1781 ( 
.A(n_1614),
.B(n_251),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1577),
.A2(n_83),
.B(n_84),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1669),
.B(n_83),
.C(n_84),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1563),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1705),
.B(n_85),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1573),
.B(n_86),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1585),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1577),
.A2(n_87),
.B(n_88),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1580),
.A2(n_87),
.B(n_89),
.Y(n_1789)
);

BUFx8_ASAP7_75t_L g1790 ( 
.A(n_1726),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_L g1791 ( 
.A(n_1711),
.B(n_89),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1695),
.B(n_90),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1580),
.B(n_91),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1717),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1657),
.B(n_92),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1580),
.B(n_1606),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1654),
.B(n_93),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1624),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1574),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1648),
.B(n_1665),
.Y(n_1800)
);

AO21x1_ASAP7_75t_L g1801 ( 
.A1(n_1682),
.A2(n_94),
.B(n_95),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1606),
.A2(n_96),
.B(n_97),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1581),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1606),
.A2(n_97),
.B(n_98),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1746),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1805)
);

NOR2x1_ASAP7_75t_L g1806 ( 
.A(n_1602),
.B(n_99),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1610),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1572),
.B(n_1584),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1604),
.A2(n_100),
.B(n_102),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1564),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1700),
.A2(n_102),
.B(n_103),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1693),
.B(n_103),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1615),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1696),
.A2(n_1750),
.B(n_1582),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1704),
.B(n_1733),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1578),
.B(n_104),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1640),
.A2(n_105),
.B(n_106),
.Y(n_1817)
);

AO21x1_ASAP7_75t_L g1818 ( 
.A1(n_1622),
.A2(n_105),
.B(n_107),
.Y(n_1818)
);

AOI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1752),
.A2(n_253),
.B(n_252),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1738),
.B(n_107),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1729),
.A2(n_108),
.B(n_109),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1605),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1735),
.A2(n_1579),
.B(n_1641),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1628),
.B(n_110),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1618),
.B(n_110),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1617),
.Y(n_1826)
);

AO21x1_ASAP7_75t_L g1827 ( 
.A1(n_1698),
.A2(n_112),
.B(n_113),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_1713),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1570),
.B(n_113),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1576),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1615),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1602),
.B(n_114),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1628),
.B(n_115),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1749),
.A2(n_115),
.B(n_116),
.Y(n_1834)
);

AND2x6_ASAP7_75t_L g1835 ( 
.A(n_1748),
.B(n_254),
.Y(n_1835)
);

NAND2x1p5_ASAP7_75t_L g1836 ( 
.A(n_1671),
.B(n_255),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1720),
.B(n_117),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1597),
.A2(n_117),
.B(n_118),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1659),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1730),
.A2(n_119),
.B(n_120),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1725),
.B(n_1662),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1679),
.B(n_121),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1590),
.A2(n_123),
.B(n_124),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1586),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1709),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1629),
.B(n_125),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1590),
.A2(n_126),
.B(n_127),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1616),
.B(n_1632),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_1581),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1743),
.B(n_128),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1714),
.B(n_129),
.Y(n_1851)
);

NOR4xp25_ASAP7_75t_L g1852 ( 
.A(n_1680),
.B(n_133),
.C(n_130),
.D(n_131),
.Y(n_1852)
);

INVx3_ASAP7_75t_L g1853 ( 
.A(n_1615),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1581),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1642),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1631),
.Y(n_1856)
);

OAI21xp33_ASAP7_75t_L g1857 ( 
.A1(n_1723),
.A2(n_130),
.B(n_134),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1706),
.A2(n_1613),
.B1(n_1744),
.B2(n_1684),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1630),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_SL g1860 ( 
.A1(n_1621),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1655),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1596),
.A2(n_137),
.B(n_138),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_SL g1863 ( 
.A(n_1672),
.B(n_256),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1587),
.A2(n_137),
.B(n_138),
.Y(n_1864)
);

O2A1O1Ixp5_ASAP7_75t_L g1865 ( 
.A1(n_1715),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1635),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1683),
.B(n_140),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1658),
.B(n_141),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1637),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1719),
.A2(n_1588),
.B(n_1732),
.Y(n_1870)
);

NOR2x1_ASAP7_75t_L g1871 ( 
.A(n_1706),
.B(n_142),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1663),
.Y(n_1872)
);

AOI21xp33_ASAP7_75t_L g1873 ( 
.A1(n_1734),
.A2(n_142),
.B(n_143),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1666),
.B(n_143),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1728),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1675),
.B(n_144),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1719),
.A2(n_144),
.B(n_146),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1678),
.B(n_146),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1681),
.B(n_147),
.Y(n_1879)
);

A2O1A1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1612),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1737),
.A2(n_1742),
.B(n_1722),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1639),
.B(n_148),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1727),
.A2(n_152),
.B1(n_149),
.B2(n_151),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1575),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1627),
.B(n_1643),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1661),
.A2(n_1753),
.B1(n_1633),
.B2(n_1625),
.Y(n_1886)
);

O2A1O1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1651),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1688),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1701),
.A2(n_153),
.B(n_154),
.Y(n_1889)
);

NAND2x1_ASAP7_75t_L g1890 ( 
.A(n_1611),
.B(n_257),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1673),
.A2(n_154),
.B(n_156),
.Y(n_1891)
);

INVx4_ASAP7_75t_L g1892 ( 
.A(n_1671),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1620),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1692),
.B(n_157),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1686),
.B(n_158),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1575),
.B(n_159),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1649),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1694),
.B(n_159),
.Y(n_1898)
);

CKINVDCx10_ASAP7_75t_R g1899 ( 
.A(n_1626),
.Y(n_1899)
);

AOI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1598),
.A2(n_263),
.B(n_259),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1686),
.B(n_160),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1691),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1600),
.A2(n_161),
.B(n_162),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1660),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1703),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1674),
.B(n_163),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1653),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1731),
.B(n_164),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1589),
.B(n_165),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1607),
.A2(n_167),
.B(n_168),
.Y(n_1910)
);

A2O1A1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1664),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1686),
.B(n_1575),
.Y(n_1912)
);

AOI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1568),
.A2(n_265),
.B(n_264),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1599),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1697),
.B(n_171),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1707),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1739),
.B(n_172),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1589),
.B(n_172),
.Y(n_1918)
);

OAI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1634),
.A2(n_173),
.B(n_175),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1593),
.B(n_173),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_SL g1921 ( 
.A(n_1593),
.B(n_266),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1780),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1760),
.A2(n_1650),
.B(n_1745),
.Y(n_1923)
);

INVx4_ASAP7_75t_L g1924 ( 
.A(n_1813),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1783),
.A2(n_1676),
.B(n_1689),
.Y(n_1925)
);

OAI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1768),
.A2(n_1819),
.B(n_1767),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1765),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1807),
.Y(n_1928)
);

OAI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1756),
.A2(n_1656),
.B(n_1670),
.Y(n_1929)
);

AOI21x1_ASAP7_75t_L g1930 ( 
.A1(n_1823),
.A2(n_1740),
.B(n_1690),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1778),
.B(n_1569),
.Y(n_1931)
);

OAI21x1_ASAP7_75t_L g1932 ( 
.A1(n_1900),
.A2(n_1777),
.B(n_1774),
.Y(n_1932)
);

OAI21x1_ASAP7_75t_L g1933 ( 
.A1(n_1809),
.A2(n_1583),
.B(n_1571),
.Y(n_1933)
);

AO31x2_ASAP7_75t_L g1934 ( 
.A1(n_1775),
.A2(n_1592),
.A3(n_1718),
.B(n_1716),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1815),
.B(n_1699),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1857),
.A2(n_1839),
.B(n_1794),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1814),
.A2(n_1667),
.B(n_1754),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1787),
.B(n_1623),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1870),
.A2(n_1667),
.B(n_1603),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1828),
.B(n_1619),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1759),
.A2(n_1603),
.B(n_1637),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1808),
.B(n_1644),
.Y(n_1942)
);

AOI21x1_ASAP7_75t_L g1943 ( 
.A1(n_1796),
.A2(n_1652),
.B(n_1609),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1871),
.A2(n_1652),
.B1(n_1687),
.B2(n_1736),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1862),
.A2(n_1646),
.B(n_1637),
.Y(n_1945)
);

AO21x2_ASAP7_75t_L g1946 ( 
.A1(n_1881),
.A2(n_1560),
.B(n_1708),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1786),
.B(n_1763),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1913),
.A2(n_1595),
.B(n_1636),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1824),
.A2(n_1833),
.B(n_1877),
.Y(n_1949)
);

A2O1A1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1858),
.A2(n_1840),
.B(n_1842),
.C(n_1919),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1826),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1822),
.B(n_1646),
.Y(n_1952)
);

AND2x2_ASAP7_75t_SL g1953 ( 
.A(n_1921),
.B(n_1611),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1761),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1865),
.A2(n_1671),
.B(n_1702),
.Y(n_1955)
);

OAI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1907),
.A2(n_1710),
.B(n_1712),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1841),
.B(n_1646),
.Y(n_1957)
);

OAI21x1_ASAP7_75t_L g1958 ( 
.A1(n_1903),
.A2(n_1910),
.B(n_1838),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1889),
.A2(n_1668),
.B(n_1736),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1854),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1909),
.B(n_1668),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1890),
.A2(n_1721),
.B(n_1668),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1820),
.B(n_178),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1836),
.A2(n_269),
.B(n_268),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1816),
.A2(n_179),
.B(n_180),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1886),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1912),
.A2(n_1793),
.B(n_1757),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1766),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1863),
.A2(n_181),
.B(n_182),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1772),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1784),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1779),
.A2(n_1788),
.B(n_1782),
.Y(n_1972)
);

OAI21x1_ASAP7_75t_L g1973 ( 
.A1(n_1864),
.A2(n_271),
.B(n_270),
.Y(n_1973)
);

AOI21xp33_ASAP7_75t_L g1974 ( 
.A1(n_1887),
.A2(n_182),
.B(n_183),
.Y(n_1974)
);

OAI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1834),
.A2(n_273),
.B(n_272),
.Y(n_1975)
);

INVxp67_ASAP7_75t_SL g1976 ( 
.A(n_1848),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1810),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1789),
.A2(n_184),
.B(n_185),
.Y(n_1978)
);

OAI21x1_ASAP7_75t_SL g1979 ( 
.A1(n_1801),
.A2(n_184),
.B(n_186),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1830),
.B(n_186),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1844),
.B(n_187),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1817),
.A2(n_187),
.B(n_188),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1855),
.B(n_188),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1802),
.A2(n_189),
.B(n_190),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1861),
.B(n_1872),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1780),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1804),
.A2(n_189),
.B(n_190),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1758),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1882),
.A2(n_195),
.B(n_192),
.C(n_194),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1762),
.A2(n_195),
.B(n_196),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1813),
.A2(n_277),
.B(n_274),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1892),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1920),
.B(n_197),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1883),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1891),
.A2(n_198),
.B(n_200),
.Y(n_1995)
);

INVx5_ASAP7_75t_L g1996 ( 
.A(n_1835),
.Y(n_1996)
);

AOI21xp33_ASAP7_75t_L g1997 ( 
.A1(n_1770),
.A2(n_201),
.B(n_202),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1792),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1888),
.B(n_1916),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1781),
.B(n_278),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1915),
.B(n_203),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1859),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1764),
.B(n_1799),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1894),
.B(n_204),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1764),
.B(n_279),
.Y(n_2005)
);

OA21x2_ASAP7_75t_L g2006 ( 
.A1(n_1773),
.A2(n_205),
.B(n_206),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1866),
.Y(n_2007)
);

AOI21xp33_ASAP7_75t_L g2008 ( 
.A1(n_1902),
.A2(n_205),
.B(n_206),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1897),
.Y(n_2009)
);

NAND2x1_ASAP7_75t_L g2010 ( 
.A(n_1892),
.B(n_207),
.Y(n_2010)
);

AO21x1_ASAP7_75t_L g2011 ( 
.A1(n_1821),
.A2(n_207),
.B(n_208),
.Y(n_2011)
);

AOI21x1_ASAP7_75t_L g2012 ( 
.A1(n_1776),
.A2(n_209),
.B(n_210),
.Y(n_2012)
);

OAI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1880),
.A2(n_210),
.B(n_211),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1825),
.B(n_211),
.Y(n_2014)
);

OAI21x1_ASAP7_75t_L g2015 ( 
.A1(n_1831),
.A2(n_283),
.B(n_282),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1856),
.B(n_212),
.Y(n_2016)
);

OAI22x1_ASAP7_75t_L g2017 ( 
.A1(n_1797),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1771),
.B(n_213),
.Y(n_2018)
);

OAI21x1_ASAP7_75t_L g2019 ( 
.A1(n_1831),
.A2(n_286),
.B(n_285),
.Y(n_2019)
);

OAI22x1_ASAP7_75t_L g2020 ( 
.A1(n_1837),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1896),
.B(n_215),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1829),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1860),
.A2(n_217),
.B(n_218),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1908),
.B(n_218),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1853),
.A2(n_292),
.B(n_289),
.Y(n_2025)
);

BUFx4_ASAP7_75t_SL g2026 ( 
.A(n_1970),
.Y(n_2026)
);

BUFx3_ASAP7_75t_L g2027 ( 
.A(n_1960),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1999),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1957),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1976),
.Y(n_2030)
);

BUFx2_ASAP7_75t_R g2031 ( 
.A(n_1952),
.Y(n_2031)
);

AOI22xp33_ASAP7_75t_L g2032 ( 
.A1(n_1936),
.A2(n_1827),
.B1(n_1818),
.B2(n_1805),
.Y(n_2032)
);

CKINVDCx6p67_ASAP7_75t_R g2033 ( 
.A(n_1996),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1934),
.Y(n_2034)
);

BUFx12f_ASAP7_75t_L g2035 ( 
.A(n_2001),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1947),
.B(n_1885),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1934),
.Y(n_2037)
);

INVx3_ASAP7_75t_L g2038 ( 
.A(n_1985),
.Y(n_2038)
);

BUFx12f_ASAP7_75t_L g2039 ( 
.A(n_1922),
.Y(n_2039)
);

INVx5_ASAP7_75t_L g2040 ( 
.A(n_1996),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1942),
.B(n_1906),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_1985),
.B(n_1846),
.Y(n_2042)
);

INVx4_ASAP7_75t_L g2043 ( 
.A(n_1996),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1992),
.Y(n_2044)
);

BUFx2_ASAP7_75t_L g2045 ( 
.A(n_1942),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_1992),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1935),
.B(n_1812),
.Y(n_2047)
);

BUFx12f_ASAP7_75t_L g2048 ( 
.A(n_1922),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1971),
.Y(n_2049)
);

BUFx2_ASAP7_75t_SL g2050 ( 
.A(n_1968),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1961),
.B(n_1940),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_1953),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1977),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1954),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1950),
.A2(n_1988),
.B1(n_1966),
.B2(n_2013),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1934),
.Y(n_2056)
);

INVx6_ASAP7_75t_SL g2057 ( 
.A(n_2005),
.Y(n_2057)
);

INVx3_ASAP7_75t_L g2058 ( 
.A(n_1924),
.Y(n_2058)
);

INVx2_ASAP7_75t_SL g2059 ( 
.A(n_2022),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1922),
.Y(n_2060)
);

BUFx12f_ASAP7_75t_L g2061 ( 
.A(n_1986),
.Y(n_2061)
);

BUFx2_ASAP7_75t_SL g2062 ( 
.A(n_1986),
.Y(n_2062)
);

INVx6_ASAP7_75t_SL g2063 ( 
.A(n_2005),
.Y(n_2063)
);

BUFx3_ASAP7_75t_L g2064 ( 
.A(n_1938),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2002),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2002),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1931),
.Y(n_2067)
);

NAND2x1p5_ASAP7_75t_L g2068 ( 
.A(n_1939),
.B(n_1853),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1980),
.B(n_1981),
.Y(n_2069)
);

BUFx2_ASAP7_75t_R g2070 ( 
.A(n_2003),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1986),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1927),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1983),
.B(n_1850),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1924),
.Y(n_2074)
);

INVxp67_ASAP7_75t_SL g2075 ( 
.A(n_1932),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1943),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1937),
.B(n_1791),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2007),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1929),
.B(n_1868),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2004),
.B(n_1874),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_2009),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1928),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1993),
.Y(n_2083)
);

BUFx3_ASAP7_75t_L g2084 ( 
.A(n_1962),
.Y(n_2084)
);

BUFx3_ASAP7_75t_L g2085 ( 
.A(n_1944),
.Y(n_2085)
);

AO21x2_ASAP7_75t_L g2086 ( 
.A1(n_2056),
.A2(n_1926),
.B(n_1979),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_SL g2087 ( 
.A1(n_2079),
.A2(n_1967),
.B(n_2012),
.Y(n_2087)
);

AOI21x1_ASAP7_75t_L g2088 ( 
.A1(n_2077),
.A2(n_1930),
.B(n_2006),
.Y(n_2088)
);

INVx3_ASAP7_75t_L g2089 ( 
.A(n_2074),
.Y(n_2089)
);

AO21x2_ASAP7_75t_L g2090 ( 
.A1(n_2075),
.A2(n_1946),
.B(n_1982),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_SL g2091 ( 
.A(n_2070),
.B(n_1963),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_2038),
.B(n_2021),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2053),
.Y(n_2093)
);

OAI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2055),
.A2(n_1969),
.B(n_1990),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_2068),
.A2(n_1923),
.B(n_1958),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2053),
.Y(n_2096)
);

NAND3xp33_ASAP7_75t_L g2097 ( 
.A(n_2032),
.B(n_1998),
.C(n_1989),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_2068),
.A2(n_1972),
.B(n_1959),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2030),
.B(n_2006),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2049),
.Y(n_2100)
);

OAI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2077),
.A2(n_1995),
.B(n_1949),
.Y(n_2101)
);

BUFx2_ASAP7_75t_L g2102 ( 
.A(n_2038),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_2074),
.Y(n_2103)
);

OAI21x1_ASAP7_75t_L g2104 ( 
.A1(n_2034),
.A2(n_1933),
.B(n_1948),
.Y(n_2104)
);

INVx6_ASAP7_75t_L g2105 ( 
.A(n_2052),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_2049),
.Y(n_2106)
);

AOI21x1_ASAP7_75t_L g2107 ( 
.A1(n_2073),
.A2(n_2014),
.B(n_2024),
.Y(n_2107)
);

OAI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_2052),
.A2(n_2000),
.B1(n_2017),
.B2(n_2020),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_2034),
.A2(n_1945),
.B(n_1955),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2065),
.Y(n_2110)
);

OA21x2_ASAP7_75t_L g2111 ( 
.A1(n_2037),
.A2(n_1997),
.B(n_1956),
.Y(n_2111)
);

AO21x2_ASAP7_75t_L g2112 ( 
.A1(n_2037),
.A2(n_1917),
.B(n_1878),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2066),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2078),
.Y(n_2114)
);

OAI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_2032),
.A2(n_1994),
.B(n_1811),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2028),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2045),
.B(n_1896),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2059),
.B(n_2016),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2083),
.A2(n_1914),
.B1(n_1798),
.B2(n_2085),
.Y(n_2119)
);

OR2x6_ASAP7_75t_L g2120 ( 
.A(n_2043),
.B(n_1941),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_2026),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_2040),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_SL g2123 ( 
.A1(n_2091),
.A2(n_2052),
.B1(n_2085),
.B2(n_2035),
.Y(n_2123)
);

BUFx4f_ASAP7_75t_SL g2124 ( 
.A(n_2121),
.Y(n_2124)
);

INVxp67_ASAP7_75t_SL g2125 ( 
.A(n_2106),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2093),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_SL g2127 ( 
.A1(n_2097),
.A2(n_2111),
.B1(n_2115),
.B2(n_2094),
.Y(n_2127)
);

BUFx6f_ASAP7_75t_L g2128 ( 
.A(n_2122),
.Y(n_2128)
);

OA21x2_ASAP7_75t_L g2129 ( 
.A1(n_2109),
.A2(n_2067),
.B(n_2047),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2096),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2110),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2112),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2112),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2113),
.Y(n_2134)
);

AOI21x1_ASAP7_75t_L g2135 ( 
.A1(n_2088),
.A2(n_2107),
.B(n_2087),
.Y(n_2135)
);

BUFx12f_ASAP7_75t_L g2136 ( 
.A(n_2118),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_2106),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2099),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_2100),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_2089),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2108),
.A2(n_2011),
.B1(n_2035),
.B2(n_2076),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2102),
.B(n_2064),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2114),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_2089),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2138),
.B(n_2059),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2132),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_2137),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2142),
.B(n_2092),
.Y(n_2148)
);

CKINVDCx20_ASAP7_75t_R g2149 ( 
.A(n_2124),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2135),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2131),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2142),
.B(n_2092),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_2128),
.Y(n_2153)
);

AO21x2_ASAP7_75t_L g2154 ( 
.A1(n_2150),
.A2(n_2135),
.B(n_2101),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2147),
.B(n_2127),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2151),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2147),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_SL g2158 ( 
.A(n_2149),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2145),
.A2(n_2141),
.B1(n_2108),
.B2(n_2123),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2157),
.B(n_2148),
.Y(n_2160)
);

A2O1A1Ixp33_ASAP7_75t_L g2161 ( 
.A1(n_2155),
.A2(n_1851),
.B(n_2018),
.C(n_2119),
.Y(n_2161)
);

AND2x4_ASAP7_75t_SL g2162 ( 
.A(n_2156),
.B(n_2149),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_2159),
.B(n_2143),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2154),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2154),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_2158),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_2157),
.B(n_2152),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2156),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2166),
.B(n_2153),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2162),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2168),
.B(n_2143),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2162),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2160),
.B(n_2153),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2167),
.Y(n_2174)
);

NOR2x1_ASAP7_75t_SL g2175 ( 
.A(n_2163),
.B(n_2050),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2165),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2161),
.B(n_2131),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2167),
.B(n_2140),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_2161),
.B(n_1899),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2170),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2172),
.B(n_2144),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2169),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2176),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_2177),
.A2(n_2164),
.B(n_1832),
.Y(n_2184)
);

INVx1_ASAP7_75t_SL g2185 ( 
.A(n_2179),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2171),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2173),
.Y(n_2187)
);

OAI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_2177),
.A2(n_1806),
.B(n_1845),
.Y(n_2188)
);

NOR3xp33_ASAP7_75t_L g2189 ( 
.A(n_2185),
.B(n_2174),
.C(n_2171),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2180),
.B(n_2178),
.Y(n_2190)
);

NOR3xp33_ASAP7_75t_L g2191 ( 
.A(n_2185),
.B(n_1785),
.C(n_1867),
.Y(n_2191)
);

INVx2_ASAP7_75t_SL g2192 ( 
.A(n_2181),
.Y(n_2192)
);

INVxp67_ASAP7_75t_L g2193 ( 
.A(n_2190),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2189),
.B(n_2182),
.Y(n_2194)
);

BUFx2_ASAP7_75t_L g2195 ( 
.A(n_2192),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2191),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2195),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2193),
.B(n_2187),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2194),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2196),
.Y(n_2200)
);

OAI21xp33_ASAP7_75t_SL g2201 ( 
.A1(n_2194),
.A2(n_2186),
.B(n_2183),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2195),
.Y(n_2202)
);

INVxp67_ASAP7_75t_SL g2203 ( 
.A(n_2197),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2198),
.Y(n_2204)
);

OAI32xp33_ASAP7_75t_L g2205 ( 
.A1(n_2201),
.A2(n_2184),
.A3(n_2188),
.B1(n_2175),
.B2(n_2083),
.Y(n_2205)
);

O2A1O1Ixp33_ASAP7_75t_SL g2206 ( 
.A1(n_2202),
.A2(n_2199),
.B(n_2200),
.C(n_2201),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2197),
.B(n_2188),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2197),
.Y(n_2208)
);

INVxp67_ASAP7_75t_SL g2209 ( 
.A(n_2197),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2197),
.B(n_2036),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2201),
.A2(n_1911),
.B(n_1893),
.Y(n_2211)
);

NAND4xp75_ASAP7_75t_L g2212 ( 
.A(n_2201),
.B(n_1755),
.C(n_1795),
.D(n_1843),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_2204),
.Y(n_2213)
);

OR2x2_ASAP7_75t_L g2214 ( 
.A(n_2203),
.B(n_2209),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2207),
.B(n_2069),
.Y(n_2215)
);

OAI21x1_ASAP7_75t_L g2216 ( 
.A1(n_2208),
.A2(n_1847),
.B(n_1965),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2206),
.Y(n_2217)
);

INVx1_ASAP7_75t_SL g2218 ( 
.A(n_2212),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2210),
.B(n_2125),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2211),
.Y(n_2220)
);

CKINVDCx20_ASAP7_75t_L g2221 ( 
.A(n_2205),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2211),
.B(n_2139),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2203),
.B(n_2054),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2204),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2204),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_2214),
.B(n_2128),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2213),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2221),
.A2(n_1800),
.B1(n_1790),
.B2(n_2146),
.Y(n_2228)
);

NAND2x1_ASAP7_75t_L g2229 ( 
.A(n_2223),
.B(n_2128),
.Y(n_2229)
);

AOI221xp5_ASAP7_75t_L g2230 ( 
.A1(n_2217),
.A2(n_1852),
.B1(n_1974),
.B2(n_2146),
.C(n_2080),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_2220),
.A2(n_2133),
.B1(n_2132),
.B2(n_2090),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2220),
.B(n_1790),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2217),
.B(n_2126),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2224),
.B(n_2054),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2215),
.Y(n_2235)
);

OAI211xp5_ASAP7_75t_L g2236 ( 
.A1(n_2225),
.A2(n_2010),
.B(n_1873),
.C(n_1879),
.Y(n_2236)
);

OAI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2218),
.A2(n_1769),
.B1(n_2023),
.B2(n_1876),
.C(n_1898),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2219),
.B(n_2126),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2222),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2227),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_2229),
.Y(n_2241)
);

AOI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2239),
.A2(n_2216),
.B1(n_2008),
.B2(n_1984),
.C(n_1987),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2234),
.Y(n_2243)
);

INVx1_ASAP7_75t_SL g2244 ( 
.A(n_2226),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2235),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2233),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2238),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2232),
.B(n_2136),
.Y(n_2248)
);

AOI21xp33_ASAP7_75t_SL g2249 ( 
.A1(n_2228),
.A2(n_219),
.B(n_220),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2237),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2236),
.B(n_2230),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_L g2252 ( 
.A(n_2231),
.B(n_2136),
.Y(n_2252)
);

INVx1_ASAP7_75t_SL g2253 ( 
.A(n_2227),
.Y(n_2253)
);

INVx1_ASAP7_75t_SL g2254 ( 
.A(n_2253),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2241),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2253),
.B(n_2064),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2240),
.Y(n_2257)
);

INVx1_ASAP7_75t_SL g2258 ( 
.A(n_2244),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2245),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2246),
.B(n_2130),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2248),
.B(n_2027),
.Y(n_2261)
);

NAND2x1_ASAP7_75t_L g2262 ( 
.A(n_2247),
.B(n_2026),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2243),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2249),
.B(n_2041),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_L g2265 ( 
.A(n_2252),
.B(n_1875),
.Y(n_2265)
);

INVx2_ASAP7_75t_SL g2266 ( 
.A(n_2250),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2251),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2242),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2253),
.B(n_2129),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2253),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2253),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2253),
.B(n_2130),
.Y(n_2272)
);

INVx3_ASAP7_75t_L g2273 ( 
.A(n_2253),
.Y(n_2273)
);

INVxp67_ASAP7_75t_L g2274 ( 
.A(n_2246),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2273),
.Y(n_2275)
);

NAND4xp75_ASAP7_75t_L g2276 ( 
.A(n_2270),
.B(n_1918),
.C(n_1901),
.D(n_1895),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2273),
.B(n_2129),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2254),
.Y(n_2278)
);

NAND3xp33_ASAP7_75t_SL g2279 ( 
.A(n_2271),
.B(n_2258),
.C(n_2259),
.Y(n_2279)
);

AOI221xp5_ASAP7_75t_L g2280 ( 
.A1(n_2267),
.A2(n_1978),
.B1(n_2132),
.B2(n_2133),
.C(n_2134),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_L g2281 ( 
.A(n_2255),
.B(n_2274),
.C(n_2257),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2261),
.B(n_2027),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2256),
.B(n_2031),
.Y(n_2283)
);

NAND4xp25_ASAP7_75t_L g2284 ( 
.A(n_2263),
.B(n_221),
.C(n_219),
.D(n_220),
.Y(n_2284)
);

NAND4xp25_ASAP7_75t_L g2285 ( 
.A(n_2265),
.B(n_224),
.C(n_222),
.D(n_223),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2272),
.Y(n_2286)
);

INVxp67_ASAP7_75t_SL g2287 ( 
.A(n_2266),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2260),
.A2(n_2128),
.B1(n_2134),
.B2(n_2048),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2269),
.Y(n_2289)
);

NOR3x1_ASAP7_75t_L g2290 ( 
.A(n_2262),
.B(n_222),
.C(n_223),
.Y(n_2290)
);

NAND4xp25_ASAP7_75t_L g2291 ( 
.A(n_2268),
.B(n_224),
.C(n_2042),
.D(n_1925),
.Y(n_2291)
);

NAND4xp25_ASAP7_75t_L g2292 ( 
.A(n_2264),
.B(n_2043),
.C(n_2092),
.D(n_2103),
.Y(n_2292)
);

AOI322xp5_ASAP7_75t_L g2293 ( 
.A1(n_2254),
.A2(n_2133),
.A3(n_2116),
.B1(n_2051),
.B2(n_2117),
.C1(n_1803),
.C2(n_1849),
.Y(n_2293)
);

INVxp67_ASAP7_75t_L g2294 ( 
.A(n_2273),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_L g2295 ( 
.A(n_2273),
.B(n_2039),
.Y(n_2295)
);

NAND4xp25_ASAP7_75t_L g2296 ( 
.A(n_2258),
.B(n_2043),
.C(n_2103),
.D(n_2117),
.Y(n_2296)
);

OAI221xp5_ASAP7_75t_SL g2297 ( 
.A1(n_2254),
.A2(n_2033),
.B1(n_2120),
.B2(n_2048),
.C(n_2039),
.Y(n_2297)
);

AOI22xp5_ASAP7_75t_SL g2298 ( 
.A1(n_2273),
.A2(n_2062),
.B1(n_1835),
.B2(n_2128),
.Y(n_2298)
);

OAI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2254),
.A2(n_2128),
.B1(n_2061),
.B2(n_2129),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_L g2300 ( 
.A(n_2273),
.B(n_2129),
.C(n_2052),
.Y(n_2300)
);

OAI211xp5_ASAP7_75t_L g2301 ( 
.A1(n_2258),
.A2(n_1964),
.B(n_2015),
.C(n_1991),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2273),
.B(n_2090),
.Y(n_2302)
);

NAND2x1_ASAP7_75t_L g2303 ( 
.A(n_2273),
.B(n_1835),
.Y(n_2303)
);

AOI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2258),
.A2(n_2025),
.B(n_2019),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2273),
.Y(n_2305)
);

AOI211xp5_ASAP7_75t_L g2306 ( 
.A1(n_2254),
.A2(n_1973),
.B(n_1975),
.C(n_2060),
.Y(n_2306)
);

NOR3xp33_ASAP7_75t_SL g2307 ( 
.A(n_2270),
.B(n_2061),
.C(n_293),
.Y(n_2307)
);

OR2x2_ASAP7_75t_L g2308 ( 
.A(n_2279),
.B(n_2086),
.Y(n_2308)
);

NOR3xp33_ASAP7_75t_L g2309 ( 
.A(n_2281),
.B(n_1869),
.C(n_2098),
.Y(n_2309)
);

NAND3x1_ASAP7_75t_L g2310 ( 
.A(n_2305),
.B(n_2058),
.C(n_2046),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2275),
.B(n_2060),
.Y(n_2311)
);

AND4x1_ASAP7_75t_L g2312 ( 
.A(n_2290),
.B(n_1835),
.C(n_2033),
.D(n_297),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_2294),
.B(n_2060),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2287),
.Y(n_2314)
);

NAND3xp33_ASAP7_75t_L g2315 ( 
.A(n_2278),
.B(n_2076),
.C(n_2111),
.Y(n_2315)
);

AOI21xp33_ASAP7_75t_SL g2316 ( 
.A1(n_2289),
.A2(n_295),
.B(n_296),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2286),
.Y(n_2317)
);

NOR2x1_ASAP7_75t_L g2318 ( 
.A(n_2284),
.B(n_2120),
.Y(n_2318)
);

NOR3xp33_ASAP7_75t_L g2319 ( 
.A(n_2295),
.B(n_1869),
.C(n_2098),
.Y(n_2319)
);

OAI221xp5_ASAP7_75t_SL g2320 ( 
.A1(n_2277),
.A2(n_2302),
.B1(n_2283),
.B2(n_2291),
.C(n_2282),
.Y(n_2320)
);

O2A1O1Ixp33_ASAP7_75t_L g2321 ( 
.A1(n_2307),
.A2(n_2120),
.B(n_2111),
.C(n_2086),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2285),
.B(n_2060),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2276),
.Y(n_2323)
);

NAND4xp75_ASAP7_75t_L g2324 ( 
.A(n_2280),
.B(n_2081),
.C(n_301),
.D(n_299),
.Y(n_2324)
);

NAND3xp33_ASAP7_75t_L g2325 ( 
.A(n_2303),
.B(n_2076),
.C(n_2071),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2292),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_2296),
.B(n_2071),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2288),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2300),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_SL g2330 ( 
.A(n_2297),
.B(n_2071),
.Y(n_2330)
);

AOI221x1_ASAP7_75t_L g2331 ( 
.A1(n_2299),
.A2(n_2046),
.B1(n_2044),
.B2(n_2058),
.C(n_2071),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2293),
.B(n_2076),
.Y(n_2332)
);

NOR3xp33_ASAP7_75t_L g2333 ( 
.A(n_2306),
.B(n_300),
.C(n_303),
.Y(n_2333)
);

O2A1O1Ixp33_ASAP7_75t_L g2334 ( 
.A1(n_2304),
.A2(n_2084),
.B(n_2029),
.C(n_2081),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2298),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2312),
.B(n_2301),
.Y(n_2336)
);

NOR3xp33_ASAP7_75t_L g2337 ( 
.A(n_2314),
.B(n_304),
.C(n_305),
.Y(n_2337)
);

NOR2x1_ASAP7_75t_L g2338 ( 
.A(n_2317),
.B(n_2044),
.Y(n_2338)
);

AOI21x1_ASAP7_75t_L g2339 ( 
.A1(n_2323),
.A2(n_2328),
.B(n_2329),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_2311),
.B(n_2122),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2311),
.Y(n_2341)
);

OR2x2_ASAP7_75t_L g2342 ( 
.A(n_2308),
.B(n_2029),
.Y(n_2342)
);

AOI222xp33_ASAP7_75t_L g2343 ( 
.A1(n_2335),
.A2(n_2326),
.B1(n_2313),
.B2(n_2327),
.C1(n_2332),
.C2(n_2322),
.Y(n_2343)
);

AOI221xp5_ASAP7_75t_L g2344 ( 
.A1(n_2320),
.A2(n_2084),
.B1(n_2122),
.B2(n_1764),
.C(n_1799),
.Y(n_2344)
);

INVx1_ASAP7_75t_SL g2345 ( 
.A(n_2324),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2316),
.B(n_2318),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2333),
.B(n_2109),
.Y(n_2347)
);

OR2x2_ASAP7_75t_L g2348 ( 
.A(n_2315),
.B(n_2095),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2325),
.B(n_2095),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2330),
.B(n_2105),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2309),
.A2(n_2105),
.B1(n_2122),
.B2(n_2040),
.Y(n_2351)
);

XOR2x2_ASAP7_75t_L g2352 ( 
.A(n_2310),
.B(n_309),
.Y(n_2352)
);

CKINVDCx14_ASAP7_75t_R g2353 ( 
.A(n_2321),
.Y(n_2353)
);

INVxp67_ASAP7_75t_L g2354 ( 
.A(n_2331),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2334),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2319),
.B(n_310),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2314),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2312),
.B(n_311),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2311),
.Y(n_2359)
);

AOI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2314),
.A2(n_2040),
.B(n_2104),
.Y(n_2360)
);

INVx1_ASAP7_75t_SL g2361 ( 
.A(n_2314),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2312),
.B(n_313),
.Y(n_2362)
);

INVx1_ASAP7_75t_SL g2363 ( 
.A(n_2314),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2314),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2314),
.Y(n_2365)
);

OR2x2_ASAP7_75t_L g2366 ( 
.A(n_2314),
.B(n_314),
.Y(n_2366)
);

OAI211xp5_ASAP7_75t_L g2367 ( 
.A1(n_2314),
.A2(n_2040),
.B(n_322),
.C(n_315),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2314),
.Y(n_2368)
);

OAI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_2308),
.A2(n_2105),
.B1(n_2063),
.B2(n_2057),
.Y(n_2369)
);

INVxp67_ASAP7_75t_L g2370 ( 
.A(n_2358),
.Y(n_2370)
);

NAND4xp25_ASAP7_75t_L g2371 ( 
.A(n_2343),
.B(n_327),
.C(n_318),
.D(n_326),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2339),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2366),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2361),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2363),
.Y(n_2375)
);

NOR2x1_ASAP7_75t_L g2376 ( 
.A(n_2357),
.B(n_330),
.Y(n_2376)
);

AO22x2_ASAP7_75t_L g2377 ( 
.A1(n_2341),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2359),
.B(n_335),
.Y(n_2378)
);

AOI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2364),
.A2(n_1799),
.B1(n_1884),
.B2(n_1904),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2365),
.A2(n_1884),
.B1(n_1905),
.B2(n_2072),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2368),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2352),
.B(n_336),
.Y(n_2382)
);

AOI22xp33_ASAP7_75t_L g2383 ( 
.A1(n_2353),
.A2(n_2345),
.B1(n_2362),
.B2(n_2336),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2346),
.B(n_337),
.Y(n_2384)
);

A2O1A1Ixp33_ASAP7_75t_SL g2385 ( 
.A1(n_2354),
.A2(n_339),
.B(n_340),
.C(n_342),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2338),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2342),
.Y(n_2387)
);

OA22x2_ASAP7_75t_L g2388 ( 
.A1(n_2355),
.A2(n_2104),
.B1(n_2063),
.B2(n_2057),
.Y(n_2388)
);

NOR2x1_ASAP7_75t_L g2389 ( 
.A(n_2367),
.B(n_343),
.Y(n_2389)
);

A2O1A1Ixp33_ASAP7_75t_SL g2390 ( 
.A1(n_2350),
.A2(n_345),
.B(n_346),
.C(n_348),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2356),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2340),
.B(n_349),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2348),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2337),
.B(n_2369),
.Y(n_2394)
);

AO22x1_ASAP7_75t_L g2395 ( 
.A1(n_2347),
.A2(n_1884),
.B1(n_351),
.B2(n_352),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2372),
.Y(n_2396)
);

NOR2x1p5_ASAP7_75t_L g2397 ( 
.A(n_2374),
.B(n_2349),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2375),
.B(n_2381),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2373),
.Y(n_2399)
);

NAND3xp33_ASAP7_75t_L g2400 ( 
.A(n_2383),
.B(n_2344),
.C(n_2360),
.Y(n_2400)
);

OA21x2_ASAP7_75t_L g2401 ( 
.A1(n_2386),
.A2(n_2351),
.B(n_350),
.Y(n_2401)
);

AOI22xp5_ASAP7_75t_L g2402 ( 
.A1(n_2370),
.A2(n_2082),
.B1(n_2072),
.B2(n_1951),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2382),
.B(n_353),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2395),
.B(n_354),
.Y(n_2404)
);

NAND3x1_ASAP7_75t_SL g2405 ( 
.A(n_2376),
.B(n_355),
.C(n_356),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2387),
.B(n_357),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2389),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2393),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2392),
.Y(n_2409)
);

XNOR2x2_ASAP7_75t_L g2410 ( 
.A(n_2384),
.B(n_359),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2391),
.B(n_2082),
.Y(n_2411)
);

OAI31xp33_ASAP7_75t_L g2412 ( 
.A1(n_2385),
.A2(n_2063),
.A3(n_2057),
.B(n_363),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2378),
.B(n_518),
.Y(n_2413)
);

NOR2x1_ASAP7_75t_L g2414 ( 
.A(n_2371),
.B(n_360),
.Y(n_2414)
);

INVx1_ASAP7_75t_SL g2415 ( 
.A(n_2394),
.Y(n_2415)
);

NAND2xp33_ASAP7_75t_SL g2416 ( 
.A(n_2390),
.B(n_361),
.Y(n_2416)
);

OR2x2_ASAP7_75t_L g2417 ( 
.A(n_2380),
.B(n_364),
.Y(n_2417)
);

AND3x4_ASAP7_75t_L g2418 ( 
.A(n_2377),
.B(n_2379),
.C(n_2388),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2377),
.B(n_517),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2372),
.Y(n_2420)
);

NOR2xp33_ASAP7_75t_L g2421 ( 
.A(n_2372),
.B(n_368),
.Y(n_2421)
);

INVx1_ASAP7_75t_SL g2422 ( 
.A(n_2372),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2372),
.Y(n_2423)
);

INVx3_ASAP7_75t_L g2424 ( 
.A(n_2398),
.Y(n_2424)
);

NAND4xp75_ASAP7_75t_L g2425 ( 
.A(n_2407),
.B(n_369),
.C(n_370),
.D(n_371),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2415),
.B(n_372),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2422),
.B(n_373),
.Y(n_2427)
);

AND5x1_ASAP7_75t_L g2428 ( 
.A(n_2412),
.B(n_375),
.C(n_377),
.D(n_379),
.E(n_380),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2408),
.B(n_381),
.Y(n_2429)
);

NAND5xp2_ASAP7_75t_L g2430 ( 
.A(n_2396),
.B(n_513),
.C(n_383),
.D(n_385),
.E(n_386),
.Y(n_2430)
);

INVxp67_ASAP7_75t_L g2431 ( 
.A(n_2419),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2410),
.Y(n_2432)
);

HB1xp67_ASAP7_75t_L g2433 ( 
.A(n_2399),
.Y(n_2433)
);

OAI211xp5_ASAP7_75t_SL g2434 ( 
.A1(n_2420),
.A2(n_382),
.B(n_387),
.C(n_388),
.Y(n_2434)
);

NAND4xp25_ASAP7_75t_SL g2435 ( 
.A(n_2423),
.B(n_389),
.C(n_390),
.D(n_391),
.Y(n_2435)
);

AOI221xp5_ASAP7_75t_L g2436 ( 
.A1(n_2400),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.C(n_397),
.Y(n_2436)
);

NAND5xp2_ASAP7_75t_L g2437 ( 
.A(n_2409),
.B(n_512),
.C(n_400),
.D(n_403),
.E(n_404),
.Y(n_2437)
);

NOR2xp33_ASAP7_75t_L g2438 ( 
.A(n_2403),
.B(n_398),
.Y(n_2438)
);

NOR4xp75_ASAP7_75t_L g2439 ( 
.A(n_2404),
.B(n_405),
.C(n_407),
.D(n_408),
.Y(n_2439)
);

NOR2x1_ASAP7_75t_L g2440 ( 
.A(n_2397),
.B(n_409),
.Y(n_2440)
);

NAND4xp25_ASAP7_75t_SL g2441 ( 
.A(n_2414),
.B(n_410),
.C(n_412),
.D(n_413),
.Y(n_2441)
);

NOR3x2_ASAP7_75t_L g2442 ( 
.A(n_2424),
.B(n_2417),
.C(n_2405),
.Y(n_2442)
);

NOR3xp33_ASAP7_75t_SL g2443 ( 
.A(n_2432),
.B(n_2421),
.C(n_2416),
.Y(n_2443)
);

INVx1_ASAP7_75t_SL g2444 ( 
.A(n_2433),
.Y(n_2444)
);

NAND4xp75_ASAP7_75t_L g2445 ( 
.A(n_2440),
.B(n_2401),
.C(n_2406),
.D(n_2413),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2424),
.Y(n_2446)
);

AOI22xp33_ASAP7_75t_SL g2447 ( 
.A1(n_2427),
.A2(n_2401),
.B1(n_2411),
.B2(n_2418),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2429),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2425),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_2431),
.B(n_2402),
.Y(n_2450)
);

NAND3x1_ASAP7_75t_L g2451 ( 
.A(n_2426),
.B(n_414),
.C(n_418),
.Y(n_2451)
);

NOR3x2_ASAP7_75t_L g2452 ( 
.A(n_2428),
.B(n_420),
.C(n_423),
.Y(n_2452)
);

NOR3xp33_ASAP7_75t_SL g2453 ( 
.A(n_2441),
.B(n_424),
.C(n_425),
.Y(n_2453)
);

NOR4xp25_ASAP7_75t_L g2454 ( 
.A(n_2444),
.B(n_2438),
.C(n_2434),
.D(n_2435),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2446),
.B(n_2436),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2452),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_SL g2457 ( 
.A1(n_2447),
.A2(n_2439),
.B1(n_2430),
.B2(n_2437),
.Y(n_2457)
);

INVx2_ASAP7_75t_SL g2458 ( 
.A(n_2448),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2445),
.B(n_426),
.Y(n_2459)
);

OR2x2_ASAP7_75t_L g2460 ( 
.A(n_2449),
.B(n_428),
.Y(n_2460)
);

NOR3xp33_ASAP7_75t_L g2461 ( 
.A(n_2450),
.B(n_429),
.C(n_431),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2458),
.Y(n_2462)
);

AND2x4_ASAP7_75t_L g2463 ( 
.A(n_2456),
.B(n_2443),
.Y(n_2463)
);

NAND4xp75_ASAP7_75t_L g2464 ( 
.A(n_2455),
.B(n_2453),
.C(n_2442),
.D(n_2454),
.Y(n_2464)
);

BUFx2_ASAP7_75t_L g2465 ( 
.A(n_2457),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2462),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2465),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_SL g2468 ( 
.A(n_2464),
.B(n_2463),
.Y(n_2468)
);

BUFx2_ASAP7_75t_L g2469 ( 
.A(n_2466),
.Y(n_2469)
);

AND2x2_ASAP7_75t_SL g2470 ( 
.A(n_2468),
.B(n_2459),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2467),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2467),
.A2(n_2460),
.B(n_2461),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2469),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2471),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2470),
.Y(n_2475)
);

OAI22xp5_ASAP7_75t_SL g2476 ( 
.A1(n_2473),
.A2(n_2472),
.B1(n_2451),
.B2(n_434),
.Y(n_2476)
);

OAI22xp33_ASAP7_75t_L g2477 ( 
.A1(n_2476),
.A2(n_2475),
.B1(n_2474),
.B2(n_439),
.Y(n_2477)
);

AOI21xp5_ASAP7_75t_L g2478 ( 
.A1(n_2477),
.A2(n_432),
.B(n_433),
.Y(n_2478)
);

AOI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2478),
.A2(n_440),
.B1(n_443),
.B2(n_445),
.Y(n_2479)
);

AOI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2479),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.Y(n_2480)
);

OAI21x1_ASAP7_75t_L g2481 ( 
.A1(n_2480),
.A2(n_449),
.B(n_450),
.Y(n_2481)
);

AOI322xp5_ASAP7_75t_L g2482 ( 
.A1(n_2481),
.A2(n_451),
.A3(n_452),
.B1(n_453),
.B2(n_457),
.C1(n_458),
.C2(n_460),
.Y(n_2482)
);

AOI22xp5_ASAP7_75t_L g2483 ( 
.A1(n_2482),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_2483)
);

O2A1O1Ixp33_ASAP7_75t_L g2484 ( 
.A1(n_2483),
.A2(n_465),
.B(n_466),
.C(n_468),
.Y(n_2484)
);

AOI211xp5_ASAP7_75t_L g2485 ( 
.A1(n_2484),
.A2(n_469),
.B(n_470),
.C(n_472),
.Y(n_2485)
);


endmodule