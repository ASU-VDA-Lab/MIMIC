module fake_netlist_1_7973_n_34 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
INVx4_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_0), .B(n_4), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_15), .B(n_0), .Y(n_20) );
NOR3xp33_ASAP7_75t_SL g21 ( .A(n_16), .B(n_1), .C(n_5), .Y(n_21) );
BUFx4f_ASAP7_75t_SL g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_19), .B(n_17), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
OAI31xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_23), .A3(n_16), .B(n_22), .Y(n_26) );
AOI21xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_18), .B(n_14), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g29 ( .A(n_27), .B(n_1), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
AOI22xp33_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_15), .B1(n_21), .B2(n_9), .Y(n_31) );
NAND3xp33_ASAP7_75t_SL g32 ( .A(n_30), .B(n_6), .C(n_8), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
AOI22xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_31), .B1(n_10), .B2(n_12), .Y(n_34) );
endmodule