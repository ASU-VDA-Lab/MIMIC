module fake_jpeg_19299_n_290 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_18),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_24),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_44),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_52),
.B1(n_61),
.B2(n_25),
.Y(n_73)
);

CKINVDCx9p33_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_24),
.B1(n_29),
.B2(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_67),
.B1(n_72),
.B2(n_41),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_42),
.C(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_70),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_27),
.B1(n_40),
.B2(n_28),
.Y(n_67)
);

O2A1O1Ixp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_42),
.B(n_35),
.C(n_30),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_78),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_42),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_32),
.B1(n_26),
.B2(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_54),
.B1(n_41),
.B2(n_43),
.Y(n_112)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_88),
.Y(n_110)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_95),
.B1(n_25),
.B2(n_77),
.Y(n_115)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_71),
.Y(n_104)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_69),
.B1(n_70),
.B2(n_66),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_62),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_77),
.B1(n_57),
.B2(n_68),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_38),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_25),
.B1(n_43),
.B2(n_58),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_64),
.B(n_70),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_118),
.B(n_94),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_96),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_64),
.B(n_79),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_111),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_72),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_122),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_19),
.B(n_23),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_82),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_93),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_17),
.B(n_15),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_34),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_54),
.B1(n_77),
.B2(n_56),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_121),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_125),
.B(n_126),
.Y(n_172)
);

CKINVDCx12_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_129),
.B(n_133),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_105),
.C(n_104),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_14),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_R g137 ( 
.A(n_111),
.B(n_84),
.Y(n_137)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_16),
.B1(n_14),
.B2(n_20),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_98),
.B(n_97),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_139),
.B(n_143),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_115),
.B(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_84),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_87),
.C(n_34),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_55),
.C(n_34),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_92),
.B(n_19),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_83),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_44),
.B(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_148),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_13),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_101),
.A2(n_15),
.B(n_21),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_20),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_132),
.B(n_134),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_138),
.B(n_145),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_171),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_116),
.C(n_123),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_166),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_142),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_103),
.A3(n_57),
.B1(n_34),
.B2(n_17),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_81),
.B1(n_103),
.B2(n_21),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_179),
.B(n_180),
.Y(n_205)
);

AOI31xp33_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_17),
.A3(n_21),
.B(n_20),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_55),
.C(n_33),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_139),
.C(n_129),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_14),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_176),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_143),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_151),
.B(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_17),
.B1(n_12),
.B2(n_20),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_181),
.B(n_20),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_201),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_205),
.B1(n_155),
.B2(n_174),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_154),
.B1(n_144),
.B2(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_129),
.C(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_199),
.C(n_204),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_147),
.B1(n_131),
.B2(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_131),
.B1(n_152),
.B2(n_81),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_195),
.B1(n_178),
.B2(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_202),
.B(n_156),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_55),
.C(n_51),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_23),
.B1(n_12),
.B2(n_10),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_195),
.B1(n_192),
.B2(n_183),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_55),
.B(n_20),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_51),
.C(n_49),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_165),
.C(n_169),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_216),
.C(n_218),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_223),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_181),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_221),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_158),
.C(n_175),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_164),
.C(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_184),
.B(n_166),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_185),
.A2(n_160),
.B1(n_23),
.B2(n_12),
.Y(n_221)
);

OAI31xp33_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_198),
.A3(n_202),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_208),
.B(n_214),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_194),
.B1(n_198),
.B2(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_234),
.B1(n_213),
.B2(n_220),
.Y(n_240)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_201),
.B1(n_197),
.B2(n_49),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_33),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_39),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_10),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_0),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_206),
.C(n_220),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_11),
.C(n_33),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_231),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_206),
.B1(n_20),
.B2(n_14),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_246),
.B1(n_236),
.B2(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_33),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_249),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_235),
.C(n_239),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_14),
.B(n_13),
.C(n_4),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_229),
.B(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_257),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_231),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_33),
.C(n_11),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_238),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_233),
.C(n_33),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_16),
.Y(n_267)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_0),
.Y(n_264)
);

AOI21x1_ASAP7_75t_SL g266 ( 
.A1(n_256),
.A2(n_247),
.B(n_249),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_274),
.B(n_255),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_272),
.B(n_268),
.C(n_265),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_11),
.B1(n_13),
.B2(n_22),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_22),
.B(n_13),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_273),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_253),
.A2(n_22),
.B(n_16),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_261),
.B(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_278),
.B(n_16),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_16),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_33),
.B1(n_4),
.B2(n_5),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_3),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_283),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_7),
.C2(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_276),
.C(n_280),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_285),
.B(n_7),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_7),
.C(n_8),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_8),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_9),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_9),
.Y(n_290)
);


endmodule