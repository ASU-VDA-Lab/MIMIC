module fake_jpeg_14905_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_17),
.B1(n_8),
.B2(n_13),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_17)
);

O2A1O1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_27),
.Y(n_28)
);

CKINVDCx6p67_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_18),
.B(n_20),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_40),
.B(n_25),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_31),
.B(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_36),
.B1(n_39),
.B2(n_25),
.Y(n_47)
);

XOR2x2_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_38),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_42),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_12),
.B1(n_7),
.B2(n_10),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_SL g53 ( 
.A(n_52),
.B(n_15),
.C(n_12),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_15),
.Y(n_54)
);


endmodule