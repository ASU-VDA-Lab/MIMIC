module fake_jpeg_22787_n_58 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_58);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_5),
.B(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_35),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_35),
.B1(n_36),
.B2(n_23),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_23),
.A2(n_30),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_41),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_39),
.B(n_50),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_46),
.B1(n_42),
.B2(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_42),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_27),
.Y(n_54)
);

OAI21x1_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B(n_43),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_40),
.B(n_45),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_44),
.B(n_29),
.Y(n_57)
);

AOI221xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_18),
.B1(n_22),
.B2(n_19),
.C(n_46),
.Y(n_58)
);


endmodule