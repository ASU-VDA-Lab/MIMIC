module fake_jpeg_2453_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx13_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_28),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_35),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_38),
.B(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_57),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_40),
.B(n_33),
.C(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_49),
.B1(n_43),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_43),
.B1(n_34),
.B2(n_36),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_59),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_37),
.B(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_20),
.B(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_34),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_43),
.C(n_38),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_76),
.C(n_80),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_54),
.B(n_33),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_83),
.B(n_3),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_33),
.C(n_15),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_30),
.C(n_29),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_3),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_92),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_71),
.B1(n_77),
.B2(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_5),
.B(n_9),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_97),
.C(n_4),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_4),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_103),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_106),
.B1(n_88),
.B2(n_12),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_94),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_85),
.C(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_106),
.B(n_104),
.C(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_115),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_99),
.B(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_110),
.C(n_111),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_118),
.B(n_116),
.Y(n_119)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_109),
.B(n_107),
.C(n_17),
.D(n_16),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_18),
.A3(n_21),
.B1(n_107),
.B2(n_11),
.C1(n_13),
.C2(n_14),
.Y(n_121)
);


endmodule