module fake_netlist_6_2864_n_1052 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1052);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1052;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_989;
wire n_843;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_87),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_79),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_107),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_45),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_47),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_99),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_52),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_74),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_7),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_55),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_34),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_119),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_97),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_2),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_130),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_75),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_33),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_81),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_51),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_104),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_59),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_145),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_68),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_183),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_144),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_169),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_129),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_50),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_116),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_91),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_100),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_39),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_53),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_30),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_16),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_1),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_203),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_153),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_184),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_58),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_69),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_201),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_26),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_215),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_209),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_140),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_28),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_205),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_174),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_10),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_106),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_185),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_18),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_40),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_66),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_105),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_29),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_110),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_148),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_77),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_57),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_216),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_22),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_131),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_175),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_90),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_30),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_137),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_76),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_141),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_167),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_128),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_115),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_89),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_31),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_22),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_154),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_126),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_158),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_272),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_234),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_244),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_256),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_225),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_248),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_226),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_263),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_227),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_240),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_228),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_284),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_230),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_233),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_231),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_232),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_0),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_270),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_285),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_247),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_238),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_261),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_236),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_242),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_247),
.B(n_0),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_241),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_246),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_288),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_291),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_245),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_251),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_302),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_254),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_304),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_315),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_R g372 ( 
.A(n_319),
.B(n_1),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_316),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_273),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_320),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_323),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_331),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_327),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_229),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_336),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_260),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_237),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_338),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_341),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_346),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g397 ( 
.A(n_324),
.B(n_300),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_348),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_349),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_327),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_357),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_358),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_R g407 ( 
.A(n_324),
.B(n_367),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_354),
.A2(n_312),
.B(n_257),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_361),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_321),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_374),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_356),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_367),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_370),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_351),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_322),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_330),
.B(n_312),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_387),
.B(n_255),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_388),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_386),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_264),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_363),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_387),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_292),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_411),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_292),
.Y(n_452)
);

OR2x6_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_258),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_268),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_382),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_259),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_389),
.B(n_301),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_412),
.B(n_389),
.Y(n_460)
);

INVx8_ASAP7_75t_L g461 ( 
.A(n_428),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_397),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_379),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_389),
.B(n_250),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_413),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_397),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_409),
.A2(n_267),
.B1(n_286),
.B2(n_299),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_384),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_419),
.B(n_424),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_425),
.B(n_239),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_409),
.A2(n_429),
.B1(n_269),
.B2(n_275),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_392),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_426),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_252),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_404),
.B(n_262),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_265),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_403),
.B(n_266),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_422),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_429),
.B(n_274),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_378),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_407),
.B(n_276),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_385),
.B(n_277),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_393),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_394),
.B(n_278),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_380),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_395),
.B(n_371),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_431),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_400),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_401),
.B(n_371),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_405),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_407),
.B(n_373),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_406),
.B(n_373),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_461),
.Y(n_511)
);

AOI221xp5_ASAP7_75t_L g512 ( 
.A1(n_439),
.A2(n_431),
.B1(n_433),
.B2(n_432),
.C(n_430),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_292),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_437),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_435),
.B(n_430),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_476),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_480),
.B(n_292),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_453),
.A2(n_477),
.B1(n_460),
.B2(n_496),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_455),
.B(n_417),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_507),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_460),
.B(n_311),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_448),
.B(n_430),
.Y(n_524)
);

NOR2x1p5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_420),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_443),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_461),
.A2(n_313),
.B(n_249),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_448),
.B(n_472),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_472),
.A2(n_292),
.B1(n_239),
.B2(n_249),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_461),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_453),
.A2(n_374),
.B1(n_420),
.B2(n_279),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_484),
.B(n_282),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_484),
.B(n_283),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_476),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_287),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_440),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_447),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_453),
.A2(n_298),
.B1(n_289),
.B2(n_290),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_496),
.B(n_462),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_465),
.B(n_293),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_500),
.A2(n_418),
.B1(n_402),
.B2(n_380),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_454),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_497),
.B(n_432),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_470),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_479),
.Y(n_545)
);

BUFx8_ASAP7_75t_L g546 ( 
.A(n_509),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_465),
.B(n_294),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_465),
.B(n_471),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_489),
.B(n_292),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_459),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_479),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_458),
.B(n_432),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_489),
.B(n_239),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_491),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_L g555 ( 
.A(n_478),
.B(n_295),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_447),
.B(n_432),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_471),
.B(n_481),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_471),
.B(n_481),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_468),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_471),
.B(n_297),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_502),
.B(n_418),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_503),
.Y(n_563)
);

NOR2x1p5_ASAP7_75t_L g564 ( 
.A(n_498),
.B(n_505),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_453),
.A2(n_309),
.B1(n_317),
.B2(n_314),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_475),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_505),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_477),
.A2(n_310),
.B1(n_308),
.B2(n_305),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_501),
.A2(n_402),
.B1(n_249),
.B2(n_239),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_491),
.Y(n_570)
);

OAI221xp5_ASAP7_75t_L g571 ( 
.A1(n_494),
.A2(n_249),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_449),
.A2(n_112),
.B1(n_223),
.B2(n_222),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_481),
.B(n_32),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_507),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_481),
.B(n_36),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_507),
.B(n_2),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_483),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_507),
.B(n_3),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_485),
.Y(n_579)
);

NOR2xp67_ASAP7_75t_L g580 ( 
.A(n_507),
.B(n_37),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_457),
.B(n_38),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_499),
.B(n_4),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_498),
.B(n_508),
.Y(n_583)
);

AOI221xp5_ASAP7_75t_L g584 ( 
.A1(n_501),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_441),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_456),
.B(n_41),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_SL g587 ( 
.A(n_482),
.B(n_6),
.C(n_8),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_498),
.B(n_42),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_487),
.B(n_43),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_510),
.B(n_9),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_457),
.B(n_44),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_504),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_467),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_441),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_528),
.A2(n_510),
.B1(n_493),
.B2(n_492),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_518),
.B(n_449),
.Y(n_596)
);

AOI21x1_ASAP7_75t_L g597 ( 
.A1(n_540),
.A2(n_488),
.B(n_486),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_511),
.A2(n_530),
.B(n_522),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_522),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_522),
.Y(n_600)
);

O2A1O1Ixp5_ASAP7_75t_L g601 ( 
.A1(n_523),
.A2(n_490),
.B(n_434),
.C(n_463),
.Y(n_601)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_547),
.A2(n_463),
.B(n_450),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_582),
.A2(n_452),
.B1(n_434),
.B2(n_492),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_516),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_511),
.A2(n_464),
.B(n_436),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_543),
.B(n_452),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_530),
.A2(n_464),
.B(n_436),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_586),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_524),
.B(n_434),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_534),
.Y(n_610)
);

AOI21x1_ASAP7_75t_L g611 ( 
.A1(n_548),
.A2(n_450),
.B(n_445),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_544),
.B(n_504),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_557),
.A2(n_464),
.B(n_436),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_558),
.A2(n_446),
.B(n_444),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_567),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_581),
.A2(n_451),
.B(n_456),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_514),
.B(n_466),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_586),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_537),
.Y(n_619)
);

NOR2x1_ASAP7_75t_L g620 ( 
.A(n_539),
.B(n_506),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_L g621 ( 
.A(n_519),
.B(n_495),
.C(n_469),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_581),
.A2(n_469),
.B(n_466),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_562),
.B(n_473),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_520),
.B(n_442),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_591),
.A2(n_442),
.B(n_473),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_545),
.A2(n_478),
.B(n_473),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_513),
.A2(n_478),
.B(n_124),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_515),
.B(n_12),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_561),
.B(n_13),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_591),
.A2(n_478),
.B(n_127),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_580),
.A2(n_478),
.B(n_125),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_536),
.B(n_14),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_583),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_551),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_541),
.B(n_478),
.C(n_16),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_529),
.A2(n_132),
.B1(n_219),
.B2(n_218),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_563),
.B(n_46),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_552),
.B(n_15),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_560),
.A2(n_133),
.B(n_217),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_532),
.A2(n_123),
.B(n_213),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_512),
.B(n_48),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_526),
.B(n_17),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_533),
.A2(n_122),
.B(n_212),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_535),
.A2(n_121),
.B(n_211),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_556),
.B(n_17),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_542),
.B(n_18),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_513),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_517),
.A2(n_134),
.B(n_210),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_549),
.A2(n_120),
.B(n_208),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_550),
.B(n_19),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_559),
.B(n_20),
.Y(n_653)
);

CKINVDCx8_ASAP7_75t_R g654 ( 
.A(n_556),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_566),
.B(n_21),
.Y(n_655)
);

AO22x1_ASAP7_75t_L g656 ( 
.A1(n_593),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_549),
.A2(n_136),
.B(n_207),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_553),
.A2(n_135),
.B(n_202),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_553),
.A2(n_118),
.B(n_200),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_634),
.B(n_531),
.Y(n_660)
);

OAI22x1_ASAP7_75t_L g661 ( 
.A1(n_612),
.A2(n_564),
.B1(n_525),
.B2(n_590),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_634),
.B(n_577),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_596),
.A2(n_517),
.B(n_588),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_608),
.B(n_537),
.Y(n_664)
);

AOI21xp33_ASAP7_75t_L g665 ( 
.A1(n_609),
.A2(n_579),
.B(n_569),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_624),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_630),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_606),
.A2(n_521),
.B(n_574),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_613),
.A2(n_575),
.B(n_573),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_625),
.Y(n_670)
);

AND3x1_ASAP7_75t_SL g671 ( 
.A(n_656),
.B(n_584),
.C(n_571),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_601),
.A2(n_554),
.B(n_585),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_608),
.B(n_594),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_622),
.A2(n_555),
.B(n_589),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_604),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_618),
.B(n_568),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_618),
.B(n_538),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_603),
.A2(n_654),
.B1(n_595),
.B2(n_620),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_605),
.A2(n_576),
.B(n_578),
.Y(n_679)
);

AO31x2_ASAP7_75t_L g680 ( 
.A1(n_595),
.A2(n_593),
.A3(n_527),
.B(n_572),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_607),
.A2(n_565),
.B(n_587),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_629),
.B(n_546),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_626),
.A2(n_598),
.B(n_616),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_599),
.B(n_592),
.Y(n_684)
);

O2A1O1Ixp5_ASAP7_75t_L g685 ( 
.A1(n_642),
.A2(n_546),
.B(n_138),
.C(n_139),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_647),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_610),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_602),
.A2(n_114),
.B(n_199),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_617),
.A2(n_113),
.B(n_198),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_627),
.A2(n_111),
.B(n_197),
.Y(n_690)
);

NOR2x1_ASAP7_75t_L g691 ( 
.A(n_619),
.B(n_49),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_619),
.B(n_54),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_633),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_628),
.A2(n_117),
.B(n_196),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_621),
.B(n_23),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_644),
.B(n_56),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_644),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_628),
.A2(n_224),
.B(n_142),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_599),
.A2(n_109),
.B1(n_194),
.B2(n_192),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_650),
.A2(n_108),
.B(n_191),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_639),
.B(n_643),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_25),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_650),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_SL g704 ( 
.A1(n_636),
.A2(n_27),
.B(n_31),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_635),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_599),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_652),
.B(n_63),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_614),
.A2(n_64),
.B(n_65),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_644),
.B(n_67),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_623),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_600),
.A2(n_70),
.B(n_71),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_600),
.A2(n_637),
.B(n_631),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_600),
.B(n_653),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_655),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_611),
.A2(n_72),
.B(n_73),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_597),
.A2(n_78),
.B(n_80),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_697),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_700),
.A2(n_649),
.B1(n_638),
.B2(n_657),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_667),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_664),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_696),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_714),
.B(n_615),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_664),
.B(n_651),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_710),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_666),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_687),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_698),
.B(n_646),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_705),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_662),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_663),
.A2(n_645),
.B(n_641),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_670),
.B(n_640),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_669),
.A2(n_632),
.B(n_658),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_698),
.A2(n_659),
.B1(n_83),
.B2(n_84),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_696),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_674),
.A2(n_82),
.B(n_85),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_701),
.B(n_86),
.Y(n_736)
);

AOI221x1_ASAP7_75t_L g737 ( 
.A1(n_703),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_686),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_675),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_660),
.B(n_195),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_667),
.B(n_95),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_693),
.B(n_96),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_694),
.A2(n_98),
.B(n_101),
.C(n_102),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_673),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_678),
.A2(n_677),
.B1(n_676),
.B2(n_713),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_682),
.B(n_190),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_695),
.B(n_103),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_692),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_692),
.Y(n_749)
);

INVx5_ASAP7_75t_L g750 ( 
.A(n_685),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_681),
.A2(n_143),
.B(n_146),
.C(n_147),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_712),
.A2(n_149),
.B(n_150),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_702),
.B(n_151),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_684),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_661),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_709),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_665),
.A2(n_159),
.B(n_160),
.C(n_162),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_704),
.B(n_163),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_690),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_707),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_668),
.A2(n_164),
.B(n_165),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_704),
.B(n_166),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_699),
.A2(n_706),
.B(n_689),
.C(n_679),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_691),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_716),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_680),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_672),
.B(n_189),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_708),
.A2(n_168),
.B(n_170),
.C(n_171),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_715),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_688),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_719),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_725),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_726),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_744),
.B(n_680),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_734),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_R g776 ( 
.A1(n_719),
.A2(n_671),
.B1(n_173),
.B2(n_177),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_728),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_758),
.A2(n_762),
.B1(n_740),
.B2(n_733),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_767),
.B(n_683),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_766),
.Y(n_780)
);

INVx4_ASAP7_75t_SL g781 ( 
.A(n_767),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_739),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_729),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_749),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_SL g785 ( 
.A1(n_758),
.A2(n_711),
.B1(n_680),
.B2(n_179),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_738),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_717),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_730),
.A2(n_172),
.B(n_178),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_770),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_723),
.Y(n_790)
);

OA21x2_ASAP7_75t_L g791 ( 
.A1(n_737),
.A2(n_732),
.B(n_731),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_769),
.Y(n_792)
);

AO21x2_ASAP7_75t_L g793 ( 
.A1(n_733),
.A2(n_180),
.B(n_181),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_748),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_724),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_734),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_L g797 ( 
.A1(n_758),
.A2(n_182),
.B1(n_187),
.B2(n_755),
.Y(n_797)
);

CKINVDCx11_ASAP7_75t_R g798 ( 
.A(n_755),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_721),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_721),
.B(n_760),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_723),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_769),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_759),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_741),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_765),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_752),
.A2(n_735),
.B(n_763),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_742),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_756),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_734),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_736),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_764),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_722),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_745),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_747),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_720),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_720),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_718),
.A2(n_727),
.B1(n_746),
.B2(n_753),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_754),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_757),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_750),
.Y(n_820)
);

INVx5_ASAP7_75t_L g821 ( 
.A(n_750),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_751),
.Y(n_822)
);

AOI21x1_ASAP7_75t_L g823 ( 
.A1(n_718),
.A2(n_761),
.B(n_750),
.Y(n_823)
);

CKINVDCx14_ASAP7_75t_R g824 ( 
.A(n_743),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_768),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_727),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_734),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_717),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_725),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_814),
.B(n_807),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_774),
.B(n_826),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_774),
.B(n_789),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_771),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_789),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_828),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_780),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_813),
.B(n_790),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_777),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_786),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_777),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_800),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_813),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_792),
.Y(n_844)
);

OA21x2_ASAP7_75t_L g845 ( 
.A1(n_806),
.A2(n_823),
.B(n_817),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_829),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_792),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_829),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_802),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_773),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_808),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_783),
.B(n_800),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_804),
.B(n_810),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_782),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_772),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_805),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_811),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_803),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_784),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_779),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_790),
.B(n_801),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_828),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_803),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_809),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_805),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_779),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_779),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_801),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_809),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_821),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_821),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_791),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_791),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_791),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_821),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_821),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_795),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_834),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_832),
.B(n_793),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_834),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_860),
.B(n_781),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_832),
.B(n_831),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_831),
.B(n_850),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_839),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_839),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_836),
.B(n_793),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_850),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_851),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_851),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_844),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_844),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_862),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_860),
.B(n_866),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_842),
.B(n_793),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_833),
.B(n_810),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_836),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_835),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_842),
.B(n_781),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_847),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_875),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_849),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_837),
.B(n_781),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_837),
.B(n_820),
.Y(n_903)
);

NOR2x1_ASAP7_75t_SL g904 ( 
.A(n_870),
.B(n_821),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_858),
.B(n_863),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_849),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_841),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_866),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_858),
.B(n_863),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_841),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_L g911 ( 
.A(n_897),
.B(n_797),
.C(n_824),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_895),
.B(n_840),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_886),
.B(n_778),
.C(n_824),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_882),
.B(n_862),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_882),
.B(n_867),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_883),
.B(n_857),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_L g917 ( 
.A(n_886),
.B(n_825),
.C(n_818),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_883),
.B(n_867),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_892),
.A2(n_818),
.B1(n_812),
.B2(n_785),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_879),
.A2(n_776),
.B1(n_819),
.B2(n_822),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_896),
.B(n_859),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_903),
.B(n_830),
.C(n_853),
.Y(n_922)
);

AOI221xp5_ASAP7_75t_L g923 ( 
.A1(n_879),
.A2(n_852),
.B1(n_855),
.B2(n_854),
.C(n_812),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_881),
.A2(n_798),
.B1(n_781),
.B2(n_820),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_903),
.B(n_845),
.C(n_798),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_894),
.A2(n_845),
.B1(n_794),
.B2(n_877),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_892),
.A2(n_795),
.B1(n_877),
.B2(n_815),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_905),
.B(n_865),
.Y(n_928)
);

OA211x2_ASAP7_75t_L g929 ( 
.A1(n_904),
.A2(n_820),
.B(n_845),
.C(n_788),
.Y(n_929)
);

AOI221xp5_ASAP7_75t_L g930 ( 
.A1(n_894),
.A2(n_787),
.B1(n_868),
.B2(n_865),
.C(n_799),
.Y(n_930)
);

NAND4xp25_ASAP7_75t_L g931 ( 
.A(n_907),
.B(n_838),
.C(n_868),
.D(n_864),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_892),
.B(n_861),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_902),
.B(n_861),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_SL g934 ( 
.A(n_898),
.B(n_787),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_905),
.B(n_838),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_915),
.B(n_893),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_921),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_912),
.B(n_910),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_928),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_916),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_917),
.B(n_909),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_935),
.B(n_893),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_918),
.B(n_893),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_933),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_914),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_932),
.B(n_904),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_922),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_934),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_931),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_926),
.B(n_893),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_930),
.Y(n_951)
);

AND2x2_ASAP7_75t_SL g952 ( 
.A(n_948),
.B(n_920),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_946),
.B(n_902),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_948),
.B(n_881),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_938),
.Y(n_955)
);

NAND3xp33_ASAP7_75t_L g956 ( 
.A(n_951),
.B(n_923),
.C(n_920),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_947),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_946),
.B(n_926),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_938),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_946),
.B(n_881),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_937),
.B(n_909),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_955),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_960),
.B(n_943),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_954),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_959),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_961),
.B(n_941),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_953),
.B(n_948),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_957),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_952),
.B(n_881),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_957),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_954),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_952),
.B(n_949),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_969),
.B(n_958),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_969),
.B(n_958),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_963),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_972),
.B(n_956),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_972),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_977),
.B(n_968),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_976),
.A2(n_967),
.B1(n_964),
.B2(n_970),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_976),
.B(n_965),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_973),
.A2(n_967),
.B1(n_964),
.B2(n_911),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_980),
.B(n_975),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_979),
.A2(n_974),
.B1(n_911),
.B2(n_913),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_978),
.Y(n_984)
);

CKINVDCx16_ASAP7_75t_R g985 ( 
.A(n_981),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_978),
.Y(n_986)
);

AOI322xp5_ASAP7_75t_L g987 ( 
.A1(n_985),
.A2(n_950),
.A3(n_962),
.B1(n_967),
.B2(n_971),
.C1(n_924),
.C2(n_945),
.Y(n_987)
);

AOI222xp33_ASAP7_75t_L g988 ( 
.A1(n_984),
.A2(n_919),
.B1(n_925),
.B2(n_927),
.C1(n_971),
.C2(n_950),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_983),
.A2(n_986),
.B(n_982),
.C(n_966),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_984),
.A2(n_940),
.B(n_796),
.C(n_939),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_985),
.B(n_775),
.C(n_796),
.Y(n_991)
);

NAND3xp33_ASAP7_75t_L g992 ( 
.A(n_984),
.B(n_827),
.C(n_900),
.Y(n_992)
);

OAI211xp5_ASAP7_75t_L g993 ( 
.A1(n_983),
.A2(n_864),
.B(n_869),
.C(n_775),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_985),
.A2(n_929),
.B1(n_900),
.B2(n_898),
.Y(n_994)
);

AOI221xp5_ASAP7_75t_L g995 ( 
.A1(n_985),
.A2(n_900),
.B1(n_910),
.B2(n_907),
.C(n_908),
.Y(n_995)
);

NOR3x1_ASAP7_75t_L g996 ( 
.A(n_993),
.B(n_876),
.C(n_871),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_L g997 ( 
.A(n_989),
.B(n_775),
.C(n_788),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_988),
.A2(n_876),
.B(n_871),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_992),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_991),
.B(n_869),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_990),
.B(n_870),
.C(n_806),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_856),
.C(n_875),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_994),
.B(n_942),
.Y(n_1003)
);

OAI211xp5_ASAP7_75t_SL g1004 ( 
.A1(n_997),
.A2(n_987),
.B(n_944),
.C(n_899),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_998),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_L g1006 ( 
.A(n_1000),
.B(n_827),
.C(n_816),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_996),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_L g1008 ( 
.A(n_1003),
.B(n_1002),
.Y(n_1008)
);

XNOR2xp5_ASAP7_75t_L g1009 ( 
.A(n_1001),
.B(n_845),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_999),
.Y(n_1011)
);

OAI211xp5_ASAP7_75t_SL g1012 ( 
.A1(n_997),
.A2(n_944),
.B(n_899),
.C(n_885),
.Y(n_1012)
);

NAND4xp25_ASAP7_75t_SL g1013 ( 
.A(n_997),
.B(n_936),
.C(n_943),
.D(n_843),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1011),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1010),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_1008),
.A2(n_900),
.B1(n_827),
.B2(n_856),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_1005),
.B(n_878),
.C(n_880),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1007),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1006),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_1004),
.B(n_878),
.C(n_880),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1012),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1009),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_1014),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1015),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1018),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_1019),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1021),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_1022),
.Y(n_1029)
);

AOI222xp33_ASAP7_75t_L g1030 ( 
.A1(n_1023),
.A2(n_827),
.B1(n_874),
.B2(n_873),
.C1(n_872),
.C2(n_936),
.Y(n_1030)
);

AND2x2_ASAP7_75t_SL g1031 ( 
.A(n_1017),
.B(n_827),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1020),
.B(n_900),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_1027),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1024),
.B(n_1016),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_1026),
.B(n_887),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_SL g1036 ( 
.A(n_1029),
.B(n_848),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1033),
.A2(n_1028),
.B1(n_1025),
.B2(n_1032),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1034),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1034),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1036),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1038),
.A2(n_1039),
.B(n_1040),
.Y(n_1041)
);

NAND5xp2_ASAP7_75t_L g1042 ( 
.A(n_1037),
.B(n_1030),
.C(n_1031),
.D(n_1035),
.E(n_843),
.Y(n_1042)
);

AOI21xp33_ASAP7_75t_SL g1043 ( 
.A1(n_1041),
.A2(n_1030),
.B(n_885),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_SL g1044 ( 
.A1(n_1042),
.A2(n_888),
.B(n_887),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1044),
.A2(n_816),
.B(n_846),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1043),
.A2(n_816),
.B1(n_908),
.B2(n_884),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_1046),
.B(n_1045),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_1046),
.A2(n_816),
.B(n_884),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_SL g1049 ( 
.A(n_1047),
.B(n_816),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1049),
.A2(n_1048),
.B1(n_889),
.B2(n_888),
.Y(n_1050)
);

OAI221xp5_ASAP7_75t_L g1051 ( 
.A1(n_1050),
.A2(n_889),
.B1(n_846),
.B2(n_848),
.C(n_890),
.Y(n_1051)
);

AOI211xp5_ASAP7_75t_L g1052 ( 
.A1(n_1051),
.A2(n_891),
.B(n_906),
.C(n_901),
.Y(n_1052)
);


endmodule