module fake_aes_7183_n_28 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
AND2x2_ASAP7_75t_L g13 ( .A(n_0), .B(n_8), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
OAI21x1_ASAP7_75t_SL g20 ( .A1(n_19), .A2(n_17), .B(n_13), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
XNOR2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_14), .Y(n_24) );
NOR2x1_ASAP7_75t_L g25 ( .A(n_24), .B(n_1), .Y(n_25) );
OA22x2_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_26) );
NOR2xp67_ASAP7_75t_L g27 ( .A(n_26), .B(n_6), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_28) );
endmodule