module fake_jpeg_29901_n_77 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_12),
.B(n_14),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_36),
.B1(n_32),
.B2(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_50),
.Y(n_56)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_20),
.Y(n_54)
);

A2O1A1O1Ixp25_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_19),
.B(n_27),
.C(n_7),
.D(n_9),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_58),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_17),
.C(n_25),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_45),
.B1(n_4),
.B2(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_11),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_16),
.B(n_22),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_67),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_66),
.C(n_55),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_55),
.B2(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_64),
.C(n_28),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_24),
.Y(n_77)
);


endmodule