module real_jpeg_6747_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_2),
.A2(n_44),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_2),
.A2(n_44),
.B1(n_281),
.B2(n_289),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_3),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_3),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_76),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_76),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_4),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_4),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_4),
.A2(n_110),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_4),
.A2(n_110),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_4),
.A2(n_110),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_5),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_5),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_197),
.B1(n_258),
.B2(n_261),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_5),
.A2(n_197),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_5),
.A2(n_197),
.B1(n_329),
.B2(n_403),
.Y(n_402)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_6),
.Y(n_129)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g425 ( 
.A(n_7),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_147),
.B1(n_151),
.B2(n_154),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_8),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_8),
.A2(n_154),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_8),
.A2(n_154),
.B1(n_208),
.B2(n_211),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_8),
.A2(n_154),
.B1(n_267),
.B2(n_366),
.Y(n_365)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_9),
.Y(n_383)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_11),
.A2(n_182),
.B1(n_183),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_11),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_11),
.B(n_252),
.C(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_11),
.B(n_136),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_11),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_11),
.B(n_83),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_11),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_12),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_12),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_12),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_12),
.Y(n_196)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_13),
.A2(n_35),
.B1(n_81),
.B2(n_164),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_14),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_14),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_14),
.A2(n_89),
.B1(n_186),
.B2(n_189),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_14),
.A2(n_89),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_14),
.A2(n_77),
.B1(n_89),
.B2(n_406),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_15),
.A2(n_46),
.B1(n_183),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_15),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_15),
.A2(n_273),
.B1(n_288),
.B2(n_293),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_15),
.A2(n_104),
.B1(n_273),
.B2(n_331),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_15),
.A2(n_116),
.B1(n_117),
.B2(n_273),
.Y(n_428)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_16),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_231),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_229),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_200),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_20),
.B(n_200),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_122),
.C(n_168),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_21),
.A2(n_22),
.B1(n_122),
.B2(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_84),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_23),
.A2(n_24),
.B(n_86),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B1(n_86),
.B2(n_121),
.Y(n_84)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_24),
.A2(n_42),
.B1(n_121),
.B2(n_417),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_25),
.A2(n_34),
.B1(n_171),
.B2(n_177),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_257),
.B(n_263),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_25),
.A2(n_241),
.B(n_263),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_25),
.A2(n_32),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_26),
.B(n_265),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_26),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_26),
.A2(n_336),
.B1(n_365),
.B2(n_368),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_26),
.A2(n_390),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_28),
.Y(n_283)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_28),
.Y(n_304)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_28),
.Y(n_369)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_29),
.Y(n_281)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_31),
.Y(n_176)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_32),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_32),
.A2(n_287),
.B(n_296),
.Y(n_286)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_41),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_42),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B1(n_75),
.B2(n_83),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_43),
.A2(n_51),
.B1(n_83),
.B2(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_46),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_46),
.B(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_47),
.Y(n_183)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_47),
.Y(n_250)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_50),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_51),
.A2(n_75),
.B1(n_83),
.B2(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_51),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_51),
.B(n_243),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_67),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_60),
.B2(n_64),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_55),
.Y(n_246)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_56),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_56),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g345 ( 
.A(n_64),
.Y(n_345)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_65),
.Y(n_244)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_67),
.A2(n_163),
.B(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_67),
.A2(n_272),
.B(n_274),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_67),
.A2(n_216),
.B1(n_272),
.B2(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_67),
.A2(n_274),
.B(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_67),
.A2(n_216),
.B1(n_405),
.B2(n_421),
.Y(n_420)
);

AOI22x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_70),
.Y(n_339)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_71),
.Y(n_254)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_83),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_108),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_96),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_88),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_90),
.B(n_241),
.Y(n_385)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_96),
.B(n_109),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_96),
.Y(n_206)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_97),
.B(n_241),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_97),
.A2(n_193),
.B1(n_194),
.B2(n_428),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_106),
.Y(n_97)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_99),
.Y(n_321)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_102),
.Y(n_226)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_108),
.A2(n_206),
.B(n_428),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_113),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_113),
.A2(n_397),
.B(n_399),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_118),
.Y(n_380)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_122),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_160),
.B(n_167),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_161),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_136),
.B1(n_145),
.B2(n_155),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_125),
.A2(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_125),
.B(n_361),
.Y(n_360)
);

AOI22x1_ASAP7_75t_L g429 ( 
.A1(n_125),
.A2(n_136),
.B1(n_361),
.B2(n_430),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_125),
.A2(n_327),
.B(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_126),
.A2(n_146),
.B1(n_185),
.B2(n_191),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_126),
.A2(n_191),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_126),
.A2(n_191),
.B1(n_359),
.B2(n_402),
.Y(n_401)
);

OR2x2_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_128),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g403 ( 
.A(n_135),
.Y(n_403)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_139),
.Y(n_346)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_147),
.B(n_382),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_201),
.CI(n_202),
.CON(n_200),
.SN(n_200)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_168),
.B(n_432),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_184),
.C(n_192),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_169),
.B(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_170),
.B(n_180),
.Y(n_440)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_171),
.Y(n_423)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_172),
.Y(n_337)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_174),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_174),
.Y(n_292)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_179),
.Y(n_341)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_181),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_184),
.B(n_192),
.Y(n_415)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_185),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_190),
.Y(n_332)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_190),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_191),
.B(n_328),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_191),
.A2(n_359),
.B(n_360),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B(n_199),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_204)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_199),
.Y(n_399)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_200),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_214),
.B2(n_228),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx8_ASAP7_75t_L g398 ( 
.A(n_210),
.Y(n_398)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_227),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_240),
.B(n_242),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_216),
.A2(n_242),
.B(n_315),
.Y(n_355)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g330 ( 
.A(n_222),
.Y(n_330)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI311xp33_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_411),
.A3(n_448),
.B1(n_466),
.C1(n_467),
.Y(n_232)
);

AOI21x1_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_372),
.B(n_410),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_350),
.B(n_371),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_309),
.B(n_349),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_277),
.B(n_308),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_255),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_238),
.B(n_255),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_247),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_239),
.A2(n_247),
.B1(n_248),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_239),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_SL g320 ( 
.A1(n_241),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g397 ( 
.A1(n_241),
.A2(n_385),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_244),
.Y(n_316)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_269),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_270),
.C(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_259),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_275),
.B2(n_276),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_299),
.B(n_307),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_285),
.B(n_298),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_297),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_297),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_335),
.B(n_340),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_305),
.Y(n_307)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_311),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_333),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_318),
.B2(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_318),
.C(n_333),
.Y(n_351)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI32xp33_ASAP7_75t_L g342 ( 
.A1(n_323),
.A2(n_343),
.A3(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_342)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_342),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_342),
.Y(n_356)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_351),
.B(n_352),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_357),
.B2(n_370),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_356),
.C(n_370),
.Y(n_373)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_363),
.C(n_364),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_373),
.B(n_374),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_394),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_375)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_376),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_386),
.B2(n_387),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_378),
.B(n_386),
.Y(n_444)
);

OAI32xp33_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_380),
.A3(n_381),
.B1(n_384),
.B2(n_385),
.Y(n_378)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_393),
.C(n_394),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_400),
.B2(n_409),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_395),
.B(n_401),
.C(n_404),
.Y(n_457)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_434),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_SL g467 ( 
.A1(n_412),
.A2(n_434),
.B(n_468),
.C(n_471),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_431),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_431),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.C(n_418),
.Y(n_413)
);

FAx1_ASAP7_75t_SL g447 ( 
.A(n_414),
.B(n_416),
.CI(n_418),
.CON(n_447),
.SN(n_447)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_426),
.C(n_429),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_422),
.Y(n_456)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_426),
.A2(n_427),
.B1(n_429),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_429),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_447),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_447),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_440),
.C(n_441),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_436),
.A2(n_437),
.B1(n_440),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.C(n_445),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_442),
.A2(n_443),
.B1(n_445),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_444),
.B(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_445),
.Y(n_454)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_447),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_461),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_469),
.B(n_470),
.Y(n_468)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_458),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_458),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.C(n_457),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_464),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_455),
.A2(n_456),
.B1(n_457),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_457),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_463),
.Y(n_469)
);


endmodule