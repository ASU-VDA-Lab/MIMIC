module fake_jpeg_3285_n_395 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_53),
.Y(n_143)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_54),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_59),
.Y(n_150)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_7),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_63),
.A2(n_72),
.B(n_75),
.Y(n_165)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_76),
.Y(n_113)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_65),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_69),
.B(n_95),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_52),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_34),
.B(n_8),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_84),
.Y(n_115)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_14),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_82),
.B(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_15),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_88),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_11),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_93),
.Y(n_116)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_89),
.B(n_99),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_13),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_91),
.B(n_100),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_96),
.B(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_30),
.A2(n_13),
.B1(n_9),
.B2(n_3),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_98),
.A2(n_18),
.B1(n_75),
.B2(n_19),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_9),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_101),
.B(n_106),
.Y(n_166)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_105),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_46),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_27),
.B(n_1),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_108),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_1),
.B(n_2),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_97),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_50),
.B(n_47),
.C(n_44),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_110),
.A2(n_166),
.B(n_163),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_32),
.B1(n_45),
.B2(n_46),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_114),
.A2(n_138),
.B1(n_151),
.B2(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_119),
.B(n_131),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_80),
.A2(n_35),
.B1(n_24),
.B2(n_37),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_123),
.A2(n_129),
.B1(n_136),
.B2(n_152),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_30),
.B1(n_21),
.B2(n_33),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_29),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_132),
.B(n_133),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_43),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_66),
.A2(n_37),
.B1(n_36),
.B2(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_36),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_55),
.A2(n_50),
.B1(n_47),
.B2(n_28),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_30),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_142),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_75),
.B(n_33),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_141),
.B(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_44),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_42),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_149),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_56),
.A2(n_33),
.B1(n_21),
.B2(n_45),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_148),
.A2(n_114),
.B1(n_153),
.B2(n_174),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_57),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_67),
.A2(n_42),
.B1(n_28),
.B2(n_45),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_77),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_77),
.A2(n_46),
.B1(n_5),
.B2(n_6),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_167),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_53),
.A2(n_1),
.B1(n_6),
.B2(n_26),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_70),
.A2(n_71),
.B1(n_83),
.B2(n_90),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_105),
.A2(n_26),
.B1(n_106),
.B2(n_98),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_58),
.A2(n_35),
.B1(n_39),
.B2(n_80),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_173),
.B1(n_133),
.B2(n_132),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_63),
.B(n_106),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_69),
.B(n_63),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_143),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_113),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_182),
.B(n_202),
.Y(n_260)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_134),
.A2(n_154),
.B(n_178),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_188),
.A2(n_235),
.B(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_118),
.B1(n_129),
.B2(n_150),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_195),
.A2(n_210),
.B1(n_215),
.B2(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_211),
.Y(n_241)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_200),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_201),
.B(n_231),
.C(n_233),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_120),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_141),
.B1(n_128),
.B2(n_119),
.Y(n_205)
);

AO22x1_ASAP7_75t_L g252 ( 
.A1(n_205),
.A2(n_221),
.B1(n_220),
.B2(n_187),
.Y(n_252)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_207),
.Y(n_255)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_208),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_222),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_118),
.B(n_117),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_217),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_118),
.A2(n_150),
.B1(n_125),
.B2(n_121),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_184),
.B1(n_189),
.B2(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_165),
.A2(n_131),
.B1(n_174),
.B2(n_153),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_219),
.B1(n_226),
.B2(n_193),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_139),
.B1(n_155),
.B2(n_124),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_116),
.B(n_122),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_224),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_124),
.A2(n_155),
.B1(n_139),
.B2(n_164),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_234),
.Y(n_268)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_144),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_110),
.A2(n_111),
.B1(n_164),
.B2(n_121),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_145),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_229),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_125),
.A2(n_111),
.B1(n_115),
.B2(n_122),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_157),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_143),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_143),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_143),
.A2(n_134),
.B(n_154),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_240),
.A2(n_259),
.B1(n_238),
.B2(n_246),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_182),
.B(n_190),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_248),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_212),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_197),
.B(n_199),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_249),
.B(n_257),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_180),
.A2(n_194),
.B1(n_221),
.B2(n_214),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_SL g307 ( 
.A1(n_250),
.A2(n_276),
.B(n_242),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_205),
.B(n_203),
.CI(n_188),
.CON(n_251),
.SN(n_251)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_251),
.B(n_266),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_252),
.A2(n_253),
.B1(n_266),
.B2(n_240),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_186),
.A2(n_235),
.B1(n_192),
.B2(n_211),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_197),
.B(n_199),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_SL g258 ( 
.A(n_220),
.B(n_211),
.C(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_262),
.C(n_268),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_191),
.B(n_225),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_271),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_223),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_196),
.B(n_222),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_263),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_229),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_185),
.A2(n_217),
.B(n_200),
.C(n_204),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_252),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_241),
.A2(n_208),
.B1(n_183),
.B2(n_179),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_279),
.A2(n_287),
.B1(n_236),
.B2(n_237),
.Y(n_319)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_239),
.A2(n_233),
.B(n_206),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_307),
.B(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_285),
.B(n_298),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_303),
.C(n_255),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_241),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_297),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_264),
.B1(n_274),
.B2(n_275),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_295),
.A2(n_296),
.B(n_242),
.Y(n_313)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_244),
.B(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_304),
.Y(n_315)
);

AOI22x1_ASAP7_75t_SL g302 ( 
.A1(n_251),
.A2(n_258),
.B1(n_267),
.B2(n_277),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_262),
.B(n_244),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_272),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_309),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_276),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_306),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_238),
.A2(n_245),
.B(n_243),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_270),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_317),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_290),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_287),
.A2(n_264),
.B1(n_242),
.B2(n_255),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_316),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_285),
.C(n_303),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_236),
.B1(n_237),
.B2(n_275),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_318),
.A2(n_319),
.B1(n_327),
.B2(n_311),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_305),
.A2(n_273),
.B1(n_298),
.B2(n_291),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_273),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_321),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_334),
.Y(n_351)
);

OA22x2_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_299),
.B1(n_292),
.B2(n_280),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_342),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_313),
.A2(n_299),
.B(n_282),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_317),
.B(n_312),
.Y(n_332)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_338),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_333),
.Y(n_358)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_301),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_337),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_321),
.A2(n_302),
.B(n_281),
.C(n_308),
.Y(n_337)
);

AOI221xp5_ASAP7_75t_L g339 ( 
.A1(n_327),
.A2(n_300),
.B1(n_279),
.B2(n_283),
.C(n_288),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_344),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_289),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_341),
.Y(n_356)
);

OAI321xp33_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_278),
.A3(n_284),
.B1(n_297),
.B2(n_309),
.C(n_326),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_319),
.B1(n_322),
.B2(n_326),
.Y(n_343)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_320),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_315),
.A2(n_324),
.B(n_325),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_346),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_359),
.C(n_360),
.Y(n_369)
);

XOR2x1_ASAP7_75t_SL g355 ( 
.A(n_345),
.B(n_330),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_329),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_310),
.C(n_325),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_324),
.C(n_311),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_354),
.A2(n_356),
.B(n_353),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_361),
.A2(n_364),
.B(n_331),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_356),
.A2(n_342),
.B1(n_349),
.B2(n_351),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_358),
.B1(n_357),
.B2(n_343),
.Y(n_378)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_365),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_352),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_350),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_366),
.B(n_368),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_344),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_336),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_358),
.B1(n_335),
.B2(n_346),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_376),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_359),
.C(n_348),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_369),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_378),
.B(n_361),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_380),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_375),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_373),
.B(n_367),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_381),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_389)
);

AOI31xp33_ASAP7_75t_SL g382 ( 
.A1(n_376),
.A2(n_337),
.A3(n_341),
.B(n_330),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_362),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_377),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_386),
.B(n_387),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_384),
.A2(n_354),
.B(n_370),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_323),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_392),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_390),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_389),
.Y(n_395)
);


endmodule