module fake_netlist_6_3255_n_808 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_808);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_808;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_47),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_13),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_127),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_36),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_68),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_12),
.B(n_55),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_8),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_117),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_4),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_34),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_94),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_119),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_27),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_114),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_16),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_77),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_74),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_18),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_168),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_87),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_9),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_135),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_37),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_95),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_26),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_137),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_99),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_13),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_51),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_20),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_5),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_62),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_54),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_33),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_104),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_5),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_130),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_61),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_98),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_128),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_32),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_0),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_183),
.B(n_0),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_1),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_227),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_21),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_22),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_204),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_R g258 ( 
.A1(n_172),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_23),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_2),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_192),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_223),
.B(n_24),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_196),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_205),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_6),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_230),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_224),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_184),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_248),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_173),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_178),
.C(n_175),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_234),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g306 ( 
.A1(n_242),
.A2(n_181),
.B(n_179),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_260),
.B(n_230),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_269),
.B(n_185),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_248),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_246),
.B(n_188),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_200),
.C(n_226),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_189),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_245),
.A2(n_191),
.B(n_222),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_251),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_243),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_269),
.B(n_193),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_262),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_244),
.B(n_195),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_249),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g327 ( 
.A1(n_236),
.A2(n_206),
.B1(n_213),
.B2(n_210),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_289),
.B(n_251),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_272),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_254),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_326),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

OR2x6_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_279),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_L g340 ( 
.A(n_288),
.B(n_278),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_254),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_311),
.B(n_254),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_311),
.B(n_256),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_267),
.Y(n_346)
);

BUFx6f_ASAP7_75t_SL g347 ( 
.A(n_288),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

AND3x1_ASAP7_75t_L g349 ( 
.A(n_281),
.B(n_273),
.C(n_258),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_280),
.B(n_256),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_307),
.B(n_313),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_256),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_298),
.B(n_270),
.Y(n_356)
);

NOR3xp33_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_257),
.C(n_271),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_267),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_322),
.B(n_255),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_270),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_270),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_306),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_259),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_327),
.B(n_264),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_316),
.B(n_198),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_306),
.B(n_275),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_299),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_320),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_306),
.B(n_250),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_288),
.B(n_328),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_283),
.B(n_250),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_288),
.A2(n_258),
.B1(n_186),
.B2(n_229),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_293),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_288),
.B(n_250),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_285),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_293),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_297),
.B(n_250),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_316),
.B(n_199),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_294),
.B(n_263),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_L g385 ( 
.A(n_308),
.B(n_202),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_318),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_294),
.B(n_263),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_301),
.B(n_263),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_301),
.B(n_265),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_320),
.B(n_208),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_318),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_321),
.B(n_265),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_308),
.B(n_265),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_321),
.B(n_265),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_317),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_362),
.A2(n_309),
.B1(n_323),
.B2(n_302),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_336),
.B(n_329),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_374),
.A2(n_300),
.B(n_329),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_346),
.B(n_317),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_362),
.A2(n_286),
.B(n_284),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_342),
.A2(n_300),
.B(n_287),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_303),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_368),
.A2(n_315),
.B(n_291),
.C(n_290),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_360),
.A2(n_300),
.B(n_287),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_364),
.A2(n_372),
.B(n_365),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_350),
.B(n_284),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_291),
.B(n_290),
.C(n_286),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_25),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_343),
.B(n_344),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_265),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_356),
.A2(n_379),
.B(n_340),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_358),
.B(n_359),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_266),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_348),
.A2(n_300),
.B(n_287),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_358),
.B(n_266),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_351),
.A2(n_277),
.B(n_266),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_345),
.A2(n_277),
.B1(n_266),
.B2(n_229),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_384),
.A2(n_277),
.B(n_266),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_357),
.B(n_277),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_387),
.A2(n_277),
.B(n_91),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_388),
.A2(n_90),
.B(n_171),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_366),
.B(n_186),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_389),
.A2(n_84),
.B(n_165),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_380),
.B(n_169),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_347),
.A2(n_83),
.B1(n_161),
.B2(n_159),
.Y(n_432)
);

O2A1O1Ixp33_ASAP7_75t_SL g433 ( 
.A1(n_365),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_357),
.B(n_378),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_393),
.A2(n_82),
.B(n_158),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_28),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_354),
.B(n_29),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_369),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_367),
.A2(n_86),
.B(n_156),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_395),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_331),
.B(n_7),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_367),
.A2(n_383),
.B(n_371),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_377),
.B(n_10),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_339),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_373),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_376),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_375),
.B(n_30),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_347),
.A2(n_92),
.B1(n_155),
.B2(n_152),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_339),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_332),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_341),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_333),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_383),
.A2(n_80),
.B(n_151),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_375),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_455)
);

NOR2x1_ASAP7_75t_L g456 ( 
.A(n_330),
.B(n_31),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_385),
.A2(n_392),
.B(n_394),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_339),
.B(n_14),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_390),
.B(n_15),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_377),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_390),
.A2(n_97),
.B(n_150),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_382),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_334),
.B(n_19),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_35),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_406),
.A2(n_349),
.B(n_352),
.Y(n_465)
);

AO31x2_ASAP7_75t_L g466 ( 
.A1(n_415),
.A2(n_409),
.A3(n_422),
.B(n_459),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_417),
.B(n_406),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_411),
.A2(n_352),
.B1(n_341),
.B2(n_40),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

AO31x2_ASAP7_75t_L g471 ( 
.A1(n_455),
.A2(n_352),
.A3(n_341),
.B(n_41),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_396),
.B(n_341),
.Y(n_472)
);

AO21x2_ASAP7_75t_L g473 ( 
.A1(n_442),
.A2(n_352),
.B(n_39),
.Y(n_473)
);

AO31x2_ASAP7_75t_L g474 ( 
.A1(n_462),
.A2(n_38),
.A3(n_42),
.B(n_44),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_429),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_45),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_407),
.B(n_46),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_414),
.A2(n_48),
.B(n_49),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_399),
.A2(n_164),
.B(n_52),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_403),
.A2(n_50),
.B1(n_53),
.B2(n_56),
.Y(n_481)
);

AO31x2_ASAP7_75t_L g482 ( 
.A1(n_398),
.A2(n_57),
.A3(n_58),
.B(n_59),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_452),
.A2(n_60),
.B(n_63),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_442),
.A2(n_64),
.B(n_65),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_434),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_412),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_418),
.B(n_70),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_452),
.A2(n_71),
.B(n_72),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_452),
.A2(n_75),
.B(n_76),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_78),
.Y(n_490)
);

AOI21x1_ASAP7_75t_SL g491 ( 
.A1(n_436),
.A2(n_79),
.B(n_93),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_450),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_449),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_397),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

NAND3xp33_ASAP7_75t_L g497 ( 
.A(n_443),
.B(n_107),
.C(n_108),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_452),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_457),
.A2(n_401),
.B(n_402),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_110),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_413),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_401),
.A2(n_111),
.B(n_112),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_405),
.A2(n_113),
.B(n_115),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_424),
.A2(n_116),
.B(n_118),
.C(n_120),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_446),
.B(n_121),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_451),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_408),
.A2(n_122),
.B(n_123),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_458),
.B(n_456),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_410),
.B(n_124),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_404),
.A2(n_125),
.B(n_126),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_453),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_439),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_419),
.A2(n_134),
.B(n_136),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_437),
.A2(n_149),
.B(n_139),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_447),
.A2(n_138),
.B(n_142),
.Y(n_516)
);

AOI21xp33_ASAP7_75t_L g517 ( 
.A1(n_460),
.A2(n_143),
.B(n_145),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_464),
.A2(n_146),
.B(n_147),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_432),
.B(n_148),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_470),
.B(n_445),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_433),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_480),
.A2(n_454),
.B1(n_439),
.B2(n_448),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_499),
.A2(n_454),
.B(n_421),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_467),
.B(n_463),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_467),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_479),
.A2(n_425),
.B(n_461),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_491),
.A2(n_427),
.B(n_430),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_492),
.B(n_423),
.Y(n_530)
);

BUFx2_ASAP7_75t_R g531 ( 
.A(n_475),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_515),
.A2(n_435),
.B(n_500),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_487),
.A2(n_507),
.B(n_503),
.Y(n_534)
);

NAND2x1p5_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_498),
.Y(n_535)
);

OAI21xp33_ASAP7_75t_L g536 ( 
.A1(n_476),
.A2(n_465),
.B(n_508),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_498),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_494),
.B(n_496),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_506),
.B(n_512),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_502),
.A2(n_484),
.B(n_511),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_501),
.B(n_509),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

CKINVDCx14_ASAP7_75t_R g544 ( 
.A(n_490),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_472),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_466),
.B(n_471),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_472),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_518),
.B(n_510),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_505),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_513),
.A2(n_510),
.B(n_473),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_520),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_514),
.A2(n_516),
.B(n_519),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_471),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_478),
.A2(n_488),
.B(n_483),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_466),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_497),
.C(n_495),
.Y(n_556)
);

OA21x2_ASAP7_75t_L g557 ( 
.A1(n_504),
.A2(n_469),
.B(n_489),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_471),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_474),
.B(n_482),
.Y(n_560)
);

CKINVDCx11_ASAP7_75t_R g561 ( 
.A(n_485),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_493),
.A2(n_481),
.B(n_474),
.Y(n_562)
);

OAI21x1_ASAP7_75t_SL g563 ( 
.A1(n_520),
.A2(n_502),
.B(n_484),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_520),
.B(n_482),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_482),
.A2(n_499),
.B(n_479),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_563),
.A2(n_520),
.B1(n_544),
.B2(n_551),
.Y(n_566)
);

AO21x2_ASAP7_75t_L g567 ( 
.A1(n_540),
.A2(n_565),
.B(n_560),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_543),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_543),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_555),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_555),
.Y(n_571)
);

INVx4_ASAP7_75t_SL g572 ( 
.A(n_551),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_545),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_526),
.Y(n_576)
);

AO21x1_ASAP7_75t_SL g577 ( 
.A1(n_553),
.A2(n_549),
.B(n_536),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_531),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_541),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_544),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_530),
.B(n_522),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_561),
.A2(n_556),
.B1(n_551),
.B2(n_523),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_537),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_521),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_521),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_542),
.B(n_547),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_521),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_539),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_565),
.A2(n_527),
.B(n_554),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_527),
.A2(n_554),
.B(n_552),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_546),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_546),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_559),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_552),
.A2(n_534),
.B(n_529),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_534),
.A2(n_529),
.B(n_533),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_559),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_548),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_524),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_522),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_558),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_535),
.Y(n_604)
);

AO21x2_ASAP7_75t_L g605 ( 
.A1(n_540),
.A2(n_550),
.B(n_562),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_603),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_582),
.B(n_551),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_568),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_568),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_584),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_564),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_569),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_583),
.A2(n_561),
.B1(n_564),
.B2(n_542),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_582),
.A2(n_564),
.B1(n_525),
.B2(n_557),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_535),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_595),
.B(n_562),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_566),
.A2(n_557),
.B1(n_537),
.B2(n_524),
.Y(n_617)
);

NOR2x1_ASAP7_75t_SL g618 ( 
.A(n_577),
.B(n_532),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_595),
.B(n_557),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_569),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_600),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_602),
.B(n_590),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_603),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_579),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_581),
.B(n_537),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_586),
.B(n_532),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_586),
.B(n_532),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_588),
.B(n_532),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_570),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_588),
.B(n_533),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_572),
.B(n_590),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_574),
.B(n_575),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_574),
.B(n_575),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_579),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_571),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_587),
.B(n_576),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_596),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_572),
.B(n_604),
.Y(n_640)
);

AOI222xp33_ASAP7_75t_L g641 ( 
.A1(n_587),
.A2(n_591),
.B1(n_578),
.B2(n_580),
.C1(n_573),
.C2(n_589),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_576),
.B(n_585),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_580),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_584),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_585),
.B(n_573),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_589),
.B(n_604),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_599),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_572),
.B(n_577),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_567),
.B(n_599),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_601),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_572),
.B(n_589),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_584),
.B(n_567),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_601),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_567),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_631),
.B(n_605),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_621),
.B(n_622),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_650),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_622),
.B(n_605),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_637),
.B(n_605),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_637),
.B(n_597),
.Y(n_661)
);

AOI222xp33_ASAP7_75t_L g662 ( 
.A1(n_613),
.A2(n_592),
.B1(n_593),
.B2(n_597),
.C1(n_598),
.C2(n_625),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_607),
.B(n_598),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_606),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_641),
.A2(n_592),
.B1(n_593),
.B2(n_607),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_650),
.B(n_653),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_608),
.Y(n_667)
);

AOI222xp33_ASAP7_75t_L g668 ( 
.A1(n_635),
.A2(n_645),
.B1(n_623),
.B2(n_606),
.C1(n_626),
.C2(n_614),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_645),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_623),
.A2(n_615),
.B1(n_646),
.B2(n_627),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_619),
.B(n_616),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_619),
.B(n_616),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_617),
.B(n_615),
.C(n_642),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_642),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_653),
.B(n_611),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_611),
.B(n_612),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_612),
.B(n_630),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_633),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_634),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_609),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_609),
.B(n_639),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_639),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_620),
.B(n_638),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_620),
.B(n_636),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_624),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_627),
.B(n_629),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_624),
.B(n_638),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_636),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_628),
.B(n_629),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_647),
.B(n_628),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_647),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_680),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_683),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_682),
.B(n_649),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_657),
.B(n_648),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_671),
.B(n_655),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_669),
.B(n_648),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_671),
.B(n_655),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_666),
.B(n_654),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_682),
.B(n_649),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_672),
.B(n_654),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_680),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_685),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_669),
.B(n_651),
.Y(n_704)
);

NAND2x1p5_ASAP7_75t_L g705 ( 
.A(n_664),
.B(n_644),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_683),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_664),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_686),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_679),
.B(n_651),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_689),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_685),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_688),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_672),
.B(n_618),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_679),
.B(n_610),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_688),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_674),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_691),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_SL g718 ( 
.A1(n_668),
.A2(n_652),
.B(n_640),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_693),
.B(n_656),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_706),
.B(n_656),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_692),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_696),
.B(n_656),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_712),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_712),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_694),
.B(n_663),
.Y(n_725)
);

OAI21xp33_ASAP7_75t_L g726 ( 
.A1(n_718),
.A2(n_670),
.B(n_665),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_696),
.B(n_656),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_715),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_710),
.B(n_676),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_716),
.B(n_666),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_692),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_714),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_721),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_730),
.B(n_675),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_732),
.A2(n_673),
.B1(n_708),
.B2(n_675),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_725),
.B(n_727),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_721),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_731),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_731),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_SL g740 ( 
.A(n_726),
.B(n_643),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_723),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_724),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_735),
.B(n_729),
.Y(n_743)
);

AOI221xp5_ASAP7_75t_L g744 ( 
.A1(n_740),
.A2(n_728),
.B1(n_719),
.B2(n_720),
.C(n_695),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_741),
.Y(n_745)
);

AOI221xp5_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_720),
.B1(n_719),
.B2(n_727),
.C(n_722),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_734),
.A2(n_673),
.B1(n_694),
.B2(n_700),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_733),
.A2(n_618),
.B(n_662),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_736),
.A2(n_694),
.B1(n_700),
.B2(n_705),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_733),
.Y(n_750)
);

OAI311xp33_ASAP7_75t_L g751 ( 
.A1(n_744),
.A2(n_662),
.A3(n_699),
.B1(n_697),
.C1(n_709),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_SL g752 ( 
.A(n_743),
.B(n_643),
.C(n_704),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_L g753 ( 
.A1(n_747),
.A2(n_739),
.B1(n_738),
.B2(n_737),
.C(n_705),
.Y(n_753)
);

OAI211xp5_ASAP7_75t_L g754 ( 
.A1(n_748),
.A2(n_746),
.B(n_745),
.C(n_750),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_749),
.B(n_722),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_700),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_754),
.B(n_713),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_755),
.B(n_713),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

NAND4xp75_ASAP7_75t_L g760 ( 
.A(n_757),
.B(n_751),
.C(n_707),
.D(n_652),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_759),
.B(n_701),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_761),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_760),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_761),
.Y(n_764)
);

NOR2x1_ASAP7_75t_L g765 ( 
.A(n_763),
.B(n_756),
.Y(n_765)
);

NAND4xp75_ASAP7_75t_L g766 ( 
.A(n_762),
.B(n_758),
.C(n_707),
.D(n_690),
.Y(n_766)
);

NOR2x1_ASAP7_75t_L g767 ( 
.A(n_763),
.B(n_715),
.Y(n_767)
);

INVxp33_ASAP7_75t_SL g768 ( 
.A(n_764),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_763),
.A2(n_690),
.B1(n_701),
.B2(n_683),
.Y(n_769)
);

NAND4xp75_ASAP7_75t_L g770 ( 
.A(n_762),
.B(n_698),
.C(n_687),
.D(n_684),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_768),
.B(n_765),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_767),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_769),
.Y(n_773)
);

XNOR2x1_ASAP7_75t_L g774 ( 
.A(n_766),
.B(n_705),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_770),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_770),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_768),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_771),
.A2(n_699),
.B1(n_660),
.B2(n_702),
.Y(n_778)
);

OAI21xp33_ASAP7_75t_L g779 ( 
.A1(n_777),
.A2(n_698),
.B(n_663),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_773),
.A2(n_640),
.B1(n_683),
.B2(n_632),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_772),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_775),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_776),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_782),
.A2(n_776),
.B1(n_774),
.B2(n_640),
.Y(n_784)
);

AOI211xp5_ASAP7_75t_L g785 ( 
.A1(n_781),
.A2(n_640),
.B(n_632),
.C(n_610),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_783),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_780),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_778),
.A2(n_717),
.B(n_711),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_779),
.B(n_717),
.Y(n_789)
);

AOI211xp5_ASAP7_75t_L g790 ( 
.A1(n_782),
.A2(n_632),
.B(n_610),
.C(n_659),
.Y(n_790)
);

OA22x2_ASAP7_75t_L g791 ( 
.A1(n_781),
.A2(n_632),
.B1(n_711),
.B2(n_703),
.Y(n_791)
);

OAI221xp5_ASAP7_75t_L g792 ( 
.A1(n_786),
.A2(n_644),
.B1(n_703),
.B2(n_702),
.C(n_661),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_788),
.Y(n_793)
);

OA22x2_ASAP7_75t_L g794 ( 
.A1(n_784),
.A2(n_691),
.B1(n_678),
.B2(n_667),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_787),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_791),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_785),
.B(n_687),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_789),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_SL g799 ( 
.A1(n_795),
.A2(n_790),
.B1(n_644),
.B2(n_610),
.Y(n_799)
);

AO21x2_ASAP7_75t_L g800 ( 
.A1(n_793),
.A2(n_681),
.B(n_684),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_796),
.A2(n_658),
.B1(n_678),
.B2(n_667),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_798),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_802),
.B(n_797),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_799),
.B(n_794),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_801),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_803),
.A2(n_792),
.B(n_800),
.Y(n_806)
);

XNOR2xp5_ASAP7_75t_L g807 ( 
.A(n_806),
.B(n_805),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_807),
.A2(n_804),
.B(n_677),
.Y(n_808)
);


endmodule