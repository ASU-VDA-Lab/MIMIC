module fake_jpeg_19514_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_47),
.Y(n_72)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_55),
.Y(n_65)
);

OR2x4_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_72),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_44),
.B1(n_53),
.B2(n_51),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_74),
.B1(n_52),
.B2(n_53),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_76),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_3),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_48),
.B1(n_42),
.B2(n_54),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_49),
.B1(n_45),
.B2(n_41),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_23),
.B1(n_37),
.B2(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_86),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_75),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_3),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_89),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_20),
.B1(n_34),
.B2(n_32),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_88),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_66),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_84),
.C(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_93),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_74),
.B(n_88),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_4),
.B(n_5),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_103),
.A3(n_97),
.B1(n_98),
.B2(n_94),
.C1(n_6),
.C2(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_5),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_97),
.B1(n_7),
.B2(n_6),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_102),
.B(n_101),
.C(n_16),
.D(n_17),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_106),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_108),
.A2(n_107),
.B(n_106),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_109),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_9),
.Y(n_112)
);

AOI31xp67_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_12),
.A3(n_18),
.B(n_21),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_24),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_38),
.B1(n_29),
.B2(n_30),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_117),
.Y(n_118)
);


endmodule