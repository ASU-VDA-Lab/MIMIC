module fake_aes_11674_n_655 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_655);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_655;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_285;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_51), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_67), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_87), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_80), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_70), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_65), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_35), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_63), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_49), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_62), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_56), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_78), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_10), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_12), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_76), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_59), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_3), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_43), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_13), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_64), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_86), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_34), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_11), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_46), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_61), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_6), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_26), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_2), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_77), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_57), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_12), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_74), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_25), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_18), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_33), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_53), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_4), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_118), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_118), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_118), .B(n_0), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_99), .B(n_1), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_118), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_101), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
XOR2xp5_ASAP7_75t_L g137 ( .A(n_105), .B(n_1), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
BUFx8_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_101), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_111), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_88), .B(n_2), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_107), .B(n_4), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_111), .B(n_5), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
BUFx2_ASAP7_75t_L g156 ( .A(n_107), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_135), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_131), .B(n_120), .Y(n_159) );
INVx1_ASAP7_75t_SL g160 ( .A(n_154), .Y(n_160) );
AND2x6_ASAP7_75t_L g161 ( .A(n_131), .B(n_95), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_131), .B(n_95), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_156), .B(n_120), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_156), .B(n_109), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_153), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
OAI221xp5_ASAP7_75t_L g174 ( .A1(n_132), .A2(n_113), .B1(n_88), .B2(n_115), .C(n_125), .Y(n_174) );
AO22x2_ASAP7_75t_L g175 ( .A1(n_153), .A2(n_97), .B1(n_127), .B2(n_126), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_138), .B(n_102), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_138), .B(n_117), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_149), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_153), .A2(n_113), .B1(n_115), .B2(n_116), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
AND2x6_ASAP7_75t_L g183 ( .A(n_153), .B(n_97), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_149), .A2(n_116), .B1(n_125), .B2(n_121), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_136), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_132), .A2(n_121), .B1(n_122), .B2(n_124), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_139), .B(n_93), .Y(n_188) );
AO22x2_ASAP7_75t_L g189 ( .A1(n_154), .A2(n_114), .B1(n_127), .B2(n_126), .Y(n_189) );
AND2x6_ASAP7_75t_L g190 ( .A(n_183), .B(n_98), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_189), .A2(n_139), .B1(n_142), .B2(n_151), .Y(n_191) );
NAND3xp33_ASAP7_75t_SL g192 ( .A(n_160), .B(n_134), .C(n_144), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_170), .B(n_139), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_172), .B(n_158), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_168), .B(n_139), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_181), .B(n_150), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_176), .B(n_142), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_162), .A2(n_155), .B(n_151), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_189), .A2(n_155), .B1(n_143), .B2(n_146), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_186), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_158), .B(n_152), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_177), .B(n_143), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_159), .B(n_146), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_159), .A2(n_148), .B1(n_106), .B2(n_150), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_183), .B(n_122), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_183), .B(n_152), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_158), .B(n_100), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_159), .B(n_152), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_158), .B(n_96), .Y(n_214) );
OR2x2_ASAP7_75t_SL g215 ( .A(n_189), .B(n_137), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_189), .A2(n_128), .B1(n_103), .B2(n_104), .Y(n_217) );
INVxp67_ASAP7_75t_L g218 ( .A(n_174), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_186), .B(n_112), .Y(n_219) );
OAI21xp33_ASAP7_75t_SL g220 ( .A1(n_164), .A2(n_98), .B(n_103), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_167), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_167), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_169), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_172), .A2(n_128), .B1(n_104), .B2(n_108), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_169), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_187), .B(n_137), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_173), .Y(n_228) );
NOR2xp67_ASAP7_75t_L g229 ( .A(n_188), .B(n_5), .Y(n_229) );
NOR2x2_ASAP7_75t_L g230 ( .A(n_175), .B(n_7), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_172), .B(n_108), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_173), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_184), .B(n_7), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_195), .A2(n_180), .B(n_186), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_198), .A2(n_175), .B1(n_183), .B2(n_165), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_201), .B(n_180), .Y(n_236) );
BUFx12f_ASAP7_75t_L g237 ( .A(n_215), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_198), .A2(n_175), .B1(n_183), .B2(n_165), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_197), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_205), .B(n_183), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_226), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_196), .B(n_161), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_226), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_198), .B(n_183), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_215), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_199), .B(n_204), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_194), .B(n_161), .Y(n_249) );
BUFx12f_ASAP7_75t_L g250 ( .A(n_233), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_218), .A2(n_182), .B(n_178), .C(n_114), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_217), .A2(n_175), .B1(n_182), .B2(n_178), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_213), .B(n_161), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_228), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
INVx5_ASAP7_75t_L g256 ( .A(n_190), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_197), .Y(n_257) );
AND2x6_ASAP7_75t_L g258 ( .A(n_209), .B(n_161), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_190), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_191), .B(n_161), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_232), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_193), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_209), .A2(n_165), .B1(n_161), .B2(n_110), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_195), .B(n_161), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_200), .B(n_165), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_212), .B(n_165), .Y(n_267) );
INVx6_ASAP7_75t_L g268 ( .A(n_202), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_190), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_210), .A2(n_165), .B1(n_119), .B2(n_123), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_208), .Y(n_271) );
INVx4_ASAP7_75t_L g272 ( .A(n_190), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_207), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_233), .A2(n_165), .B1(n_179), .B2(n_171), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_216), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_190), .B(n_8), .Y(n_276) );
INVx3_ASAP7_75t_SL g277 ( .A(n_258), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_248), .A2(n_220), .B(n_225), .C(n_231), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_247), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_241), .Y(n_280) );
AND2x6_ASAP7_75t_L g281 ( .A(n_238), .B(n_210), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_241), .A2(n_231), .B(n_211), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_246), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_255), .B(n_221), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_243), .A2(n_203), .B(n_229), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_272), .B(n_256), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_243), .B(n_203), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_244), .A2(n_203), .B(n_223), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_255), .B(n_222), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_244), .A2(n_214), .B(n_216), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_259), .Y(n_291) );
BUFx8_ASAP7_75t_L g292 ( .A(n_258), .Y(n_292) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_236), .A2(n_136), .B(n_140), .Y(n_293) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_254), .A2(n_140), .B(n_141), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_254), .A2(n_190), .B(n_219), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_252), .A2(n_140), .B(n_141), .Y(n_296) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_261), .A2(n_141), .B(n_145), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_245), .A2(n_145), .B(n_147), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_237), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_261), .Y(n_300) );
CKINVDCx11_ASAP7_75t_R g301 ( .A(n_237), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_250), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_234), .A2(n_145), .B(n_147), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_238), .A2(n_206), .B1(n_230), .B2(n_202), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_250), .A2(n_227), .B1(n_192), .B2(n_230), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_251), .A2(n_147), .B(n_179), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_267), .A2(n_166), .B(n_179), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_235), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_262), .B(n_227), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_249), .A2(n_171), .B(n_166), .C(n_185), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_310), .A2(n_262), .B1(n_271), .B2(n_260), .C(n_274), .Y(n_312) );
BUFx12f_ASAP7_75t_L g313 ( .A(n_292), .Y(n_313) );
AOI22xp33_ASAP7_75t_SL g314 ( .A1(n_305), .A2(n_260), .B1(n_258), .B2(n_242), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_300), .B(n_271), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_309), .A2(n_270), .B1(n_264), .B2(n_273), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_303), .Y(n_317) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_306), .A2(n_270), .B1(n_240), .B2(n_253), .C(n_276), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_305), .A2(n_265), .B1(n_266), .B2(n_258), .Y(n_319) );
INVx4_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_310), .A2(n_265), .B1(n_266), .B2(n_275), .C(n_239), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g322 ( .A1(n_309), .A2(n_265), .B1(n_258), .B2(n_272), .C1(n_263), .C2(n_275), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_280), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g324 ( .A1(n_290), .A2(n_275), .B(n_273), .Y(n_324) );
AO31x2_ASAP7_75t_L g325 ( .A1(n_290), .A2(n_273), .A3(n_239), .B(n_263), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_281), .A2(n_265), .B1(n_258), .B2(n_272), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_301), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_281), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_287), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_284), .A2(n_289), .B1(n_280), .B2(n_300), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g331 ( .A1(n_278), .A2(n_272), .B1(n_263), .B2(n_257), .C(n_268), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_287), .B(n_257), .Y(n_332) );
OAI221xp5_ASAP7_75t_SL g333 ( .A1(n_278), .A2(n_166), .B1(n_171), .B2(n_10), .C(n_13), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_303), .B(n_258), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_284), .B(n_269), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_281), .A2(n_268), .B1(n_269), .B2(n_259), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_289), .A2(n_269), .B1(n_259), .B2(n_256), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_311), .A2(n_269), .B(n_259), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_330), .B(n_281), .Y(n_341) );
OR2x6_ASAP7_75t_L g342 ( .A(n_330), .B(n_296), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_323), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_329), .B(n_288), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_339), .B(n_281), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_339), .B(n_281), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_332), .B(n_288), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_323), .B(n_281), .Y(n_348) );
CKINVDCx11_ASAP7_75t_R g349 ( .A(n_313), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_325), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_317), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g353 ( .A1(n_319), .A2(n_302), .B(n_283), .C(n_279), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_332), .B(n_288), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_317), .B(n_297), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_315), .B(n_328), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_315), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_325), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_298), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_340), .B(n_297), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_340), .B(n_291), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_325), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_321), .B(n_297), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_335), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_312), .B(n_282), .Y(n_368) );
OAI211xp5_ASAP7_75t_L g369 ( .A1(n_353), .A2(n_349), .B(n_314), .C(n_343), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_350), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_354), .B(n_335), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_343), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_313), .B1(n_316), .B2(n_318), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_341), .A2(n_313), .B1(n_346), .B2(n_345), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_347), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_357), .A2(n_316), .B1(n_322), .B2(n_326), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_358), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_354), .B(n_324), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_358), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_347), .B(n_324), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_357), .B(n_299), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_359), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_345), .B(n_336), .Y(n_384) );
OAI33xp33_ASAP7_75t_L g385 ( .A1(n_359), .A2(n_365), .A3(n_362), .B1(n_348), .B2(n_341), .B3(n_368), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_362), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_356), .A2(n_322), .B1(n_292), .B2(n_320), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_344), .B(n_333), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_356), .B(n_334), .Y(n_391) );
BUFx4f_ASAP7_75t_L g392 ( .A(n_344), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_352), .Y(n_393) );
NAND3xp33_ASAP7_75t_SL g394 ( .A(n_365), .B(n_327), .C(n_320), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_364), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_331), .B(n_320), .C(n_295), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_348), .B(n_282), .C(n_295), .D(n_320), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_345), .A2(n_292), .B1(n_334), .B2(n_298), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_346), .A2(n_292), .B1(n_298), .B2(n_337), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_367), .B(n_298), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_346), .B(n_296), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_350), .B(n_296), .Y(n_402) );
INVx5_ASAP7_75t_SL g403 ( .A(n_342), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_386), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_372), .B(n_367), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_372), .B(n_352), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_383), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_371), .B(n_355), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_377), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_378), .B(n_360), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_371), .B(n_355), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_377), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_378), .B(n_360), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_381), .B(n_8), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_375), .B(n_360), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_380), .B(n_361), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_389), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_389), .B(n_342), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_395), .B(n_342), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_395), .B(n_370), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_380), .B(n_401), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_370), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_401), .B(n_361), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_373), .A2(n_342), .B1(n_366), .B2(n_368), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_386), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_384), .B(n_342), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_393), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_384), .B(n_342), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_384), .B(n_363), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_392), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_390), .B(n_366), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_390), .B(n_363), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_369), .B(n_9), .Y(n_443) );
NAND3xp33_ASAP7_75t_SL g444 ( .A(n_373), .B(n_286), .C(n_14), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_384), .B(n_363), .Y(n_445) );
INVx4_ASAP7_75t_L g446 ( .A(n_392), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_392), .B(n_363), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_402), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g451 ( .A(n_388), .B(n_9), .C(n_14), .D(n_15), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_374), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_376), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_418), .B(n_403), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_426), .B(n_403), .Y(n_456) );
AOI221x1_ASAP7_75t_L g457 ( .A1(n_451), .A2(n_394), .B1(n_397), .B2(n_337), .C(n_338), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
AOI221x1_ASAP7_75t_L g459 ( .A1(n_451), .A2(n_397), .B1(n_391), .B2(n_385), .C(n_291), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_414), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_414), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_426), .B(n_403), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_453), .B(n_376), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_427), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_415), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_415), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_419), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_448), .B(n_388), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_449), .B(n_403), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_428), .B(n_399), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_398), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_449), .B(n_396), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_408), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_453), .B(n_15), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_421), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_420), .B(n_293), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_440), .B(n_16), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_404), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_420), .B(n_293), .Y(n_480) );
INVxp33_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_412), .B(n_16), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_417), .B(n_17), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_444), .B(n_297), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_412), .B(n_17), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_424), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_446), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_450), .B(n_293), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_409), .B(n_18), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_450), .B(n_293), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_450), .B(n_304), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_416), .B(n_19), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_413), .B(n_19), .Y(n_494) );
XNOR2xp5_ASAP7_75t_L g495 ( .A(n_452), .B(n_20), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_416), .B(n_20), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_421), .B(n_21), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_452), .A2(n_285), .B1(n_307), .B2(n_297), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_404), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_404), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_441), .B(n_21), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_443), .B(n_22), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_425), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_425), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_411), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_441), .B(n_22), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_429), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_429), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_442), .B(n_23), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_424), .B(n_23), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_405), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_405), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_433), .B(n_304), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_502), .A2(n_442), .B(n_406), .C(n_439), .Y(n_514) );
AOI21xp33_ASAP7_75t_SL g515 ( .A1(n_495), .A2(n_439), .B(n_422), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_488), .A2(n_446), .B1(n_422), .B2(n_411), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_483), .A2(n_430), .B(n_411), .C(n_423), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_479), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_485), .A2(n_446), .B(n_407), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_495), .A2(n_446), .B(n_431), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_484), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_484), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_503), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g524 ( .A1(n_459), .A2(n_448), .B(n_447), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_481), .B(n_448), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_456), .B(n_433), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_503), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_488), .Y(n_528) );
AOI31xp33_ASAP7_75t_SL g529 ( .A1(n_510), .A2(n_423), .A3(n_405), .B(n_448), .Y(n_529) );
AOI211xp5_ASAP7_75t_L g530 ( .A1(n_472), .A2(n_436), .B(n_447), .C(n_437), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_456), .B(n_436), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_464), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_510), .A2(n_431), .B1(n_438), .B2(n_432), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_468), .A2(n_445), .B1(n_437), .B2(n_438), .Y(n_534) );
AOI21xp33_ASAP7_75t_L g535 ( .A1(n_475), .A2(n_434), .B(n_432), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_459), .B(n_434), .C(n_445), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_478), .B(n_285), .C(n_307), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_455), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g539 ( .A1(n_481), .A2(n_285), .B(n_307), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_487), .B(n_24), .Y(n_540) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_470), .A2(n_304), .B(n_308), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_468), .A2(n_294), .B1(n_277), .B2(n_268), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_470), .B(n_24), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_490), .B(n_25), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_458), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_460), .Y(n_546) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_457), .A2(n_308), .B(n_26), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_471), .B(n_308), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_461), .Y(n_549) );
AOI322xp5_ASAP7_75t_L g550 ( .A1(n_471), .A2(n_291), .A3(n_256), .B1(n_269), .B2(n_259), .C1(n_294), .C2(n_277), .Y(n_550) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_497), .B(n_294), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_465), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_466), .Y(n_553) );
AOI21xp33_ASAP7_75t_SL g554 ( .A1(n_497), .A2(n_286), .B(n_28), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_457), .A2(n_286), .B(n_294), .Y(n_555) );
AOI21xp33_ASAP7_75t_L g556 ( .A1(n_501), .A2(n_294), .B(n_29), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_463), .B(n_185), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_472), .B(n_467), .Y(n_558) );
AOI211x1_ASAP7_75t_L g559 ( .A1(n_482), .A2(n_496), .B(n_493), .C(n_486), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g560 ( .A1(n_506), .A2(n_27), .B(n_30), .C(n_31), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_504), .Y(n_561) );
AOI21xp33_ASAP7_75t_SL g562 ( .A1(n_490), .A2(n_32), .B(n_36), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_507), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_508), .Y(n_564) );
OAI322xp33_ASAP7_75t_L g565 ( .A1(n_494), .A2(n_185), .A3(n_291), .B1(n_39), .B2(n_40), .C1(n_41), .C2(n_42), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_558), .B(n_473), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_521), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_530), .B(n_476), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_522), .Y(n_569) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_520), .A2(n_468), .B(n_494), .C(n_509), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_520), .A2(n_501), .B(n_474), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_532), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_533), .B(n_480), .Y(n_573) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_543), .B(n_488), .C(n_505), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_528), .B(n_462), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_526), .B(n_462), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_540), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g578 ( .A1(n_515), .A2(n_505), .B(n_469), .C(n_454), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_523), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_524), .A2(n_513), .B1(n_454), .B2(n_480), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_531), .B(n_513), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_517), .A2(n_469), .B(n_477), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_527), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_518), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_548), .B(n_477), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_533), .B(n_512), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_534), .B(n_512), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_514), .B(n_535), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_554), .A2(n_511), .B(n_500), .C(n_499), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_528), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_538), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_519), .B(n_511), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_545), .Y(n_593) );
OAI211xp5_ASAP7_75t_L g594 ( .A1(n_559), .A2(n_498), .B(n_499), .C(n_500), .Y(n_594) );
XOR2x2_ASAP7_75t_L g595 ( .A(n_544), .B(n_492), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_519), .B(n_492), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_546), .B(n_479), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_489), .B(n_491), .Y(n_598) );
NOR3xp33_ASAP7_75t_SL g599 ( .A(n_565), .B(n_37), .C(n_38), .Y(n_599) );
AOI211xp5_ASAP7_75t_SL g600 ( .A1(n_516), .A2(n_491), .B(n_489), .C(n_47), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_549), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_572), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_588), .A2(n_536), .B1(n_563), .B2(n_553), .C(n_561), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_SL g604 ( .A1(n_578), .A2(n_562), .B(n_529), .C(n_556), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_585), .B(n_564), .Y(n_605) );
XNOR2x2_ASAP7_75t_L g606 ( .A(n_595), .B(n_551), .Y(n_606) );
XNOR2xp5_ASAP7_75t_L g607 ( .A(n_595), .B(n_552), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_600), .A2(n_560), .B(n_542), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_588), .Y(n_609) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_590), .B(n_547), .Y(n_610) );
AOI211x1_ASAP7_75t_SL g611 ( .A1(n_582), .A2(n_555), .B(n_557), .C(n_529), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_589), .A2(n_547), .B(n_555), .Y(n_612) );
AO22x1_ASAP7_75t_L g613 ( .A1(n_571), .A2(n_537), .B1(n_539), .B2(n_550), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_577), .A2(n_541), .B1(n_185), .B2(n_291), .C(n_256), .Y(n_614) );
AOI211x1_ASAP7_75t_SL g615 ( .A1(n_568), .A2(n_291), .B(n_185), .C(n_48), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_574), .A2(n_268), .B1(n_256), .B2(n_185), .Y(n_616) );
AO22x2_ASAP7_75t_L g617 ( .A1(n_590), .A2(n_44), .B1(n_45), .B2(n_50), .Y(n_617) );
XNOR2x1_ASAP7_75t_L g618 ( .A(n_575), .B(n_52), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_580), .A2(n_256), .B1(n_55), .B2(n_58), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g620 ( .A(n_570), .B(n_54), .C(n_60), .D(n_66), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_567), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_569), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_594), .A2(n_68), .B(n_69), .C(n_71), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_609), .A2(n_607), .B1(n_608), .B2(n_602), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_604), .A2(n_592), .B(n_599), .C(n_573), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_605), .Y(n_626) );
NOR2xp33_ASAP7_75t_R g627 ( .A(n_618), .B(n_566), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g628 ( .A(n_611), .B(n_599), .C(n_592), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_603), .B(n_586), .C(n_593), .Y(n_629) );
NAND3xp33_ASAP7_75t_SL g630 ( .A(n_623), .B(n_598), .C(n_596), .Y(n_630) );
OAI211xp5_ASAP7_75t_L g631 ( .A1(n_620), .A2(n_587), .B(n_591), .C(n_601), .Y(n_631) );
OAI211xp5_ASAP7_75t_SL g632 ( .A1(n_615), .A2(n_579), .B(n_583), .C(n_597), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_621), .B(n_587), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_622), .B(n_575), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_606), .Y(n_635) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_628), .B(n_610), .Y(n_636) );
NAND3x1_ASAP7_75t_SL g637 ( .A(n_635), .B(n_614), .C(n_613), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_624), .A2(n_612), .B1(n_616), .B2(n_575), .Y(n_638) );
OR5x1_ASAP7_75t_L g639 ( .A(n_631), .B(n_617), .C(n_619), .D(n_576), .E(n_581), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_633), .B(n_584), .Y(n_640) );
NAND2x1p5_ASAP7_75t_L g641 ( .A(n_634), .B(n_617), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_626), .B(n_581), .Y(n_642) );
NOR3xp33_ASAP7_75t_SL g643 ( .A(n_638), .B(n_631), .C(n_625), .Y(n_643) );
XOR2xp5_ASAP7_75t_L g644 ( .A(n_641), .B(n_630), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_640), .Y(n_645) );
NOR4xp75_ASAP7_75t_L g646 ( .A(n_637), .B(n_627), .C(n_629), .D(n_632), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_645), .Y(n_647) );
NOR4xp25_ASAP7_75t_L g648 ( .A(n_646), .B(n_639), .C(n_636), .D(n_642), .Y(n_648) );
XNOR2x1_ASAP7_75t_L g649 ( .A(n_644), .B(n_584), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_647), .A2(n_643), .B(n_73), .C(n_75), .Y(n_650) );
OAI22xp5_ASAP7_75t_SL g651 ( .A1(n_648), .A2(n_643), .B1(n_79), .B2(n_81), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_650), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_652), .A2(n_651), .B1(n_649), .B2(n_648), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_653), .A2(n_72), .B(n_82), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_655) );
endmodule