module fake_jpeg_15369_n_369 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_369);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_369;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_9),
.B(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_38),
.B(n_52),
.Y(n_110)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_40),
.B(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_59),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_25),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_36),
.B(n_37),
.C(n_18),
.Y(n_83)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_25),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_27),
.B(n_13),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_12),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_92),
.Y(n_117)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_49),
.B1(n_55),
.B2(n_48),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_74),
.A2(n_76),
.B1(n_84),
.B2(n_85),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_52),
.C(n_64),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_93),
.C(n_10),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_36),
.B1(n_26),
.B2(n_37),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_38),
.A2(n_47),
.B1(n_40),
.B2(n_43),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_80),
.A2(n_114),
.B1(n_71),
.B2(n_90),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_83),
.B(n_105),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_33),
.B1(n_14),
.B2(n_18),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_88),
.B(n_103),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_111),
.B1(n_112),
.B2(n_51),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_22),
.C(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_34),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_59),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_30),
.B1(n_28),
.B2(n_14),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_97),
.A2(n_106),
.B1(n_113),
.B2(n_11),
.Y(n_147)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_62),
.B(n_30),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_28),
.B1(n_12),
.B2(n_31),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_58),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_45),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_62),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_113)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_124),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_73),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_51),
.B1(n_50),
.B2(n_62),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_125),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_126),
.A2(n_147),
.B1(n_132),
.B2(n_153),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_81),
.B(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_133),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_148),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_59),
.B1(n_3),
.B2(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_132),
.A2(n_137),
.B1(n_143),
.B2(n_155),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_1),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_75),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_7),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_138),
.B(n_141),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_9),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_10),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_125),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_10),
.B1(n_11),
.B2(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_72),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_145),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_11),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_69),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_90),
.A2(n_11),
.B1(n_114),
.B2(n_70),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_149),
.A2(n_153),
.B1(n_134),
.B2(n_168),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_126),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_73),
.C(n_108),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_142),
.C(n_150),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_156),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_71),
.A2(n_101),
.B1(n_112),
.B2(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_69),
.B(n_104),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_87),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_160),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_158),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_77),
.A2(n_86),
.B1(n_94),
.B2(n_96),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_159),
.A2(n_168),
.B1(n_152),
.B2(n_118),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_100),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_86),
.B1(n_94),
.B2(n_96),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_141),
.B(n_140),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_88),
.B(n_80),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_139),
.C(n_119),
.Y(n_177)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_170),
.B(n_188),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_173),
.A2(n_212),
.B1(n_191),
.B2(n_195),
.Y(n_232)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_180),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_176),
.B(n_177),
.Y(n_253)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_211),
.B1(n_213),
.B2(n_205),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_185),
.A2(n_190),
.B1(n_197),
.B2(n_206),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_158),
.C(n_213),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_190),
.B(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_137),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_204),
.Y(n_226)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_155),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_210),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_117),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_202),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_130),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_172),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_123),
.B(n_146),
.Y(n_210)
);

AO22x1_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_120),
.B1(n_154),
.B2(n_158),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_123),
.A2(n_120),
.B1(n_154),
.B2(n_158),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_120),
.A2(n_164),
.B1(n_125),
.B2(n_142),
.Y(n_213)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_228),
.B1(n_254),
.B2(n_230),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_236),
.C(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_187),
.B1(n_193),
.B2(n_185),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_231),
.B1(n_241),
.B2(n_222),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_225),
.A2(n_193),
.B(n_192),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_169),
.Y(n_227)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_183),
.B(n_211),
.C(n_192),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_228),
.A2(n_215),
.B(n_241),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_229),
.A2(n_250),
.B(n_226),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_184),
.B1(n_176),
.B2(n_172),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_232),
.A2(n_245),
.B1(n_243),
.B2(n_246),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_179),
.Y(n_233)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_234),
.B(n_247),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_237),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_194),
.C(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_170),
.B(n_188),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_202),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_201),
.B1(n_208),
.B2(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_243),
.B(n_248),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_191),
.A2(n_186),
.B1(n_203),
.B2(n_214),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_191),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_180),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_254),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_171),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_171),
.B(n_193),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_219),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_264),
.C(n_269),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_257),
.A2(n_260),
.B(n_268),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_226),
.A2(n_222),
.B(n_229),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_262),
.A2(n_260),
.B1(n_271),
.B2(n_261),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_231),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_230),
.A2(n_217),
.B1(n_251),
.B2(n_228),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_275),
.B1(n_277),
.B2(n_272),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_217),
.A2(n_228),
.B(n_251),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_228),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_253),
.C(n_237),
.Y(n_270)
);

HAxp5_ASAP7_75t_SL g299 ( 
.A(n_270),
.B(n_272),
.CON(n_299),
.SN(n_299)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_253),
.C(n_224),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_284),
.C(n_282),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_221),
.A2(n_216),
.B(n_218),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_238),
.B1(n_239),
.B2(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_250),
.A2(n_244),
.B(n_246),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_283),
.B(n_259),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_226),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_223),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_305),
.C(n_273),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_276),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_294),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_286),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_279),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_255),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_267),
.B(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_283),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_304),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_271),
.C(n_284),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_306),
.A2(n_296),
.B1(n_301),
.B2(n_294),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_278),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_308),
.A2(n_293),
.B1(n_296),
.B2(n_310),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_269),
.A2(n_268),
.B(n_257),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_281),
.Y(n_310)
);

INVx11_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_309),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_265),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_266),
.B1(n_264),
.B2(n_274),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_316),
.C(n_326),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_280),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_300),
.B(n_259),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_317),
.B(n_307),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_304),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_298),
.B(n_289),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_319),
.B(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_288),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_295),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_307),
.Y(n_326)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_288),
.B1(n_311),
.B2(n_297),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_335),
.B(n_331),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_314),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_312),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_SL g339 ( 
.A1(n_328),
.A2(n_299),
.A3(n_313),
.B1(n_308),
.B2(n_303),
.C1(n_297),
.C2(n_311),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_339),
.B(n_343),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_341),
.A2(n_318),
.B(n_320),
.Y(n_348)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_330),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_291),
.Y(n_343)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_345),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_348),
.B(n_350),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_335),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_332),
.A2(n_329),
.B(n_319),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_315),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_353),
.B(n_340),
.C(n_338),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_346),
.A2(n_334),
.B1(n_342),
.B2(n_324),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_359),
.C(n_352),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_352),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_347),
.B(n_344),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_361),
.C(n_357),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_351),
.B(n_356),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_363),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_366),
.B(n_355),
.C(n_348),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_362),
.B(n_364),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_353),
.Y(n_369)
);


endmodule