module real_jpeg_2773_n_16 (n_5, n_4, n_8, n_0, n_12, n_378, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_378;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_1),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_1),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_1),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_1),
.B(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_3),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_3),
.B(n_33),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_38),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_53),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_3),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_3),
.B(n_42),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_3),
.B(n_71),
.Y(n_308)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_4),
.B(n_42),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_4),
.B(n_71),
.Y(n_254)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_5),
.B(n_53),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_5),
.B(n_38),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_60),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_68),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_11),
.B(n_42),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_11),
.B(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_11),
.B(n_33),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_11),
.B(n_53),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_60),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_11),
.B(n_68),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_13),
.B(n_68),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_13),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_13),
.B(n_60),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_71),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_13),
.B(n_33),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_13),
.B(n_53),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_13),
.B(n_38),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_13),
.B(n_30),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_14),
.B(n_68),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_14),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_14),
.B(n_42),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_14),
.B(n_33),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_42),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_15),
.B(n_53),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_15),
.B(n_60),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_15),
.B(n_71),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_358),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_156),
.B(n_357),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_19),
.B(n_134),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_82),
.C(n_101),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_20),
.B(n_82),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_63),
.B2(n_81),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_21),
.B(n_64),
.C(n_73),
.Y(n_155)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_47),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_23),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_32),
.C(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_28),
.B(n_37),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_29),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_29),
.B(n_39),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_29),
.B(n_171),
.Y(n_289)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_66),
.C(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_32),
.A2(n_34),
.B1(n_66),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_32),
.A2(n_34),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_32),
.B(n_188),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_33),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_35),
.A2(n_36),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_35),
.B(n_288),
.C(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_37),
.B(n_171),
.Y(n_194)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_39),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_40),
.A2(n_47),
.B1(n_48),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_40),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.C(n_46),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_41),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_46),
.Y(n_119)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_55),
.B2(n_62),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_50),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_49),
.A2(n_50),
.B1(n_125),
.B2(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_49),
.B(n_227),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_56),
.C(n_59),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_50),
.B(n_85),
.C(n_88),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_52),
.B(n_171),
.Y(n_198)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_56),
.A2(n_57),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_60),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_73),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.C(n_70),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_66),
.A2(n_108),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_66),
.B(n_244),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_67),
.A2(n_109),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_68),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_69),
.A2(n_70),
.B1(n_80),
.B2(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_70),
.B(n_74),
.C(n_77),
.Y(n_148)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_71),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_79),
.B(n_123),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_91),
.C(n_92),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_84),
.A2(n_85),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_84),
.A2(n_85),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_85),
.B(n_238),
.C(n_239),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_85),
.B(n_138),
.C(n_141),
.Y(n_370)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_88),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_100),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_111),
.C(n_113),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_98),
.C(n_100),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_96),
.A2(n_97),
.B1(n_113),
.B2(n_114),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_101),
.A2(n_102),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_120),
.C(n_131),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_103),
.A2(n_104),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.C(n_115),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_105),
.B(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_109),
.B(n_150),
.C(n_152),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_110),
.B(n_115),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_111),
.B(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_112),
.B(n_266),
.Y(n_372)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_120),
.B(n_131),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.C(n_129),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_121),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.C(n_125),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_122),
.A2(n_125),
.B1(n_227),
.B2(n_301),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_122),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_123),
.B(n_126),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_123),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_124),
.A2(n_299),
.B1(n_300),
.B2(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_124),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_124),
.A2(n_137),
.B1(n_138),
.B2(n_299),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_125),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_328)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_134),
.B(n_360),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_134),
.B(n_360),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_146),
.CI(n_155),
.CON(n_134),
.SN(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_136),
.B(n_144),
.C(n_145),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_138),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_138),
.B(n_280),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_148),
.B(n_149),
.C(n_154),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

AOI321xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_334),
.A3(n_346),
.B1(n_351),
.B2(n_356),
.C(n_378),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_291),
.C(n_330),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_258),
.B(n_290),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_230),
.B(n_257),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_210),
.B(n_229),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_191),
.B(n_209),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_173),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.C(n_172),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_164),
.A2(n_165),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_183),
.C(n_187),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_221),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_186),
.B1(n_187),
.B2(n_190),
.Y(n_182)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_200),
.B(n_208),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_196),
.B(n_199),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_201),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_212),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_222),
.C(n_223),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_217),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_232),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_246),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_247),
.C(n_248),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_240),
.B2(n_241),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_242),
.C(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_256),
.Y(n_248)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_254),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_259),
.B(n_260),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_277),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_275),
.B2(n_276),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_263),
.B(n_276),
.C(n_277),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_272),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_273),
.C(n_274),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_269),
.C(n_271),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_285),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_306),
.C(n_309),
.Y(n_326)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_283),
.C(n_285),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g352 ( 
.A1(n_292),
.A2(n_353),
.B(n_354),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_319),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_293),
.B(n_319),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_310),
.C(n_311),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_297),
.C(n_304),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_303),
.B2(n_304),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_308),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_311),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_316),
.C(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_329),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_323),
.C(n_329),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_326),
.C(n_327),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_332),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_343),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_335),
.B(n_343),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.C(n_342),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_339),
.Y(n_350)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_347),
.A2(n_352),
.B(n_355),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_348),
.B(n_349),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_375),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_374),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);


endmodule