module real_aes_6312_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_762;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g237 ( .A1(n_0), .A2(n_238), .B(n_239), .C(n_243), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_1), .B(n_179), .Y(n_244) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_3), .B(n_151), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_4), .A2(n_137), .B(n_142), .C(n_505), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_5), .A2(n_132), .B(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_6), .A2(n_132), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_7), .B(n_179), .Y(n_549) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_8), .A2(n_167), .B(n_183), .Y(n_182) );
AND2x6_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_10), .A2(n_137), .B(n_142), .C(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g487 ( .A(n_11), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_12), .B(n_42), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_12), .B(n_42), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_13), .B(n_242), .Y(n_507) );
INVx1_ASAP7_75t_L g161 ( .A(n_14), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_15), .B(n_151), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_16), .A2(n_152), .B(n_495), .C(n_497), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_17), .B(n_179), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_18), .A2(n_468), .B1(n_746), .B2(n_752), .C1(n_755), .C2(n_756), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_19), .B(n_216), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_20), .A2(n_142), .B(n_193), .C(n_212), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_21), .A2(n_191), .B(n_241), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_22), .B(n_242), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_23), .A2(n_104), .B1(n_114), .B2(n_762), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_24), .B(n_242), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_25), .Y(n_534) );
INVx1_ASAP7_75t_L g526 ( .A(n_26), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_27), .A2(n_142), .B(n_186), .C(n_193), .Y(n_185) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_29), .Y(n_503) );
INVx1_ASAP7_75t_L g583 ( .A(n_30), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_31), .A2(n_132), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g135 ( .A(n_32), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_33), .A2(n_140), .B(n_155), .C(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_34), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_35), .A2(n_241), .B(n_546), .C(n_548), .Y(n_545) );
INVxp67_ASAP7_75t_L g584 ( .A(n_36), .Y(n_584) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_37), .A2(n_47), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_38), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_39), .A2(n_142), .B(n_193), .C(n_525), .Y(n_524) );
CKINVDCx14_ASAP7_75t_R g544 ( .A(n_40), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_41), .A2(n_46), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_41), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_43), .A2(n_243), .B(n_485), .C(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_44), .B(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_45), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_46), .Y(n_750) );
INVx1_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
OAI321xp33_ASAP7_75t_L g120 ( .A1(n_48), .A2(n_121), .A3(n_455), .B1(n_461), .B2(n_462), .C(n_464), .Y(n_120) );
INVx1_ASAP7_75t_L g461 ( .A(n_48), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_49), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_50), .B(n_132), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_51), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_52), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_53), .A2(n_140), .B(n_145), .C(n_155), .Y(n_139) );
INVx1_ASAP7_75t_L g240 ( .A(n_54), .Y(n_240) );
INVx1_ASAP7_75t_L g146 ( .A(n_55), .Y(n_146) );
INVx1_ASAP7_75t_L g515 ( .A(n_56), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_57), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_58), .B(n_132), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_59), .Y(n_219) );
CKINVDCx14_ASAP7_75t_R g483 ( .A(n_60), .Y(n_483) );
INVx1_ASAP7_75t_L g138 ( .A(n_61), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_62), .B(n_132), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_63), .B(n_179), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_64), .A2(n_173), .B(n_175), .C(n_177), .Y(n_172) );
INVx1_ASAP7_75t_L g160 ( .A(n_65), .Y(n_160) );
INVx1_ASAP7_75t_SL g547 ( .A(n_66), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_68), .B(n_151), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_69), .B(n_179), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_70), .B(n_152), .Y(n_254) );
INVx1_ASAP7_75t_L g537 ( .A(n_71), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_72), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_73), .B(n_148), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_74), .A2(n_142), .B(n_155), .C(n_225), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_75), .Y(n_171) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_77), .A2(n_132), .B(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_78), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_79), .A2(n_132), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_80), .A2(n_210), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g493 ( .A(n_81), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_82), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_83), .B(n_147), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_84), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_84), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_85), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_86), .A2(n_132), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g496 ( .A(n_87), .Y(n_496) );
INVx2_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g506 ( .A(n_89), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_90), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_91), .B(n_242), .Y(n_255) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_92), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g457 ( .A(n_92), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g474 ( .A(n_92), .Y(n_474) );
OR2x2_ASAP7_75t_L g745 ( .A(n_92), .B(n_459), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_93), .A2(n_142), .B(n_155), .C(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_94), .B(n_132), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_95), .Y(n_202) );
INVxp67_ASAP7_75t_L g176 ( .A(n_96), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_97), .B(n_167), .Y(n_488) );
INVx2_ASAP7_75t_L g518 ( .A(n_98), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_99), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g226 ( .A(n_100), .Y(n_226) );
INVx1_ASAP7_75t_L g250 ( .A(n_101), .Y(n_250) );
AND2x2_ASAP7_75t_L g162 ( .A(n_102), .B(n_157), .Y(n_162) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g763 ( .A(n_107), .Y(n_763) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g459 ( .A(n_110), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_466), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g761 ( .A(n_118), .Y(n_761) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_121), .B(n_463), .Y(n_462) );
XOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_125), .A2(n_470), .B1(n_475), .B2(n_742), .Y(n_469) );
INVx4_ASAP7_75t_L g759 ( .A(n_125), .Y(n_759) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR5x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_328), .C(n_406), .D(n_430), .E(n_447), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_194), .B(n_245), .C(n_305), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
AND2x2_ASAP7_75t_L g259 ( .A(n_129), .B(n_165), .Y(n_259) );
INVx5_ASAP7_75t_SL g287 ( .A(n_129), .Y(n_287) );
AND2x2_ASAP7_75t_L g323 ( .A(n_129), .B(n_308), .Y(n_323) );
OR2x2_ASAP7_75t_L g362 ( .A(n_129), .B(n_164), .Y(n_362) );
OR2x2_ASAP7_75t_L g393 ( .A(n_129), .B(n_284), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_129), .B(n_297), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_129), .B(n_284), .Y(n_441) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_162), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_139), .B(n_157), .Y(n_130) );
BUFx2_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_133), .B(n_137), .Y(n_251) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx1_ASAP7_75t_L g192 ( .A(n_135), .Y(n_192) );
INVx1_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
INVx1_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_136), .Y(n_242) );
INVx4_ASAP7_75t_SL g156 ( .A(n_137), .Y(n_156) );
BUFx3_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_141), .A2(n_156), .B(n_171), .C(n_172), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_141), .A2(n_156), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_141), .A2(n_156), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_141), .A2(n_156), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_141), .A2(n_156), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_141), .A2(n_156), .B(n_544), .C(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_SL g579 ( .A1(n_141), .A2(n_156), .B(n_580), .C(n_581), .Y(n_579) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_143), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .C(n_153), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_147), .A2(n_153), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp5_ASAP7_75t_L g505 ( .A1(n_147), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_147), .A2(n_508), .B(n_537), .C(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_151), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g238 ( .A(n_151), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_151), .A2(n_215), .B(n_526), .C(n_527), .Y(n_525) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_151), .A2(n_174), .B1(n_583), .B2(n_584), .Y(n_582) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_152), .B(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g243 ( .A(n_154), .Y(n_243) );
INVx1_ASAP7_75t_L g497 ( .A(n_154), .Y(n_497) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_157), .A2(n_199), .B(n_200), .Y(n_198) );
INVx2_ASAP7_75t_L g217 ( .A(n_157), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_157), .A2(n_481), .B(n_488), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_157), .A2(n_251), .B(n_523), .C(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g168 ( .A(n_158), .B(n_159), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AND2x2_ASAP7_75t_L g440 ( .A(n_163), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
OR2x2_ASAP7_75t_L g303 ( .A(n_164), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_181), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_165), .B(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_165), .Y(n_296) );
INVx3_ASAP7_75t_L g311 ( .A(n_165), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_165), .B(n_181), .Y(n_335) );
OR2x2_ASAP7_75t_L g344 ( .A(n_165), .B(n_287), .Y(n_344) );
AND2x2_ASAP7_75t_L g348 ( .A(n_165), .B(n_308), .Y(n_348) );
AND2x2_ASAP7_75t_L g354 ( .A(n_165), .B(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g391 ( .A(n_165), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_165), .B(n_248), .Y(n_405) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_178), .Y(n_165) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_166), .A2(n_491), .B(n_498), .Y(n_490) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_166), .A2(n_513), .B(n_519), .Y(n_512) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_166), .A2(n_542), .B(n_549), .Y(n_541) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_167), .A2(n_184), .B(n_185), .Y(n_183) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g258 ( .A(n_168), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_173), .A2(n_226), .B(n_227), .C(n_228), .Y(n_225) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_174), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_174), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g215 ( .A(n_177), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_177), .B(n_582), .Y(n_581) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_179), .A2(n_234), .B(n_244), .Y(n_233) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_180), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_180), .A2(n_223), .B(n_231), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_180), .B(n_232), .Y(n_231) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_180), .A2(n_249), .B(n_256), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_180), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_180), .B(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_180), .A2(n_533), .B(n_539), .Y(n_532) );
OR2x2_ASAP7_75t_L g297 ( .A(n_181), .B(n_248), .Y(n_297) );
AND2x2_ASAP7_75t_L g308 ( .A(n_181), .B(n_284), .Y(n_308) );
AND2x2_ASAP7_75t_L g320 ( .A(n_181), .B(n_311), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_181), .B(n_248), .Y(n_343) );
INVx1_ASAP7_75t_SL g355 ( .A(n_181), .Y(n_355) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g247 ( .A(n_182), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_182), .B(n_287), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B(n_190), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_190), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
AND2x2_ASAP7_75t_L g268 ( .A(n_196), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_196), .B(n_221), .Y(n_272) );
AND2x2_ASAP7_75t_L g275 ( .A(n_196), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_196), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g300 ( .A(n_196), .B(n_291), .Y(n_300) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_196), .Y(n_319) );
AND2x2_ASAP7_75t_L g340 ( .A(n_196), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g350 ( .A(n_196), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g396 ( .A(n_196), .B(n_279), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_196), .B(n_302), .Y(n_423) );
INVx5_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g293 ( .A(n_197), .Y(n_293) );
AND2x2_ASAP7_75t_L g359 ( .A(n_197), .B(n_291), .Y(n_359) );
AND2x2_ASAP7_75t_L g443 ( .A(n_197), .B(n_311), .Y(n_443) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_204), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_206), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_206), .Y(n_432) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_221), .Y(n_206) );
AND2x2_ASAP7_75t_L g262 ( .A(n_207), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g271 ( .A(n_207), .B(n_269), .Y(n_271) );
INVx5_ASAP7_75t_L g279 ( .A(n_207), .Y(n_279) );
AND2x2_ASAP7_75t_L g302 ( .A(n_207), .B(n_233), .Y(n_302) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_207), .Y(n_339) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_211), .B(n_216), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_217), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_220), .A2(n_502), .B(n_509), .Y(n_501) );
INVx1_ASAP7_75t_L g380 ( .A(n_221), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_221), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g413 ( .A(n_221), .B(n_279), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_221), .A2(n_336), .B(n_443), .C(n_444), .Y(n_442) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_233), .Y(n_221) );
BUFx2_ASAP7_75t_L g263 ( .A(n_222), .Y(n_263) );
INVx2_ASAP7_75t_L g267 ( .A(n_222), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g548 ( .A(n_229), .Y(n_548) );
INVx2_ASAP7_75t_L g269 ( .A(n_233), .Y(n_269) );
AND2x2_ASAP7_75t_L g276 ( .A(n_233), .B(n_267), .Y(n_276) );
AND2x2_ASAP7_75t_L g367 ( .A(n_233), .B(n_279), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_241), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g485 ( .A(n_242), .Y(n_485) );
INVx2_ASAP7_75t_L g508 ( .A(n_243), .Y(n_508) );
AOI211x1_ASAP7_75t_SL g245 ( .A1(n_246), .A2(n_260), .B(n_273), .C(n_298), .Y(n_245) );
INVx1_ASAP7_75t_L g364 ( .A(n_246), .Y(n_364) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_259), .Y(n_246) );
INVx5_ASAP7_75t_SL g284 ( .A(n_248), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_248), .B(n_354), .Y(n_353) );
AOI311xp33_ASAP7_75t_L g372 ( .A1(n_248), .A2(n_373), .A3(n_375), .B(n_376), .C(n_382), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_248), .A2(n_320), .B(n_408), .C(n_411), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_252), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_251), .A2(n_503), .B(n_504), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_251), .A2(n_534), .B(n_535), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g576 ( .A(n_258), .Y(n_576) );
INVxp67_ASAP7_75t_L g327 ( .A(n_259), .Y(n_327) );
NAND4xp25_ASAP7_75t_SL g260 ( .A(n_261), .B(n_264), .C(n_270), .D(n_272), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_261), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g318 ( .A(n_262), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_265), .B(n_271), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_265), .B(n_278), .Y(n_398) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_266), .B(n_279), .Y(n_416) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g291 ( .A(n_267), .Y(n_291) );
INVxp67_ASAP7_75t_L g326 ( .A(n_268), .Y(n_326) );
AND2x4_ASAP7_75t_L g278 ( .A(n_269), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g352 ( .A(n_269), .B(n_291), .Y(n_352) );
INVx1_ASAP7_75t_L g379 ( .A(n_269), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_269), .B(n_366), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_270), .B(n_340), .Y(n_360) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_271), .B(n_293), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_271), .B(n_340), .Y(n_439) );
INVx1_ASAP7_75t_L g450 ( .A(n_272), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B(n_280), .C(n_288), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g292 ( .A(n_276), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g330 ( .A(n_276), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
AND2x2_ASAP7_75t_L g289 ( .A(n_278), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_278), .B(n_340), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_278), .B(n_359), .Y(n_383) );
OR2x2_ASAP7_75t_L g299 ( .A(n_279), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_279), .B(n_291), .Y(n_346) );
AND2x2_ASAP7_75t_L g403 ( .A(n_279), .B(n_359), .Y(n_403) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_279), .Y(n_410) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_281), .A2(n_293), .B1(n_415), .B2(n_417), .C(n_420), .Y(n_414) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g304 ( .A(n_284), .B(n_287), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_284), .B(n_354), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_284), .B(n_311), .Y(n_419) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g404 ( .A(n_286), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g418 ( .A(n_286), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_287), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g315 ( .A(n_287), .B(n_308), .Y(n_315) );
AND2x2_ASAP7_75t_L g385 ( .A(n_287), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_287), .B(n_334), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_287), .B(n_435), .Y(n_434) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_292), .B(n_294), .Y(n_288) );
INVx2_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g341 ( .A(n_291), .Y(n_341) );
OR2x2_ASAP7_75t_L g345 ( .A(n_293), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g448 ( .A(n_293), .B(n_416), .Y(n_448) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AOI21xp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_301), .B(n_303), .Y(n_298) );
INVx1_ASAP7_75t_L g452 ( .A(n_299), .Y(n_452) );
INVx2_ASAP7_75t_SL g366 ( .A(n_300), .Y(n_366) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_303), .A2(n_384), .B(n_448), .C(n_449), .Y(n_447) );
OAI322xp33_ASAP7_75t_SL g316 ( .A1(n_304), .A2(n_317), .A3(n_320), .B1(n_321), .B2(n_322), .C1(n_324), .C2(n_327), .Y(n_316) );
INVx2_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_312), .B1(n_313), .B2(n_315), .C(n_316), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp33_ASAP7_75t_SL g382 ( .A1(n_307), .A2(n_383), .B1(n_384), .B2(n_387), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_308), .B(n_311), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_308), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g381 ( .A(n_310), .B(n_343), .Y(n_381) );
INVx1_ASAP7_75t_L g371 ( .A(n_311), .Y(n_371) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_315), .A2(n_425), .B(n_427), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g349 ( .A1(n_317), .A2(n_350), .B(n_353), .Y(n_349) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp67_ASAP7_75t_SL g378 ( .A(n_319), .B(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_319), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g435 ( .A(n_320), .Y(n_435) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g328 ( .A(n_329), .B(n_356), .C(n_372), .D(n_388), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_337), .C(n_349), .Y(n_329) );
INVx1_ASAP7_75t_L g421 ( .A(n_330), .Y(n_421) );
AND2x2_ASAP7_75t_L g369 ( .A(n_331), .B(n_352), .Y(n_369) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_336), .B(n_371), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_342), .B1(n_345), .B2(n_347), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_339), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g387 ( .A(n_340), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_340), .A2(n_379), .B(n_402), .C(n_404), .Y(n_401) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g386 ( .A(n_343), .Y(n_386) );
INVx1_ASAP7_75t_L g446 ( .A(n_344), .Y(n_446) );
NAND2xp33_ASAP7_75t_SL g436 ( .A(n_345), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g375 ( .A(n_354), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_361), .C(n_363), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_368), .B2(n_370), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_366), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_371), .B(n_392), .Y(n_454) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI21xp33_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_380), .B(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_394), .B1(n_397), .B2(n_399), .C(n_401), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_404), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_420) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_414), .C(n_424), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B(n_433), .C(n_442), .Y(n_430) );
INVx1_ASAP7_75t_L g451 ( .A(n_431), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_438), .B2(n_440), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_452), .B2(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g463 ( .A(n_457), .Y(n_463) );
NOR2x2_ASAP7_75t_L g754 ( .A(n_458), .B(n_474), .Y(n_754) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g473 ( .A(n_459), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g465 ( .A(n_463), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_464), .B(n_467), .C(n_760), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI22x1_ASAP7_75t_SL g757 ( .A1(n_470), .A2(n_742), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g758 ( .A(n_475), .Y(n_758) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_672), .Y(n_475) );
NAND5xp2_ASAP7_75t_L g476 ( .A(n_477), .B(n_587), .C(n_619), .D(n_636), .E(n_659), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_520), .B1(n_550), .B2(n_554), .C(n_558), .Y(n_477) );
INVx1_ASAP7_75t_L g699 ( .A(n_478), .Y(n_699) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_499), .Y(n_478) );
AND3x2_ASAP7_75t_L g674 ( .A(n_479), .B(n_501), .C(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_480), .B(n_556), .Y(n_555) );
BUFx3_ASAP7_75t_L g565 ( .A(n_480), .Y(n_565) );
AND2x2_ASAP7_75t_L g569 ( .A(n_480), .B(n_511), .Y(n_569) );
INVx2_ASAP7_75t_L g596 ( .A(n_480), .Y(n_596) );
OR2x2_ASAP7_75t_L g607 ( .A(n_480), .B(n_512), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_480), .B(n_500), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_480), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g686 ( .A(n_480), .B(n_512), .Y(n_686) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_489), .Y(n_568) );
AND2x2_ASAP7_75t_L g627 ( .A(n_489), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_489), .B(n_500), .Y(n_646) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g557 ( .A(n_490), .B(n_500), .Y(n_557) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
AND2x2_ASAP7_75t_L g613 ( .A(n_490), .B(n_512), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_490), .B(n_499), .C(n_596), .Y(n_638) );
AND2x2_ASAP7_75t_L g703 ( .A(n_490), .B(n_501), .Y(n_703) );
AND2x2_ASAP7_75t_L g737 ( .A(n_490), .B(n_500), .Y(n_737) );
INVxp67_ASAP7_75t_L g566 ( .A(n_499), .Y(n_566) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_500), .B(n_596), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_500), .B(n_627), .Y(n_635) );
AND2x2_ASAP7_75t_L g685 ( .A(n_500), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g713 ( .A(n_500), .Y(n_713) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g620 ( .A(n_501), .B(n_613), .Y(n_620) );
BUFx3_ASAP7_75t_L g652 ( .A(n_501), .Y(n_652) );
INVx2_ASAP7_75t_L g628 ( .A(n_511), .Y(n_628) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_512), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_520), .A2(n_688), .B1(n_690), .B2(n_691), .Y(n_687) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
AND2x2_ASAP7_75t_L g550 ( .A(n_521), .B(n_551), .Y(n_550) );
INVx3_ASAP7_75t_SL g561 ( .A(n_521), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_521), .B(n_591), .Y(n_623) );
OR2x2_ASAP7_75t_L g642 ( .A(n_521), .B(n_531), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_521), .B(n_599), .Y(n_647) );
AND2x2_ASAP7_75t_L g650 ( .A(n_521), .B(n_592), .Y(n_650) );
AND2x2_ASAP7_75t_L g662 ( .A(n_521), .B(n_541), .Y(n_662) );
AND2x2_ASAP7_75t_L g678 ( .A(n_521), .B(n_532), .Y(n_678) );
AND2x4_ASAP7_75t_L g681 ( .A(n_521), .B(n_552), .Y(n_681) );
OR2x2_ASAP7_75t_L g698 ( .A(n_521), .B(n_634), .Y(n_698) );
OR2x2_ASAP7_75t_L g729 ( .A(n_521), .B(n_574), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_521), .B(n_657), .Y(n_731) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
AND2x2_ASAP7_75t_L g605 ( .A(n_530), .B(n_572), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_530), .B(n_592), .Y(n_724) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_541), .Y(n_530) );
AND2x2_ASAP7_75t_L g560 ( .A(n_531), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g599 ( .A(n_531), .B(n_574), .Y(n_599) );
AND2x2_ASAP7_75t_L g617 ( .A(n_531), .B(n_552), .Y(n_617) );
OR2x2_ASAP7_75t_L g634 ( .A(n_531), .B(n_592), .Y(n_634) );
INVx2_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g553 ( .A(n_532), .Y(n_553) );
AND2x2_ASAP7_75t_L g657 ( .A(n_532), .B(n_541), .Y(n_657) );
INVx2_ASAP7_75t_L g552 ( .A(n_541), .Y(n_552) );
INVx1_ASAP7_75t_L g669 ( .A(n_541), .Y(n_669) );
AND2x2_ASAP7_75t_L g719 ( .A(n_541), .B(n_561), .Y(n_719) );
AND2x2_ASAP7_75t_L g571 ( .A(n_551), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g603 ( .A(n_551), .B(n_561), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_551), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g590 ( .A(n_552), .B(n_561), .Y(n_590) );
OR2x2_ASAP7_75t_L g706 ( .A(n_553), .B(n_680), .Y(n_706) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_556), .B(n_686), .Y(n_692) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_557), .A2(n_649), .A3(n_651), .B1(n_653), .B2(n_654), .Y(n_648) );
OR2x2_ASAP7_75t_L g665 ( .A(n_557), .B(n_607), .Y(n_665) );
OAI21xp33_ASAP7_75t_SL g690 ( .A1(n_557), .A2(n_567), .B(n_595), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B1(n_567), .B2(n_570), .Y(n_558) );
INVxp33_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_560), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_561), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_561), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g716 ( .A(n_561), .B(n_657), .Y(n_716) );
OR2x2_ASAP7_75t_L g740 ( .A(n_561), .B(n_634), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g723 ( .A1(n_562), .A2(n_622), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g600 ( .A(n_564), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_564), .B(n_569), .Y(n_618) );
AND2x2_ASAP7_75t_L g640 ( .A(n_565), .B(n_613), .Y(n_640) );
INVx1_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
OR2x2_ASAP7_75t_L g658 ( .A(n_565), .B(n_592), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_568), .B(n_607), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_569), .A2(n_589), .B1(n_594), .B2(n_598), .Y(n_588) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_572), .A2(n_631), .B1(n_638), .B2(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g715 ( .A(n_572), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_574), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g734 ( .A(n_574), .B(n_617), .Y(n_734) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .B(n_585), .Y(n_574) );
INVx1_ASAP7_75t_L g593 ( .A(n_575), .Y(n_593) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OA21x2_ASAP7_75t_L g592 ( .A1(n_578), .A2(n_586), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_600), .B1(n_601), .B2(n_606), .C(n_608), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_590), .B(n_592), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_590), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g609 ( .A(n_591), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_591), .A2(n_697), .B(n_698), .C(n_699), .Y(n_696) );
AND2x2_ASAP7_75t_L g701 ( .A(n_591), .B(n_681), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_SL g739 ( .A1(n_591), .A2(n_680), .B(n_740), .C(n_741), .Y(n_739) );
BUFx3_ASAP7_75t_L g631 ( .A(n_592), .Y(n_631) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_595), .B(n_652), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g714 ( .A1(n_595), .A2(n_715), .B(n_717), .C(n_723), .Y(n_714) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVxp67_ASAP7_75t_L g675 ( .A(n_597), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_599), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g619 ( .A1(n_603), .A2(n_620), .B(n_621), .C(n_629), .Y(n_619) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g704 ( .A(n_607), .Y(n_704) );
OR2x2_ASAP7_75t_L g721 ( .A(n_607), .B(n_651), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_615), .B2(n_618), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_610), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
OR2x2_ASAP7_75t_L g708 ( .A(n_612), .B(n_652), .Y(n_708) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g663 ( .A(n_613), .B(n_653), .Y(n_663) );
INVx1_ASAP7_75t_L g671 ( .A(n_614), .Y(n_671) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_617), .B(n_631), .Y(n_679) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_627), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g736 ( .A(n_628), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_635), .Y(n_629) );
INVx1_ASAP7_75t_L g666 ( .A(n_630), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_631), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_631), .B(n_662), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_631), .B(n_657), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_631), .B(n_678), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_631), .A2(n_641), .B(n_681), .C(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_641), .B1(n_643), .B2(n_647), .C(n_648), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_645), .B(n_653), .Y(n_727) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g738 ( .A1(n_647), .A2(n_662), .B(n_664), .C(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_650), .B(n_657), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_651), .B(n_704), .Y(n_741) );
CKINVDCx16_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
INVxp33_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g667 ( .A1(n_656), .A2(n_668), .B(n_670), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_656), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_657), .B(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B1(n_664), .B2(n_666), .C(n_667), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_663), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g697 ( .A(n_669), .Y(n_697) );
NAND5xp2_ASAP7_75t_L g672 ( .A(n_673), .B(n_700), .C(n_714), .D(n_725), .E(n_738), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B(n_683), .C(n_696), .Y(n_673) );
INVx2_ASAP7_75t_SL g720 ( .A(n_674), .Y(n_720) );
NAND4xp25_ASAP7_75t_SL g676 ( .A(n_677), .B(n_679), .C(n_680), .D(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_682), .A2(n_684), .B(n_687), .C(n_693), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_685), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_685), .A2(n_726), .B1(n_728), .B2(n_730), .C(n_732), .Y(n_725) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_SL g700 ( .A1(n_701), .A2(n_702), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_700) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_708), .A2(n_731), .B1(n_733), .B2(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_746), .Y(n_755) );
CKINVDCx16_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
endmodule