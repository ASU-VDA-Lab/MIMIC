module real_jpeg_4100_n_29 (n_17, n_8, n_0, n_21, n_168, n_2, n_10, n_175, n_9, n_12, n_24, n_166, n_170, n_6, n_28, n_171, n_169, n_167, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_26, n_27, n_20, n_19, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_10;
input n_175;
input n_9;
input n_12;
input n_24;
input n_166;
input n_170;
input n_6;
input n_28;
input n_171;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_131;
wire n_47;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_1),
.B(n_49),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_3),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_4),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_4),
.B(n_72),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_122),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_6),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_7),
.B(n_108),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_9),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_9),
.B(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_9),
.B(n_32),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_9),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_10),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_11),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_148),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_13),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_14),
.B(n_53),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_15),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_15),
.B(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_69),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_17),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_18),
.B(n_59),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_19),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_20),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_21),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_23),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_23),
.B(n_43),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_24),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_24),
.B(n_131),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_26),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_27),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_28),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_154),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_38),
.B(n_153),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_34),
.B(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_36),
.B(n_93),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_143),
.B(n_150),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_124),
.B(n_137),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_64),
.B(n_112),
.C(n_121),
.Y(n_40)
);

NOR4xp25_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.C(n_52),
.D(n_58),
.Y(n_41)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_45),
.B(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_47),
.Y(n_162)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_52),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_55),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_55),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_55),
.B(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_88),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_107),
.B(n_111),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_99),
.B(n_106),
.Y(n_65)
);

AO221x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_74),
.B1(n_96),
.B2(n_97),
.C(n_98),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_81),
.B(n_95),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_80),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B(n_94),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_90),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_105),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B(n_118),
.C(n_119),
.D(n_120),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_133),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_133),
.B(n_138),
.C(n_141),
.D(n_142),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_136),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_163),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_166),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_167),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_168),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_169),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_170),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_171),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_172),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_173),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_174),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_175),
.Y(n_109)
);


endmodule