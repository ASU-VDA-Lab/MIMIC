module fake_jpeg_24124_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_72),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_26),
.Y(n_102)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_76),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_40),
.B(n_41),
.C(n_44),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_81),
.B1(n_88),
.B2(n_28),
.Y(n_120)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_82),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_42),
.B(n_18),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_34),
.B1(n_18),
.B2(n_30),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_34),
.B1(n_19),
.B2(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_97),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_93),
.B1(n_56),
.B2(n_62),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_44),
.B1(n_40),
.B2(n_20),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_50),
.B1(n_62),
.B2(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_108),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_105),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_131),
.B1(n_96),
.B2(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_111),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_75),
.Y(n_111)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_120),
.B1(n_20),
.B2(n_24),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_121),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_33),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_92),
.B(n_23),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_25),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_79),
.B1(n_97),
.B2(n_50),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_87),
.B1(n_20),
.B2(n_24),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_28),
.B1(n_19),
.B2(n_31),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_94),
.B1(n_83),
.B2(n_82),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_137),
.B1(n_140),
.B2(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_123),
.B1(n_111),
.B2(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_151),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_98),
.B(n_99),
.C(n_76),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_131),
.A3(n_127),
.B1(n_121),
.B2(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_156),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_31),
.B(n_73),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_26),
.B(n_29),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_101),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_48),
.C(n_46),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_119),
.C(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_35),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_105),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_113),
.Y(n_168)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_160),
.A2(n_175),
.B1(n_144),
.B2(n_112),
.Y(n_213)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_161),
.B(n_172),
.Y(n_202)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_183),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_102),
.B1(n_113),
.B2(n_125),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_178),
.B1(n_189),
.B2(n_144),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_109),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_155),
.B(n_138),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_104),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_24),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_181),
.C(n_48),
.Y(n_206)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_173),
.B(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_100),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_141),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_113),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_180),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_128),
.B1(n_116),
.B2(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_128),
.C(n_114),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_142),
.B(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_17),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_116),
.B1(n_23),
.B2(n_27),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_150),
.B1(n_152),
.B2(n_144),
.Y(n_193)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_188),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_119),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_119),
.B1(n_27),
.B2(n_29),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_162),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_184),
.A2(n_148),
.B1(n_151),
.B2(n_135),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_217),
.B1(n_185),
.B2(n_175),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_193),
.A2(n_213),
.B1(n_221),
.B2(n_163),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_207),
.B(n_219),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_133),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_35),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_210),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_216),
.C(n_220),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_20),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_181),
.Y(n_215)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_118),
.C(n_155),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_159),
.A2(n_118),
.B1(n_32),
.B2(n_33),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_169),
.Y(n_218)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_33),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_118),
.C(n_46),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_159),
.B1(n_164),
.B2(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_245),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_182),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_160),
.B1(n_186),
.B2(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_32),
.C(n_17),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_240),
.C(n_206),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_24),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_201),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_220),
.A2(n_200),
.B1(n_217),
.B2(n_198),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_247),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_249),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_207),
.B(n_204),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_191),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_251),
.B(n_232),
.Y(n_282)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_257),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_203),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_261),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_223),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_228),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_230),
.B(n_236),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_268),
.B1(n_229),
.B2(n_245),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_225),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_199),
.C(n_195),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_264),
.B(n_239),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_221),
.B(n_211),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_247),
.B1(n_242),
.B2(n_202),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_233),
.A2(n_208),
.B(n_190),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_279),
.B(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_193),
.B1(n_224),
.B2(n_246),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_283),
.B1(n_258),
.B2(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_256),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_281),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_240),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_242),
.B1(n_244),
.B2(n_226),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_258),
.B1(n_255),
.B2(n_253),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_9),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_267),
.Y(n_290)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_268),
.B1(n_264),
.B2(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_248),
.C(n_261),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_298),
.C(n_270),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_249),
.B(n_205),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_9),
.B(n_14),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_280),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_252),
.C(n_194),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_309),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_281),
.C(n_284),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_308),
.C(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_300),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_9),
.C(n_13),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_7),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_7),
.C(n_13),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_312),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_7),
.C(n_12),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_295),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_315),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_294),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_301),
.B(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_289),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_325),
.B(n_326),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_299),
.B(n_304),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_6),
.B(n_11),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_320),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_10),
.B1(n_11),
.B2(n_16),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_322),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_322),
.C(n_314),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_323),
.B(n_16),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_333),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_331),
.Y(n_336)
);

OAI311xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_335),
.A3(n_330),
.B1(n_16),
.C1(n_5),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_0),
.B(n_3),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_3),
.B(n_4),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_4),
.C(n_5),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_5),
.Y(n_342)
);


endmodule