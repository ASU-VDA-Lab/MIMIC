module fake_netlist_6_820_n_1258 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1258);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1258;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_809;
wire n_220;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_41),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_47),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_94),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_89),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_71),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_28),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_114),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_77),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_27),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_28),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_87),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_14),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_107),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_127),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_105),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_97),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_22),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_78),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_120),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_96),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_42),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_148),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_57),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_2),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_122),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_79),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_149),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_130),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_117),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_211),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_188),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_189),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_190),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_193),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_196),
.Y(n_254)
);

BUFx2_ASAP7_75t_SL g255 ( 
.A(n_218),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_199),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_202),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_204),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_206),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_205),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_236),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_217),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_225),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_179),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_214),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_244),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_251),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_253),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_254),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_259),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_260),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_263),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_263),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_239),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_264),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_257),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_243),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_255),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_255),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_257),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_267),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_267),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_318),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_315),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_315),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_317),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_317),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_275),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_312),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_273),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_279),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_280),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_276),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_316),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_290),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_316),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_282),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_284),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_293),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_288),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_293),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_314),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_273),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_287),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_299),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_291),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

NOR2x1_ASAP7_75t_L g375 ( 
.A(n_321),
.B(n_291),
.Y(n_375)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

BUFx8_ASAP7_75t_SL g377 ( 
.A(n_335),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_332),
.B(n_296),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_270),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_194),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_286),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_197),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_324),
.B(n_287),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_292),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_297),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_349),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_298),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_325),
.B(n_203),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_327),
.B(n_286),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_286),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_319),
.B(n_298),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

BUFx12f_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_286),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_340),
.B(n_207),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_342),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_345),
.Y(n_406)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_319),
.B(n_299),
.Y(n_409)
);

BUFx8_ASAP7_75t_SL g410 ( 
.A(n_362),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_322),
.B(n_301),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g415 ( 
.A1(n_403),
.A2(n_363),
.B(n_348),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_395),
.A2(n_351),
.B(n_350),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_346),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_410),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_369),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_371),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_382),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g426 ( 
.A(n_385),
.B(n_219),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_396),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_382),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_383),
.Y(n_432)
);

BUFx8_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_401),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_398),
.B(n_401),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_322),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_389),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_413),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_398),
.B(n_401),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_387),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_390),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

OAI22x1_ASAP7_75t_L g446 ( 
.A1(n_412),
.A2(n_367),
.B1(n_366),
.B2(n_343),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_398),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g453 ( 
.A(n_385),
.B(n_198),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_370),
.B(n_352),
.Y(n_455)
);

BUFx12f_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_397),
.A2(n_313),
.B(n_310),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_384),
.A2(n_368),
.B1(n_329),
.B2(n_330),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_379),
.B(n_329),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_330),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_375),
.B(n_212),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_380),
.B(n_301),
.Y(n_469)
);

CKINVDCx6p67_ASAP7_75t_R g470 ( 
.A(n_402),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_379),
.A2(n_231),
.B(n_313),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_410),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

AND2x2_ASAP7_75t_SL g474 ( 
.A(n_394),
.B(n_198),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_404),
.B(n_342),
.Y(n_476)
);

CKINVDCx6p67_ASAP7_75t_R g477 ( 
.A(n_386),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_377),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_366),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_201),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_399),
.B(n_367),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_377),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

OAI22x1_ASAP7_75t_SL g485 ( 
.A1(n_391),
.A2(n_339),
.B1(n_358),
.B2(n_357),
.Y(n_485)
);

AND2x2_ASAP7_75t_SL g486 ( 
.A(n_391),
.B(n_198),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

OA21x2_ASAP7_75t_L g488 ( 
.A1(n_407),
.A2(n_308),
.B(n_195),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_407),
.B(n_302),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

BUFx8_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

OR2x2_ASAP7_75t_SL g493 ( 
.A(n_391),
.B(n_343),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_411),
.A2(n_209),
.B(n_208),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_392),
.B(n_357),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_392),
.B(n_358),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_392),
.B(n_364),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_364),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_434),
.B(n_392),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_473),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_428),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_432),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_443),
.B(n_302),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_469),
.B(n_422),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_420),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_483),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_306),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_480),
.B(n_306),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_483),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_420),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_433),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_482),
.B(n_185),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_423),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_R g530 ( 
.A(n_489),
.B(n_180),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_427),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_433),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_425),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_442),
.B(n_374),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_456),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_464),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_447),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_456),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_495),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_422),
.B(n_198),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_441),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_442),
.B(n_374),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_470),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_419),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_470),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_482),
.B(n_438),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_472),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_419),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_419),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_466),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_464),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_459),
.B(n_462),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_472),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_485),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_526),
.B(n_496),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_499),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_519),
.B(n_496),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_524),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_524),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_529),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_529),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_545),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_462),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_557),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_512),
.B(n_497),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_551),
.B(n_497),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_501),
.B(n_495),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_509),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_516),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_426),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_527),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_557),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_505),
.Y(n_582)
);

NOR2x1p5_ASAP7_75t_L g583 ( 
.A(n_539),
.B(n_477),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_531),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_556),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_548),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_532),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_549),
.B(n_426),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_498),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_553),
.B(n_438),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_554),
.B(n_442),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_535),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_500),
.B(n_478),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_507),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_538),
.Y(n_598)
);

INVx8_ASAP7_75t_L g599 ( 
.A(n_535),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_540),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_597),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_583),
.B(n_539),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_599),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_571),
.B(n_477),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_582),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_591),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_587),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_587),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_515),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_591),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_562),
.B(n_495),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_579),
.B(n_504),
.Y(n_612)
);

BUFx6f_ASAP7_75t_SL g613 ( 
.A(n_582),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_599),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_597),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_599),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_595),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_598),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_574),
.B(n_544),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_599),
.B(n_436),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_599),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_582),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_575),
.B(n_436),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_564),
.B(n_528),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_600),
.B(n_596),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_594),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_596),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_590),
.B(n_481),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_594),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_598),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_577),
.B(n_556),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_592),
.A2(n_446),
.B1(n_475),
.B2(n_478),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_577),
.A2(n_446),
.B1(n_463),
.B2(n_468),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_594),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_573),
.A2(n_476),
.B1(n_460),
.B2(n_465),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_595),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_594),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_593),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_577),
.B(n_530),
.Y(n_639)
);

AO21x2_ASAP7_75t_L g640 ( 
.A1(n_576),
.A2(n_418),
.B(n_471),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_600),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_600),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_577),
.B(n_513),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_563),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_563),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_582),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_582),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_593),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_576),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_593),
.B(n_444),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_566),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_593),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_570),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_578),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_580),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_584),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_565),
.B(n_513),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_589),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_589),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_572),
.B(n_555),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_565),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_567),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_570),
.B(n_508),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_567),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_568),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_572),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_585),
.A2(n_467),
.B1(n_525),
.B2(n_503),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_568),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_585),
.B(n_476),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_586),
.B(n_537),
.Y(n_674)
);

OAI21xp33_ASAP7_75t_SL g675 ( 
.A1(n_569),
.A2(n_453),
.B(n_474),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_581),
.B(n_449),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_581),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_586),
.B(n_476),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_588),
.B(n_489),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_569),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_581),
.B(n_546),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_588),
.A2(n_453),
.B1(n_474),
.B2(n_486),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_588),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

AND2x6_ASAP7_75t_L g685 ( 
.A(n_577),
.B(n_513),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_579),
.B(n_449),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_601),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_606),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_610),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_635),
.B(n_517),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_627),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_649),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_653),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_514),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_656),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_624),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_657),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_659),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_661),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_662),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_658),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_617),
.B(n_560),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_636),
.B(n_467),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_658),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_625),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_617),
.B(n_467),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_679),
.B(n_521),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_667),
.B(n_455),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_625),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_622),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_641),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_631),
.B(n_455),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_642),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_664),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_628),
.B(n_521),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_615),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_675),
.A2(n_502),
.B(n_439),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_618),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_631),
.B(n_455),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_612),
.B(n_559),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_630),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_684),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_668),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_675),
.A2(n_502),
.B(n_486),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_686),
.B(n_517),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_669),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_674),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_672),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_635),
.A2(n_471),
.B(n_418),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_648),
.B(n_517),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_644),
.Y(n_731)
);

XNOR2xp5_ASAP7_75t_L g732 ( 
.A(n_609),
.B(n_515),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_612),
.B(n_559),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_645),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_651),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_R g736 ( 
.A(n_629),
.B(n_547),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_605),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_665),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_666),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_666),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_622),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_670),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_670),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_648),
.B(n_523),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_677),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_680),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_682),
.B(n_547),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_632),
.A2(n_458),
.B(n_494),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_677),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_663),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_663),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_655),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_683),
.Y(n_754)
);

INVx3_ASAP7_75t_R g755 ( 
.A(n_608),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_683),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_647),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_611),
.B(n_520),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_683),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_676),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_686),
.B(n_523),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_676),
.Y(n_762)
);

INVxp33_ASAP7_75t_L g763 ( 
.A(n_607),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_673),
.B(n_520),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_639),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_619),
.Y(n_766)
);

INVxp33_ASAP7_75t_L g767 ( 
.A(n_678),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_619),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_602),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_622),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_640),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_681),
.B(n_542),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_640),
.Y(n_773)
);

OR2x2_ASAP7_75t_SL g774 ( 
.A(n_753),
.B(n_633),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_766),
.B(n_632),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_768),
.B(n_652),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_715),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_696),
.B(n_720),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_733),
.B(n_552),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_688),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_736),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_727),
.B(n_652),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_726),
.B(n_623),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_767),
.B(n_603),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_689),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_694),
.B(n_603),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_707),
.B(n_552),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_771),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_763),
.B(n_561),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_701),
.B(n_623),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_704),
.B(n_705),
.Y(n_791)
);

NOR3xp33_ASAP7_75t_L g792 ( 
.A(n_758),
.B(n_682),
.C(n_461),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_709),
.B(n_623),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_691),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_751),
.B(n_671),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_692),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_765),
.B(n_614),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_772),
.B(n_614),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_693),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_752),
.B(n_681),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_710),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_695),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_730),
.B(n_616),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_697),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_698),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_749),
.B(n_621),
.C(n_616),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_730),
.B(n_621),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_699),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_L g809 ( 
.A(n_702),
.B(n_626),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_725),
.B(n_626),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_690),
.B(n_550),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_757),
.B(n_522),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_700),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_725),
.B(n_761),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_710),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_761),
.B(n_634),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_716),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_760),
.B(n_634),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_762),
.B(n_637),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_718),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_721),
.B(n_637),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_745),
.B(n_638),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_748),
.A2(n_769),
.B1(n_602),
.B2(n_724),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_714),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_749),
.B(n_479),
.C(n_523),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_732),
.B(n_522),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_711),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_722),
.B(n_650),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_723),
.B(n_650),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_713),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_728),
.B(n_602),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_687),
.B(n_731),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_734),
.B(n_650),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_735),
.B(n_638),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_738),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_764),
.B(n_533),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_739),
.B(n_646),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_748),
.A2(n_533),
.B1(n_620),
.B2(n_541),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_706),
.B(n_184),
.C(n_179),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_740),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_754),
.B(n_620),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_710),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_770),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_741),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_745),
.B(n_605),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_703),
.B(n_708),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_712),
.A2(n_229),
.B1(n_232),
.B2(n_184),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_737),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_814),
.B(n_773),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_780),
.Y(n_850)
);

NAND3xp33_ASAP7_75t_SL g851 ( 
.A(n_825),
.B(n_724),
.C(n_719),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_824),
.B(n_743),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_777),
.B(n_809),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_824),
.B(n_744),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_785),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_810),
.B(n_747),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_841),
.B(n_717),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_825),
.A2(n_232),
.B(n_233),
.C(n_229),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_794),
.B(n_756),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_804),
.B(n_759),
.Y(n_860)
);

AND2x2_ASAP7_75t_SL g861 ( 
.A(n_811),
.B(n_737),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_816),
.B(n_746),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_778),
.B(n_755),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_775),
.B(n_750),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_796),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_781),
.B(n_770),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_823),
.B(n_770),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_792),
.A2(n_823),
.B1(n_806),
.B2(n_839),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_790),
.B(n_690),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_837),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_841),
.B(n_742),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_795),
.B(n_742),
.C(n_729),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_838),
.A2(n_493),
.B1(n_620),
.B2(n_605),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_SL g874 ( 
.A1(n_774),
.A2(n_836),
.B1(n_779),
.B2(n_787),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_799),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_793),
.B(n_690),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_817),
.B(n_690),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_820),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_831),
.B(n_729),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_835),
.B(n_660),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_801),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_786),
.B(n_493),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_791),
.B(n_660),
.Y(n_883)
);

NOR2x1p5_ASAP7_75t_L g884 ( 
.A(n_783),
.B(n_536),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_782),
.B(n_660),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_788),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_792),
.A2(n_685),
.B1(n_643),
.B2(n_542),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_829),
.B(n_828),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_801),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_848),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_802),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_833),
.B(n_646),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_818),
.B(n_660),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_805),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_819),
.B(n_643),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_808),
.B(n_643),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_848),
.B(n_536),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_813),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_827),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_776),
.B(n_643),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_830),
.B(n_800),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_806),
.A2(n_847),
.B(n_784),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_840),
.B(n_685),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_R g904 ( 
.A(n_812),
.B(n_541),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_834),
.B(n_646),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_844),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_832),
.B(n_821),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_822),
.B(n_479),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_801),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_788),
.Y(n_910)
);

AND2x6_ASAP7_75t_SL g911 ( 
.A(n_789),
.B(n_826),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_846),
.B(n_798),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_815),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_803),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_797),
.A2(n_685),
.B1(n_542),
.B2(n_613),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_807),
.A2(n_847),
.B1(n_845),
.B2(n_685),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_842),
.A2(n_434),
.B(n_451),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_843),
.B(n_0),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_814),
.B(n_0),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_814),
.B(n_1),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_841),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_825),
.A2(n_435),
.B1(n_448),
.B2(n_445),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_823),
.A2(n_613),
.B1(n_494),
.B2(n_234),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_814),
.B(n_1),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_814),
.B(n_2),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_780),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_814),
.B(n_3),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_801),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_890),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_858),
.A2(n_434),
.B(n_451),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_928),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_874),
.A2(n_235),
.B1(n_234),
.B2(n_233),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_SL g933 ( 
.A(n_868),
.B(n_235),
.C(n_215),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_891),
.Y(n_934)
);

INVx5_ASAP7_75t_L g935 ( 
.A(n_857),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_850),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_861),
.B(n_435),
.Y(n_937)
);

OR2x6_ASAP7_75t_L g938 ( 
.A(n_857),
.B(n_505),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_928),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_894),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_910),
.B(n_3),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_921),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_855),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_898),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_909),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_853),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_899),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_924),
.B(n_5),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_890),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_865),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_875),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_914),
.B(n_505),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_886),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_926),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_906),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_849),
.B(n_5),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_871),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_897),
.A2(n_494),
.B(n_488),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_873),
.A2(n_543),
.B1(n_488),
.B2(n_437),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_902),
.B(n_435),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_852),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_888),
.B(n_505),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_851),
.A2(n_434),
.B(n_451),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_849),
.B(n_6),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_857),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_878),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_907),
.B(n_6),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_913),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_852),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_859),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_860),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_888),
.B(n_7),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_881),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_889),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_854),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_856),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_901),
.B(n_7),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_854),
.B(n_8),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_918),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_862),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_867),
.B(n_510),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_911),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_870),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_864),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_903),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_888),
.B(n_9),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_863),
.B(n_9),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_933),
.A2(n_902),
.B(n_925),
.C(n_924),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_984),
.B(n_872),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_933),
.A2(n_873),
.B(n_908),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_982),
.A2(n_923),
.B(n_912),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_960),
.A2(n_866),
.B(n_869),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_982),
.B(n_904),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_954),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_980),
.B(n_879),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_931),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_954),
.Y(n_997)
);

NOR2x1p5_ASAP7_75t_SL g998 ( 
.A(n_975),
.B(n_879),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_935),
.B(n_892),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_963),
.A2(n_876),
.B(n_882),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_963),
.A2(n_925),
.B(n_927),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_976),
.B(n_877),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_953),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_930),
.A2(n_937),
.B(n_932),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_932),
.A2(n_920),
.B(n_919),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_SL g1006 ( 
.A(n_939),
.B(n_883),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_945),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_948),
.A2(n_905),
.B(n_896),
.C(n_895),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_969),
.B(n_893),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_930),
.A2(n_887),
.B(n_917),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_969),
.B(n_900),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_979),
.B(n_885),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_981),
.A2(n_916),
.B1(n_915),
.B2(n_922),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_948),
.A2(n_964),
.B(n_956),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_956),
.A2(n_880),
.B(n_884),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_950),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_983),
.B(n_10),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_941),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_987),
.A2(n_10),
.B(n_11),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_964),
.A2(n_488),
.B(n_216),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_961),
.B(n_11),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_978),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_961),
.B(n_934),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_967),
.A2(n_220),
.B(n_213),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_941),
.A2(n_415),
.B(n_457),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_985),
.B(n_12),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_972),
.A2(n_221),
.B(n_222),
.C(n_223),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_945),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_953),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_979),
.B(n_13),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_986),
.A2(n_224),
.B(n_226),
.C(n_228),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_L g1032 ( 
.A(n_967),
.B(n_490),
.C(n_15),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_936),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_981),
.A2(n_510),
.B1(n_511),
.B2(n_534),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_935),
.B(n_491),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_978),
.A2(n_415),
.B(n_435),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_945),
.Y(n_1037)
);

AND3x2_ASAP7_75t_L g1038 ( 
.A(n_942),
.B(n_15),
.C(n_16),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_985),
.B(n_16),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_977),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_977),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_985),
.B(n_943),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_979),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_959),
.A2(n_534),
.B1(n_511),
.B2(n_510),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_938),
.A2(n_415),
.B(n_437),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_935),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_946),
.B(n_20),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_938),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_951),
.B(n_23),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_966),
.B(n_24),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_935),
.B(n_25),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_929),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_965),
.A2(n_938),
.B(n_955),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_940),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_1007),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1016),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1033),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_996),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_994),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_1007),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_997),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1003),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1029),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1043),
.B(n_965),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1032),
.A2(n_990),
.B1(n_991),
.B2(n_1046),
.Y(n_1065)
);

AND2x6_ASAP7_75t_L g1066 ( 
.A(n_1051),
.B(n_962),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_996),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1022),
.A2(n_965),
.B(n_962),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_1007),
.Y(n_1069)
);

OA21x2_ASAP7_75t_L g1070 ( 
.A1(n_1053),
.A2(n_947),
.B(n_944),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1054),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1043),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1070),
.A2(n_1052),
.B(n_1037),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_1067),
.B(n_996),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_SL g1075 ( 
.A1(n_1064),
.A2(n_1051),
.B(n_1021),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_SL g1076 ( 
.A(n_1064),
.B(n_993),
.Y(n_1076)
);

OAI22x1_ASAP7_75t_L g1077 ( 
.A1(n_1065),
.A2(n_1018),
.B1(n_1047),
.B2(n_1028),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1065),
.B(n_1014),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1058),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1062),
.B(n_1063),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1068),
.B(n_1001),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_1072),
.A2(n_989),
.B(n_1004),
.C(n_1000),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_SL g1083 ( 
.A1(n_1067),
.A2(n_1040),
.B(n_1041),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1072),
.B(n_999),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_L g1085 ( 
.A1(n_1059),
.A2(n_1010),
.B(n_999),
.C(n_1019),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1069),
.A2(n_988),
.B(n_1024),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1069),
.A2(n_1005),
.B(n_1048),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1062),
.B(n_1023),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1063),
.B(n_1049),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1056),
.B(n_1011),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1055),
.B(n_995),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1055),
.B(n_1012),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1070),
.A2(n_1015),
.B(n_1020),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1055),
.A2(n_998),
.B(n_1030),
.C(n_992),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1070),
.A2(n_1017),
.B(n_1027),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1066),
.A2(n_1036),
.B(n_1031),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1060),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_1097),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_L g1099 ( 
.A(n_1078),
.B(n_1066),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1084),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1080),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1080),
.Y(n_1102)
);

AO21x2_ASAP7_75t_L g1103 ( 
.A1(n_1093),
.A2(n_1061),
.B(n_1059),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1076),
.B(n_1060),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1100),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1103),
.A2(n_1083),
.B(n_1081),
.Y(n_1106)
);

BUFx2_ASAP7_75t_R g1107 ( 
.A(n_1105),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1106),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1107),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1108),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1110),
.Y(n_1111)
);

INVxp33_ASAP7_75t_L g1112 ( 
.A(n_1109),
.Y(n_1112)
);

OA21x2_ASAP7_75t_L g1113 ( 
.A1(n_1111),
.A2(n_1082),
.B(n_1104),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1112),
.B(n_1079),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1112),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_1101),
.Y(n_1116)
);

AOI222xp33_ASAP7_75t_L g1117 ( 
.A1(n_1115),
.A2(n_1099),
.B1(n_1077),
.B2(n_1102),
.C1(n_1104),
.C2(n_1100),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1113),
.B(n_1100),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1118),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1116),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1120),
.B(n_1100),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1119),
.A2(n_1103),
.B1(n_1098),
.B2(n_1099),
.C(n_1087),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1121),
.B(n_1113),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1122),
.B(n_1117),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1124),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1126),
.A2(n_1098),
.B1(n_1089),
.B2(n_1084),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1125),
.B(n_1098),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1128),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1127),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1129),
.B(n_1098),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1130),
.B(n_1103),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1129),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_1132),
.B(n_25),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1133),
.B(n_1060),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1131),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1135),
.Y(n_1137)
);

AND2x2_ASAP7_75t_SL g1138 ( 
.A(n_1136),
.B(n_1089),
.Y(n_1138)
);

XOR2x2_ASAP7_75t_L g1139 ( 
.A(n_1138),
.B(n_1134),
.Y(n_1139)
);

XOR2x2_ASAP7_75t_L g1140 ( 
.A(n_1137),
.B(n_1038),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1140),
.B(n_1139),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1140),
.B(n_1086),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1142),
.B(n_1074),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1141),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1143),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1144),
.B(n_1092),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1146),
.Y(n_1147)
);

CKINVDCx16_ASAP7_75t_R g1148 ( 
.A(n_1145),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1147),
.Y(n_1149)
);

OAI322xp33_ASAP7_75t_L g1150 ( 
.A1(n_1148),
.A2(n_1095),
.A3(n_1088),
.B1(n_30),
.B2(n_31),
.C1(n_26),
.C2(n_29),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1147),
.B(n_1073),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_SL g1152 ( 
.A(n_1149),
.B(n_1085),
.C(n_1094),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

OAI32xp33_ASAP7_75t_L g1154 ( 
.A1(n_1150),
.A2(n_1088),
.A3(n_1090),
.B1(n_1061),
.B2(n_1026),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1153),
.A2(n_1096),
.B(n_1091),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1152),
.Y(n_1156)
);

AOI222xp33_ASAP7_75t_L g1157 ( 
.A1(n_1156),
.A2(n_1154),
.B1(n_29),
.B2(n_30),
.C1(n_31),
.C2(n_26),
.Y(n_1157)
);

OAI321xp33_ASAP7_75t_L g1158 ( 
.A1(n_1155),
.A2(n_1039),
.A3(n_1050),
.B1(n_1071),
.B2(n_1057),
.C(n_1075),
.Y(n_1158)
);

AND2x4_ASAP7_75t_SL g1159 ( 
.A(n_1157),
.B(n_1056),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1158),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1160),
.B(n_32),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1159),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1161),
.A2(n_316),
.B(n_1057),
.C(n_1071),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1162),
.A2(n_1070),
.B1(n_1066),
.B2(n_491),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1163),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1164),
.A2(n_33),
.B(n_34),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1166),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1165),
.Y(n_1168)
);

OAI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1166),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.C(n_44),
.Y(n_1169)
);

NOR3xp33_ASAP7_75t_SL g1170 ( 
.A(n_1168),
.B(n_45),
.C(n_46),
.Y(n_1170)
);

OAI211xp5_ASAP7_75t_L g1171 ( 
.A1(n_1169),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1171)
);

NAND4xp25_ASAP7_75t_L g1172 ( 
.A(n_1167),
.B(n_51),
.C(n_52),
.D(n_53),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_SL g1173 ( 
.A(n_1172),
.B(n_491),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1171),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_SL g1175 ( 
.A(n_1173),
.B(n_1170),
.C(n_58),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1174),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_1175),
.Y(n_1177)
);

NOR3x1_ASAP7_75t_L g1178 ( 
.A(n_1176),
.B(n_64),
.C(n_65),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1177),
.A2(n_1066),
.B1(n_1035),
.B2(n_68),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1178),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1180),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1179),
.A2(n_1066),
.B1(n_67),
.B2(n_69),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1181),
.B(n_66),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1182),
.Y(n_1184)
);

NOR4xp25_ASAP7_75t_L g1185 ( 
.A(n_1184),
.B(n_70),
.C(n_72),
.D(n_73),
.Y(n_1185)
);

OAI311xp33_ASAP7_75t_L g1186 ( 
.A1(n_1183),
.A2(n_74),
.A3(n_75),
.B1(n_76),
.C1(n_81),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1184),
.B(n_82),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1186),
.A2(n_83),
.B(n_84),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1185),
.A2(n_1187),
.B1(n_88),
.B2(n_90),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1185),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1190),
.Y(n_1191)
);

NOR4xp25_ASAP7_75t_L g1192 ( 
.A(n_1189),
.B(n_85),
.C(n_91),
.D(n_92),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1191),
.B(n_1188),
.Y(n_1193)
);

OR2x2_ASAP7_75t_SL g1194 ( 
.A(n_1192),
.B(n_93),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_1193),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1194),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1195),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1196),
.Y(n_1198)
);

NOR2x1_ASAP7_75t_L g1199 ( 
.A(n_1198),
.B(n_103),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1197),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1200),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1199),
.B(n_104),
.C(n_106),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1201),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1202),
.B(n_108),
.C(n_110),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1201),
.B(n_111),
.C(n_112),
.Y(n_1205)
);

AOI32xp33_ASAP7_75t_L g1206 ( 
.A1(n_1203),
.A2(n_113),
.A3(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_1206)
);

NOR2x1_ASAP7_75t_L g1207 ( 
.A(n_1204),
.B(n_124),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1205),
.Y(n_1208)
);

NAND2x1_ASAP7_75t_L g1209 ( 
.A(n_1208),
.B(n_1066),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1207),
.B(n_125),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1210),
.A2(n_1206),
.B(n_129),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1209),
.A2(n_126),
.B(n_132),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1211),
.B(n_133),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_1212),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_R g1215 ( 
.A(n_1211),
.B(n_138),
.Y(n_1215)
);

AO22x2_ASAP7_75t_SL g1216 ( 
.A1(n_1215),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1213),
.A2(n_1214),
.B1(n_973),
.B2(n_974),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1213),
.A2(n_1066),
.B1(n_152),
.B2(n_153),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1217),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1217),
.A2(n_973),
.B1(n_949),
.B2(n_929),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1219),
.A2(n_973),
.B1(n_949),
.B2(n_437),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1220),
.A2(n_448),
.B1(n_437),
.B2(n_445),
.Y(n_1223)
);

AOI211xp5_ASAP7_75t_L g1224 ( 
.A1(n_1221),
.A2(n_150),
.B(n_155),
.C(n_156),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1219),
.A2(n_534),
.B1(n_511),
.B2(n_510),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1219),
.A2(n_448),
.B1(n_445),
.B2(n_1052),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1219),
.A2(n_448),
.B1(n_445),
.B2(n_534),
.Y(n_1227)
);

AOI211xp5_ASAP7_75t_L g1228 ( 
.A1(n_1219),
.A2(n_157),
.B(n_158),
.C(n_159),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1219),
.A2(n_511),
.B1(n_546),
.B2(n_416),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1219),
.A2(n_546),
.B1(n_429),
.B2(n_416),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1219),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1219),
.A2(n_429),
.B1(n_416),
.B2(n_168),
.Y(n_1232)
);

OAI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1219),
.A2(n_164),
.B1(n_167),
.B2(n_169),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1219),
.A2(n_172),
.B(n_173),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1234),
.A2(n_174),
.B(n_175),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1224),
.A2(n_176),
.B(n_177),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1231),
.A2(n_178),
.B(n_958),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1232),
.A2(n_1034),
.B(n_968),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1222),
.B(n_416),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1233),
.A2(n_429),
.B(n_425),
.C(n_431),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1225),
.B(n_1229),
.Y(n_1241)
);

AOI22x1_ASAP7_75t_L g1242 ( 
.A1(n_1226),
.A2(n_429),
.B1(n_431),
.B2(n_492),
.Y(n_1242)
);

XOR2xp5_ASAP7_75t_L g1243 ( 
.A(n_1230),
.B(n_1013),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1241),
.A2(n_1227),
.B(n_1223),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1239),
.A2(n_1240),
.B(n_1237),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1235),
.A2(n_1228),
.B(n_487),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1242),
.B(n_374),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1236),
.B(n_376),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1243),
.B(n_376),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1245),
.A2(n_1238),
.B1(n_952),
.B2(n_1042),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1244),
.A2(n_431),
.B1(n_952),
.B2(n_543),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1249),
.A2(n_543),
.B1(n_431),
.B2(n_1044),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1250),
.B(n_1246),
.Y(n_1253)
);

AOI221xp5_ASAP7_75t_L g1254 ( 
.A1(n_1253),
.A2(n_1248),
.B1(n_1247),
.B2(n_1251),
.C(n_1252),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1254),
.A2(n_1008),
.B(n_1006),
.Y(n_1255)
);

AOI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1255),
.A2(n_965),
.B(n_957),
.Y(n_1256)
);

AOI211xp5_ASAP7_75t_L g1257 ( 
.A1(n_1256),
.A2(n_1045),
.B(n_1009),
.C(n_1002),
.Y(n_1257)
);

AOI211xp5_ASAP7_75t_L g1258 ( 
.A1(n_1257),
.A2(n_971),
.B(n_970),
.C(n_1025),
.Y(n_1258)
);


endmodule