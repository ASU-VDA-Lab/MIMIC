module fake_jpeg_4876_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_17),
.B1(n_22),
.B2(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_32),
.B1(n_16),
.B2(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_50),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_51),
.B1(n_40),
.B2(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_50),
.C(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_70),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_40),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_39),
.C(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_64),
.C(n_71),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_20),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_56),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_77),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_39),
.C(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_61),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_89),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_67),
.B(n_70),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_79),
.B1(n_75),
.B2(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_88),
.B1(n_89),
.B2(n_94),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_102),
.B(n_34),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_76),
.C(n_74),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_104),
.C(n_102),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_39),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_44),
.C(n_35),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_88),
.B1(n_84),
.B2(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

AOI321xp33_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_114),
.A3(n_112),
.B1(n_24),
.B2(n_23),
.C(n_9),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_72),
.B1(n_37),
.B2(n_20),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_69),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_113),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_44),
.C(n_19),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_0),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_44),
.C(n_24),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_98),
.B(n_100),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_118),
.B(n_116),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_9),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_124),
.B(n_7),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_7),
.B(n_1),
.C(n_3),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_3),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_0),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_4),
.B(n_5),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_133),
.A2(n_6),
.B(n_23),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_5),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_132),
.Y(n_137)
);


endmodule