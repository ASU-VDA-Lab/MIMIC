module fake_jpeg_1383_n_54 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_54);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_10),
.Y(n_20)
);

CKINVDCx9p33_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_25),
.Y(n_26)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_20),
.C(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_19),
.B1(n_16),
.B2(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_25),
.B1(n_19),
.B2(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_20),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_31),
.B1(n_5),
.B2(n_6),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_34),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_8),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_37),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_4),
.B1(n_12),
.B2(n_13),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_14),
.B(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_48),
.C(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_50),
.C(n_42),
.Y(n_54)
);


endmodule