module fake_aes_7833_n_15 (n_3, n_1, n_2, n_0, n_15);
input n_3;
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
BUFx10_ASAP7_75t_L g4 ( .A(n_3), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_1), .Y(n_5) );
NOR2xp33_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_5), .B(n_2), .Y(n_7) );
NOR2xp33_ASAP7_75t_L g8 ( .A(n_7), .B(n_4), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
OR2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
BUFx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
BUFx2_ASAP7_75t_SL g15 ( .A(n_14), .Y(n_15) );
endmodule