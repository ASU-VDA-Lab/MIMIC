module fake_aes_12223_n_658 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_658);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_658;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_66), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_24), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_27), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_49), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_14), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_8), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_59), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_34), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_64), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_58), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_9), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_17), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_13), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_42), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_37), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_77), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_16), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_65), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_30), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_4), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_4), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_46), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_17), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_72), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_61), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_15), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_74), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_23), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_20), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_10), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_10), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_21), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_26), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_40), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_5), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_2), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_106), .B(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_90), .Y(n_124) );
NOR2x1_ASAP7_75t_L g125 ( .A(n_90), .B(n_0), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_106), .B(n_1), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_115), .B(n_1), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
XOR2xp5_ASAP7_75t_L g130 ( .A(n_97), .B(n_2), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_94), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_98), .B(n_3), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_92), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_94), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_101), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_115), .B(n_5), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_78), .Y(n_139) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_81), .A2(n_39), .B(n_75), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_81), .Y(n_142) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_92), .A2(n_38), .B(n_73), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_83), .B(n_6), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_112), .B(n_6), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_78), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_112), .B(n_7), .Y(n_147) );
BUFx12f_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
NOR2xp67_ASAP7_75t_L g150 ( .A(n_85), .B(n_7), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_94), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_85), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_79), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_86), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_86), .Y(n_156) );
NAND2xp33_ASAP7_75t_L g157 ( .A(n_94), .B(n_41), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_94), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_132), .B(n_107), .Y(n_162) );
XOR2x2_ASAP7_75t_SL g163 ( .A(n_122), .B(n_83), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_122), .B(n_113), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_128), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_138), .B(n_82), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_138), .B(n_82), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_141), .B(n_121), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_122), .B(n_99), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_122), .A2(n_104), .B1(n_111), .B2(n_91), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_122), .B(n_88), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_132), .B(n_105), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_138), .A2(n_120), .B1(n_108), .B2(n_91), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_141), .B(n_119), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_137), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_127), .B(n_102), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_154), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_127), .B(n_102), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_128), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_126), .B(n_88), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_126), .B(n_114), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_133), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_141), .B(n_119), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_134), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_141), .B(n_118), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_141), .B(n_118), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_163), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_167), .B(n_126), .Y(n_206) );
AND3x2_ASAP7_75t_SL g207 ( .A(n_163), .B(n_130), .C(n_183), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_167), .B(n_126), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_161), .Y(n_211) );
INVxp67_ASAP7_75t_L g212 ( .A(n_185), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_161), .B(n_198), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_161), .B(n_126), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_174), .Y(n_216) );
OR2x6_ASAP7_75t_L g217 ( .A(n_198), .B(n_132), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_198), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_186), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_173), .B(n_148), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_198), .B(n_176), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_168), .B(n_129), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_178), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_178), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_168), .B(n_129), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_184), .B(n_135), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_179), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_162), .A2(n_145), .B1(n_147), .B2(n_155), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_191), .B(n_145), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_179), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_188), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_162), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_184), .B(n_130), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_187), .B(n_135), .Y(n_238) );
BUFx4f_ASAP7_75t_L g239 ( .A(n_162), .Y(n_239) );
INVx5_ASAP7_75t_L g240 ( .A(n_162), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_188), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_187), .B(n_142), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_162), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_191), .B(n_142), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_190), .B(n_155), .Y(n_245) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_176), .B(n_145), .Y(n_246) );
INVx4_ASAP7_75t_L g247 ( .A(n_162), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_190), .B(n_152), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_177), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_162), .B(n_152), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_192), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_177), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_180), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_177), .B(n_145), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_249), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_220), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_229), .B(n_175), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_209), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_247), .B(n_177), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_240), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_238), .B(n_180), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_220), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_247), .B(n_176), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_215), .A2(n_164), .B(n_172), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_253), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_206), .A2(n_144), .B(n_201), .C(n_182), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_242), .B(n_224), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_247), .B(n_193), .Y(n_269) );
BUFx12f_ASAP7_75t_L g270 ( .A(n_219), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_209), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_251), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_208), .A2(n_199), .B(n_192), .C(n_195), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_255), .A2(n_180), .B1(n_147), .B2(n_152), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_222), .B(n_181), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_251), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_240), .B(n_181), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_215), .A2(n_166), .B(n_169), .Y(n_279) );
OR2x6_ASAP7_75t_L g280 ( .A(n_220), .B(n_148), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_205), .A2(n_180), .B1(n_137), .B2(n_148), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_255), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_232), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_SL g285 ( .A1(n_250), .A2(n_202), .B(n_196), .C(n_110), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_212), .B(n_130), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_255), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_219), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_235), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_244), .A2(n_144), .B(n_199), .C(n_195), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_231), .A2(n_147), .B1(n_180), .B2(n_152), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_235), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_228), .B(n_180), .Y(n_293) );
NOR3xp33_ASAP7_75t_L g294 ( .A(n_227), .B(n_125), .C(n_114), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_211), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_211), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_222), .B(n_180), .Y(n_297) );
AOI22xp33_ASAP7_75t_SL g298 ( .A1(n_205), .A2(n_147), .B1(n_180), .B2(n_116), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_245), .A2(n_147), .B(n_156), .C(n_152), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_217), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_239), .A2(n_156), .B1(n_150), .B2(n_166), .Y(n_301) );
NAND2x1_ASAP7_75t_L g302 ( .A(n_217), .B(n_124), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_289), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_268), .B(n_233), .Y(n_304) );
OAI211xp5_ASAP7_75t_L g305 ( .A1(n_298), .A2(n_150), .B(n_237), .C(n_125), .Y(n_305) );
AOI21xp33_ASAP7_75t_SL g306 ( .A1(n_288), .A2(n_207), .B(n_246), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_286), .B(n_248), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_290), .A2(n_143), .B(n_140), .Y(n_308) );
AO31x2_ASAP7_75t_L g309 ( .A1(n_273), .A2(n_134), .A3(n_158), .B(n_153), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_256), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_301), .A2(n_143), .B(n_140), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_273), .A2(n_143), .B(n_216), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_262), .A2(n_221), .B(n_203), .Y(n_314) );
OAI22xp33_ASAP7_75t_SL g315 ( .A1(n_281), .A2(n_207), .B1(n_217), .B2(n_116), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_266), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_299), .A2(n_140), .B(n_246), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_275), .A2(n_217), .B1(n_233), .B2(n_252), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_300), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_259), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_267), .A2(n_233), .B(n_239), .C(n_241), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_265), .A2(n_140), .B(n_156), .Y(n_322) );
INVx5_ASAP7_75t_L g323 ( .A(n_257), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_298), .B(n_241), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_271), .Y(n_325) );
OA21x2_ASAP7_75t_L g326 ( .A1(n_279), .A2(n_105), .B(n_110), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_275), .A2(n_218), .B1(n_223), .B2(n_239), .Y(n_327) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_302), .A2(n_140), .B(n_156), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_291), .A2(n_156), .B(n_252), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_293), .A2(n_204), .B(n_210), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_258), .B(n_213), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_264), .A2(n_225), .B(n_226), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
AO21x2_ASAP7_75t_L g334 ( .A1(n_285), .A2(n_134), .B(n_89), .Y(n_334) );
OAI21x1_ASAP7_75t_L g335 ( .A1(n_264), .A2(n_234), .B(n_230), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_323), .B(n_269), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_313), .A2(n_285), .B(n_297), .Y(n_338) );
AOI21xp5_ASAP7_75t_SL g339 ( .A1(n_321), .A2(n_254), .B(n_280), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g340 ( .A1(n_305), .A2(n_294), .B1(n_284), .B2(n_274), .C(n_297), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g341 ( .A1(n_315), .A2(n_269), .B1(n_270), .B2(n_300), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_306), .A2(n_294), .B1(n_315), .B2(n_305), .C(n_304), .Y(n_342) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_324), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_304), .B(n_278), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g345 ( .A1(n_318), .A2(n_307), .B1(n_306), .B2(n_331), .C(n_327), .Y(n_345) );
AO31x2_ASAP7_75t_L g346 ( .A1(n_310), .A2(n_153), .A3(n_158), .B(n_123), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_318), .A2(n_278), .B1(n_260), .B2(n_283), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_331), .A2(n_287), .B1(n_274), .B2(n_260), .C(n_123), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_311), .A2(n_280), .B1(n_272), .B2(n_277), .C(n_276), .Y(n_350) );
OAI221xp5_ASAP7_75t_SL g351 ( .A1(n_324), .A2(n_280), .B1(n_95), .B2(n_100), .C(n_89), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_311), .A2(n_223), .B1(n_295), .B2(n_124), .C(n_214), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_323), .B(n_254), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_310), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_323), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_316), .B(n_263), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_313), .A2(n_158), .B(n_153), .Y(n_357) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_314), .A2(n_124), .B(n_295), .C(n_128), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_310), .A2(n_254), .B1(n_243), .B2(n_236), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_316), .B(n_263), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_312), .A2(n_95), .B(n_93), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_354), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_354), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_362), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_362), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_361), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_349), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_361), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_355), .B(n_323), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_336), .B(n_303), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_337), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_361), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_343), .B(n_303), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_346), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_344), .B(n_325), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_345), .B(n_319), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_355), .B(n_325), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_340), .A2(n_314), .B1(n_333), .B2(n_320), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_356), .B(n_320), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_341), .B(n_103), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_342), .A2(n_124), .B1(n_100), .B2(n_96), .C(n_93), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_346), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_348), .A2(n_333), .B1(n_334), .B2(n_329), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_356), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_357), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_356), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_360), .B(n_333), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_363), .B(n_309), .Y(n_395) );
OAI31xp33_ASAP7_75t_L g396 ( .A1(n_384), .A2(n_351), .A3(n_350), .B(n_347), .Y(n_396) );
OAI21xp33_ASAP7_75t_L g397 ( .A1(n_374), .A2(n_96), .B(n_109), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_363), .B(n_309), .Y(n_398) );
OAI33xp33_ASAP7_75t_L g399 ( .A1(n_374), .A2(n_109), .A3(n_107), .B1(n_11), .B2(n_12), .B3(n_13), .Y(n_399) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_385), .B(n_358), .C(n_338), .Y(n_400) );
OAI211xp5_ASAP7_75t_SL g401 ( .A1(n_371), .A2(n_87), .B(n_117), .C(n_339), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_364), .B(n_309), .Y(n_402) );
OAI33xp33_ASAP7_75t_L g403 ( .A1(n_378), .A2(n_8), .A3(n_9), .B1(n_11), .B2(n_12), .B3(n_14), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_377), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_364), .B(n_309), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_389), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_368), .B(n_309), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_376), .B(n_360), .Y(n_408) );
AOI33xp33_ASAP7_75t_L g409 ( .A1(n_376), .A2(n_360), .A3(n_352), .B1(n_19), .B2(n_16), .B3(n_18), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_365), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_368), .B(n_381), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_386), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_365), .B(n_309), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_366), .B(n_357), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_387), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_367), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_387), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_366), .B(n_326), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_372), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_378), .A2(n_358), .B1(n_339), .B2(n_353), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_375), .B(n_326), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_367), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_369), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_369), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_380), .A2(n_329), .B1(n_334), .B2(n_330), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_372), .A2(n_124), .B(n_326), .C(n_353), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_382), .B(n_326), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_375), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g432 ( .A1(n_372), .A2(n_317), .B(n_136), .C(n_151), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_382), .B(n_334), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_372), .B(n_334), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_373), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_370), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_403), .A2(n_392), .B1(n_390), .B2(n_393), .C(n_383), .Y(n_437) );
NOR2xp67_ASAP7_75t_L g438 ( .A(n_422), .B(n_373), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_419), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_436), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_395), .B(n_383), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_407), .B(n_389), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_412), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_414), .B(n_390), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_395), .B(n_391), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_391), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_394), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_396), .B(n_392), .C(n_393), .D(n_388), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_415), .B(n_370), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_407), .B(n_370), .Y(n_451) );
OAI322xp33_ASAP7_75t_L g452 ( .A1(n_404), .A2(n_388), .A3(n_136), .B1(n_151), .B2(n_131), .C1(n_18), .C2(n_19), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_404), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_370), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_408), .B(n_330), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_436), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_397), .A2(n_157), .B(n_317), .Y(n_457) );
AND2x4_ASAP7_75t_SL g458 ( .A(n_411), .B(n_257), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_402), .B(n_136), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_410), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_413), .Y(n_462) );
NOR3xp33_ASAP7_75t_SL g463 ( .A(n_399), .B(n_214), .C(n_359), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_413), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_402), .B(n_335), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_397), .A2(n_157), .B1(n_131), .B2(n_151), .C(n_159), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_418), .B(n_131), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_419), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_405), .B(n_131), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_405), .B(n_131), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_420), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_416), .B(n_131), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g476 ( .A(n_436), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_430), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_416), .B(n_151), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_401), .A2(n_335), .B1(n_332), .B2(n_312), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_431), .B(n_426), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_426), .B(n_323), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_427), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_433), .B(n_151), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_433), .B(n_151), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_431), .Y(n_485) );
OAI33xp33_ASAP7_75t_L g486 ( .A1(n_423), .A2(n_197), .A3(n_194), .B1(n_170), .B2(n_159), .B3(n_151), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_427), .B(n_419), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_425), .B(n_151), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_430), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g490 ( .A(n_424), .B(n_323), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_425), .B(n_332), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_409), .B(n_308), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_425), .B(n_308), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_439), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_489), .B(n_421), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_440), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_443), .Y(n_497) );
NOR2xp33_ASAP7_75t_SL g498 ( .A(n_476), .B(n_421), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_489), .B(n_434), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_438), .A2(n_429), .B(n_432), .C(n_400), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_477), .B(n_435), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_481), .B(n_424), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_441), .B(n_435), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_452), .B(n_400), .C(n_428), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_485), .B(n_435), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_490), .Y(n_507) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_481), .B(n_417), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_482), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_441), .B(n_406), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_445), .B(n_406), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_483), .B(n_417), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_451), .B(n_406), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_439), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g516 ( .A(n_449), .B(n_428), .C(n_159), .D(n_170), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_442), .B(n_406), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_481), .B(n_406), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_442), .B(n_406), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_469), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_456), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_445), .B(n_328), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_448), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_460), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_447), .B(n_322), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_460), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_453), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_447), .B(n_328), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_454), .B(n_322), .Y(n_529) );
NOR2xp67_ASAP7_75t_L g530 ( .A(n_480), .B(n_323), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_454), .B(n_483), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_487), .B(n_25), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_484), .B(n_28), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_469), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_461), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_484), .B(n_29), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_463), .A2(n_236), .B(n_240), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_487), .B(n_31), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_444), .B(n_32), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_471), .B(n_33), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_471), .B(n_35), .Y(n_542) );
INVxp33_ASAP7_75t_L g543 ( .A(n_490), .Y(n_543) );
INVxp33_ASAP7_75t_L g544 ( .A(n_490), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_468), .B(n_282), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_472), .B(n_36), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_472), .B(n_43), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_462), .B(n_44), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_474), .B(n_45), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_464), .Y(n_550) );
AOI321xp33_ASAP7_75t_L g551 ( .A1(n_504), .A2(n_450), .A3(n_492), .B1(n_451), .B2(n_437), .C(n_478), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_550), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_530), .B(n_480), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_497), .B(n_478), .C(n_474), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_506), .B(n_466), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_506), .B(n_473), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_496), .B(n_475), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_512), .B(n_470), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_496), .B(n_455), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_500), .A2(n_479), .B(n_468), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_550), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g562 ( .A1(n_516), .A2(n_457), .B1(n_467), .B2(n_493), .C(n_491), .Y(n_562) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_540), .A2(n_488), .B(n_491), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_521), .A2(n_486), .B(n_488), .C(n_170), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_509), .Y(n_565) );
NAND3x2_ASAP7_75t_L g566 ( .A(n_531), .B(n_47), .C(n_48), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_499), .A2(n_458), .B1(n_282), .B2(n_257), .Y(n_567) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_508), .B(n_458), .Y(n_568) );
OAI211xp5_ASAP7_75t_L g569 ( .A1(n_507), .A2(n_261), .B(n_236), .C(n_240), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_513), .B(n_53), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_521), .B(n_55), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_503), .B(n_56), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_503), .B(n_57), .Y(n_573) );
OAI32xp33_ASAP7_75t_L g574 ( .A1(n_543), .A2(n_261), .A3(n_243), .B1(n_63), .B2(n_67), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_531), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_514), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_524), .A2(n_197), .B1(n_194), .B2(n_160), .C(n_200), .Y(n_577) );
INVxp33_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_505), .B(n_197), .C(n_194), .D(n_218), .Y(n_579) );
AOI21xp33_ASAP7_75t_L g580 ( .A1(n_543), .A2(n_60), .B(n_62), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_526), .A2(n_254), .B1(n_160), .B2(n_200), .C(n_257), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_544), .A2(n_282), .B1(n_236), .B2(n_240), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_523), .B(n_68), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_527), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_544), .B(n_70), .Y(n_585) );
AO22x1_ASAP7_75t_L g586 ( .A1(n_495), .A2(n_282), .B1(n_76), .B2(n_71), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_532), .B(n_160), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g588 ( .A1(n_548), .A2(n_166), .B(n_169), .C(n_189), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_536), .Y(n_589) );
BUFx2_ASAP7_75t_SL g590 ( .A(n_533), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_494), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_556), .B(n_510), .Y(n_593) );
INVx2_ASAP7_75t_SL g594 ( .A(n_575), .Y(n_594) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_578), .A2(n_502), .B(n_549), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_559), .B(n_510), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_552), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_561), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_555), .B(n_511), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_592), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_565), .B(n_511), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_591), .Y(n_602) );
AND3x4_ASAP7_75t_L g603 ( .A(n_568), .B(n_533), .C(n_514), .Y(n_603) );
AOI222xp33_ASAP7_75t_L g604 ( .A1(n_560), .A2(n_529), .B1(n_539), .B2(n_522), .C1(n_528), .C2(n_501), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_584), .B(n_529), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_557), .B(n_518), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_589), .B(n_522), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_553), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_572), .B(n_533), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_551), .A2(n_547), .B1(n_546), .B2(n_541), .C(n_519), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_563), .B(n_571), .C(n_576), .D(n_562), .Y(n_612) );
OAI31xp33_ASAP7_75t_L g613 ( .A1(n_579), .A2(n_549), .A3(n_542), .B(n_537), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_558), .B(n_528), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_573), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_587), .Y(n_616) );
INVxp67_ASAP7_75t_L g617 ( .A(n_587), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_580), .B(n_538), .C(n_534), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_611), .A2(n_563), .B1(n_590), .B2(n_570), .C(n_539), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_595), .A2(n_580), .B(n_585), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_617), .B(n_520), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_605), .B(n_519), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_597), .Y(n_623) );
AOI322xp5_ASAP7_75t_L g624 ( .A1(n_611), .A2(n_542), .A3(n_534), .B1(n_537), .B2(n_570), .C1(n_583), .C2(n_567), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_613), .A2(n_588), .B(n_569), .C(n_564), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_612), .A2(n_566), .B(n_581), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_598), .Y(n_627) );
NOR3x1_ASAP7_75t_L g628 ( .A(n_594), .B(n_586), .C(n_517), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_617), .A2(n_574), .B(n_525), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_618), .A2(n_582), .B(n_577), .Y(n_630) );
AOI21xp33_ASAP7_75t_SL g631 ( .A1(n_603), .A2(n_545), .B(n_525), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_604), .A2(n_494), .B(n_535), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_616), .B(n_515), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_621), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_632), .A2(n_608), .B(n_606), .Y(n_635) );
OA211x2_ASAP7_75t_L g636 ( .A1(n_626), .A2(n_603), .B(n_596), .C(n_601), .Y(n_636) );
AOI21xp33_ASAP7_75t_L g637 ( .A1(n_630), .A2(n_625), .B(n_620), .Y(n_637) );
NAND3xp33_ASAP7_75t_SL g638 ( .A(n_631), .B(n_618), .C(n_609), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_628), .B(n_600), .Y(n_639) );
NAND5xp2_ASAP7_75t_L g640 ( .A(n_619), .B(n_610), .C(n_609), .D(n_545), .E(n_607), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_633), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_624), .A2(n_615), .B1(n_600), .B2(n_593), .C(n_614), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_637), .B(n_638), .C(n_642), .Y(n_643) );
OAI222xp33_ASAP7_75t_R g644 ( .A1(n_636), .A2(n_627), .B1(n_623), .B2(n_629), .C1(n_602), .C2(n_622), .Y(n_644) );
AND2x4_ASAP7_75t_SL g645 ( .A(n_639), .B(n_520), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_634), .B(n_599), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_641), .B(n_633), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_646), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_645), .B(n_638), .Y(n_649) );
NAND5xp2_ASAP7_75t_L g650 ( .A(n_643), .B(n_644), .C(n_635), .D(n_640), .E(n_545), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_648), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_649), .A2(n_647), .B1(n_515), .B2(n_535), .Y(n_652) );
OAI22xp5_ASAP7_75t_SL g653 ( .A1(n_651), .A2(n_649), .B1(n_650), .B2(n_189), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_652), .A2(n_160), .B1(n_200), .B2(n_189), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_655), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_654), .B1(n_200), .B2(n_160), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_160), .B1(n_169), .B2(n_200), .C(n_637), .Y(n_658) );
endmodule