module fake_jpeg_12213_n_368 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_368);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_368;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g134 ( 
.A(n_54),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_60),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_61),
.Y(n_110)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_7),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_79),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g138 ( 
.A(n_75),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_78),
.Y(n_140)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_5),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_45),
.B(n_5),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_83),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_23),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_9),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_44),
.Y(n_135)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_95),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_26),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_36),
.B(n_13),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g179 ( 
.A(n_101),
.B(n_102),
.Y(n_179)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_46),
.CON(n_102),
.SN(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_74),
.B1(n_81),
.B2(n_27),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_105),
.A2(n_120),
.B1(n_121),
.B2(n_144),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_18),
.C(n_26),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_108),
.A2(n_117),
.B(n_119),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_26),
.B1(n_38),
.B2(n_31),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_112),
.A2(n_89),
.B(n_95),
.C(n_63),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_56),
.A2(n_24),
.B1(n_36),
.B2(n_38),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_38),
.B1(n_31),
.B2(n_28),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_31),
.B1(n_28),
.B2(n_19),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_65),
.A2(n_24),
.B1(n_28),
.B2(n_19),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_132),
.B1(n_142),
.B2(n_143),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_19),
.B1(n_46),
.B2(n_21),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_141),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_80),
.B(n_1),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_67),
.A2(n_44),
.B1(n_39),
.B2(n_29),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_72),
.A2(n_39),
.B1(n_29),
.B2(n_21),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_96),
.B(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_147),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_77),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_86),
.B1(n_4),
.B2(n_54),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_152),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_138),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_157),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_88),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_54),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_110),
.B1(n_130),
.B2(n_136),
.Y(n_198)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_174),
.B1(n_188),
.B2(n_190),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_10),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_10),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_187),
.Y(n_195)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_117),
.A2(n_95),
.A3(n_63),
.B1(n_12),
.B2(n_48),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_134),
.C(n_127),
.Y(n_221)
);

CKINVDCx9p33_ASAP7_75t_R g173 ( 
.A(n_102),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_107),
.A2(n_61),
.B1(n_12),
.B2(n_51),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_61),
.B1(n_131),
.B2(n_98),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_186),
.B1(n_148),
.B2(n_129),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_99),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_119),
.B1(n_104),
.B2(n_144),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_128),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_182),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_183),
.Y(n_220)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_116),
.B1(n_108),
.B2(n_126),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_114),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_115),
.A2(n_130),
.B1(n_150),
.B2(n_132),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_122),
.B(n_112),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_115),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_123),
.B1(n_127),
.B2(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_203),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_173),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_133),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_206),
.B1(n_212),
.B2(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_104),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_171),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_129),
.B1(n_150),
.B2(n_111),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_221),
.A2(n_151),
.B1(n_179),
.B2(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_167),
.A2(n_186),
.B1(n_181),
.B2(n_151),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_187),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_156),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_158),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_235),
.A2(n_237),
.B(n_242),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_218),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_152),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_185),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_202),
.Y(n_239)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_163),
.B(n_167),
.C(n_193),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_213),
.B(n_207),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_153),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_168),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_248),
.C(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_215),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_179),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_204),
.B1(n_212),
.B2(n_221),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_254),
.B1(n_263),
.B2(n_270),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_195),
.B1(n_194),
.B2(n_203),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_260),
.B(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_194),
.C(n_201),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_231),
.C(n_227),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_216),
.B1(n_199),
.B2(n_201),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_227),
.A2(n_199),
.B1(n_213),
.B2(n_222),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_240),
.B1(n_233),
.B2(n_244),
.Y(n_278)
);

AOI22x1_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_215),
.B1(n_184),
.B2(n_191),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_222),
.B1(n_219),
.B2(n_205),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_226),
.B(n_224),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_290),
.B(n_267),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_262),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_276),
.C(n_282),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_285),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_268),
.B(n_225),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_277),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_279),
.B1(n_287),
.B2(n_288),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_265),
.B1(n_251),
.B2(n_261),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_234),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_232),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_286),
.C(n_254),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_264),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_236),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_229),
.B1(n_230),
.B2(n_239),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_226),
.B1(n_246),
.B2(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_257),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_267),
.B(n_263),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_292),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_270),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_256),
.B(n_215),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_258),
.B1(n_250),
.B2(n_257),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_298),
.B1(n_279),
.B2(n_278),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_266),
.B1(n_249),
.B2(n_252),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_252),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_304),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_266),
.C(n_249),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_242),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_286),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_318),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_301),
.B1(n_299),
.B2(n_297),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_276),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_314),
.B(n_306),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_284),
.C(n_274),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_315),
.B(n_291),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_283),
.B1(n_287),
.B2(n_289),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_272),
.B1(n_290),
.B2(n_256),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_296),
.C(n_304),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_328),
.C(n_334),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_295),
.Y(n_326)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_326),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_309),
.A2(n_294),
.B(n_298),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_247),
.B(n_161),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_331),
.A2(n_247),
.B1(n_256),
.B2(n_217),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_318),
.B1(n_313),
.B2(n_315),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_303),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_316),
.B1(n_308),
.B2(n_309),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_336),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_237),
.B1(n_321),
.B2(n_311),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_343),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_323),
.B(n_326),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_341),
.A2(n_190),
.B(n_175),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_330),
.A2(n_208),
.B1(n_192),
.B2(n_205),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_345),
.A2(n_336),
.B1(n_341),
.B2(n_333),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_339),
.B(n_328),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_349),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_342),
.B(n_325),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_208),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_334),
.C(n_333),
.Y(n_349)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_355),
.A2(n_356),
.B(n_166),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_344),
.A2(n_335),
.B(n_343),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_357),
.B(n_350),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_357),
.B(n_353),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_358),
.A2(n_165),
.B(n_164),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_354),
.A2(n_350),
.B1(n_192),
.B2(n_162),
.Y(n_359)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_359),
.A2(n_360),
.B(n_361),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_362),
.B(n_177),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_134),
.C(n_177),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_366),
.B(n_363),
.C(n_134),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_111),
.Y(n_368)
);


endmodule