module fake_netlist_6_643_n_2147 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2147);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2147;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_1),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_84),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_3),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_47),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_56),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_143),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_90),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_44),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_96),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_146),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_179),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_105),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_82),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_6),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_205),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_51),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_139),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_77),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

BUFx2_ASAP7_75t_SL g246 ( 
.A(n_192),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_2),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_154),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_173),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_97),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_64),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_21),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_98),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_212),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_163),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_124),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_158),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_171),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_165),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_12),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_67),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_31),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_122),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_64),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_57),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_137),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_91),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_164),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_63),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_83),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_144),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_18),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_86),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_194),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_4),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_142),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_99),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_24),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_76),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_186),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_120),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_69),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_115),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_6),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_27),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_172),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_61),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_216),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_108),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_114),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_147),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_131),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_183),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_58),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_59),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_196),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_80),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_140),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_161),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_1),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_152),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_79),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_81),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_88),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_180),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_19),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_199),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_29),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_5),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_33),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_61),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_201),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_37),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_44),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_198),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_11),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_69),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_50),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_193),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_141),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_155),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_134),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_16),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_89),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_102),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_93),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_118),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_31),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_34),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_136),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_42),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_92),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_184),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_74),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_85),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_77),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_187),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_24),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_22),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_185),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_191),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_4),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_34),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_209),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_56),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_126),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_20),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_162),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_0),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_16),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_197),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_0),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_95),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_13),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_167),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_202),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_21),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_175),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_190),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_109),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_78),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_207),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_20),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_35),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_52),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_48),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_50),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_128),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_49),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_78),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_58),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_38),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_133),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_70),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_217),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_53),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_22),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_57),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_75),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_63),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_119),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_39),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_9),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_113),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_23),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_138),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_55),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_33),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_151),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_49),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_129),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_160),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_74),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_206),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_35),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_211),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_14),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_116),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_170),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_42),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_107),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_29),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_8),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_75),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_117),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_76),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_66),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_159),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_9),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_150),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_188),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_156),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_30),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_48),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_195),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_62),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_121),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_215),
.Y(n_428)
);

BUFx8_ASAP7_75t_SL g429 ( 
.A(n_59),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_242),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_429),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_261),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_272),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_247),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_247),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_220),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_229),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_247),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_295),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_331),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_247),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_247),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_222),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_232),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_222),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_340),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_234),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_222),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_301),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_253),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_298),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_277),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_277),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_384),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_301),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_235),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_240),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_251),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_228),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_252),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_218),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_269),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_228),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_230),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_263),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_264),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_230),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_265),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_250),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_250),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_256),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_256),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_275),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_266),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_279),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_221),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_329),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_280),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_329),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_297),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_266),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_372),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_223),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_270),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_270),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_225),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_271),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_237),
.B(n_2),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_271),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_281),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_281),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_285),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_296),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_296),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_300),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_300),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_268),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_289),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_391),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_304),
.B(n_3),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_303),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_304),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_268),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_239),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_318),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_318),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_319),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_351),
.B(n_7),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_351),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_243),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_319),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_248),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_324),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_324),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_327),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_406),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_327),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_306),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_328),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_299),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_309),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_328),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_268),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_311),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_338),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_314),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_317),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_325),
.Y(n_529)
);

INVxp33_ASAP7_75t_L g530 ( 
.A(n_338),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_330),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_334),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_336),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_337),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_254),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_257),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_353),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_353),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_342),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_359),
.Y(n_540)
);

BUFx8_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_434),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_521),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_510),
.A2(n_241),
.B1(n_321),
.B2(n_258),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_435),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_435),
.B(n_404),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_509),
.B(n_404),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_438),
.B(n_260),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_443),
.B(n_298),
.Y(n_550)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_438),
.A2(n_226),
.B(n_219),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_441),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_449),
.B(n_455),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_521),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_441),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_442),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_521),
.Y(n_559)
);

AND3x2_ASAP7_75t_L g560 ( 
.A(n_478),
.B(n_236),
.C(n_224),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_442),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_445),
.B(n_260),
.Y(n_563)
);

INVxp33_ASAP7_75t_SL g564 ( 
.A(n_436),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_445),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_443),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_451),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_448),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_477),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_448),
.B(n_320),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_460),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_452),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_464),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_452),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_464),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_489),
.B(n_268),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_453),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_465),
.B(n_224),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_465),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_468),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_470),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_454),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_471),
.B(n_347),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_471),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_519),
.Y(n_589)
);

OA21x2_ASAP7_75t_L g590 ( 
.A1(n_458),
.A2(n_226),
.B(n_219),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_458),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_473),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_473),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_475),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_475),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_482),
.B(n_428),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_482),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_485),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_480),
.B(n_485),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_486),
.B(n_236),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_486),
.B(n_427),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_488),
.B(n_320),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_488),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_491),
.B(n_278),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_484),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_491),
.B(n_354),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_487),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_326),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_492),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_494),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_505),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_495),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_495),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_496),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_496),
.B(n_358),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_497),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_511),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_503),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_503),
.B(n_278),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_506),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_507),
.B(n_363),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_507),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_508),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_508),
.B(n_282),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_512),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_498),
.A2(n_333),
.B1(n_360),
.B2(n_390),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_567),
.B(n_450),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_542),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_587),
.B(n_513),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_542),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_548),
.B(n_437),
.Y(n_636)
);

INVxp33_ASAP7_75t_L g637 ( 
.A(n_558),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_599),
.B(n_246),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_599),
.B(n_444),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_543),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_567),
.B(n_450),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_548),
.A2(n_501),
.B1(n_398),
.B2(n_413),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_567),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_543),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_629),
.B(n_430),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_543),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_560),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_613),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_599),
.B(n_447),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_613),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_613),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_564),
.B(n_463),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_545),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_560),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_613),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_545),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_558),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_587),
.B(n_456),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_590),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_565),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_565),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_565),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_615),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_578),
.A2(n_501),
.B1(n_398),
.B2(n_413),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_564),
.B(n_463),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_607),
.B(n_481),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_546),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_543),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_569),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_546),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_596),
.B(n_457),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_544),
.B(n_483),
.C(n_481),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_552),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_615),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_615),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_568),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_615),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_552),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_R g683 ( 
.A(n_569),
.B(n_431),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_596),
.B(n_459),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_569),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_555),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_607),
.B(n_483),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_605),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_553),
.B(n_461),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_556),
.Y(n_693)
);

BUFx4f_ASAP7_75t_L g694 ( 
.A(n_551),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_578),
.A2(n_237),
.B1(n_326),
.B2(n_359),
.Y(n_695)
);

NOR2x1p5_ASAP7_75t_L g696 ( 
.A(n_547),
.B(n_373),
.Y(n_696)
);

AND3x1_ASAP7_75t_L g697 ( 
.A(n_553),
.B(n_381),
.C(n_373),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_556),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_601),
.B(n_466),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_541),
.B(n_467),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_541),
.B(n_469),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_613),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_578),
.A2(n_387),
.B1(n_389),
.B2(n_381),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_615),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_601),
.B(n_474),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_606),
.B(n_476),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_615),
.Y(n_708)
);

AND2x2_ASAP7_75t_SL g709 ( 
.A(n_551),
.B(n_282),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_578),
.A2(n_389),
.B1(n_392),
.B2(n_387),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_606),
.B(n_536),
.C(n_535),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_554),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_620),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_561),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_554),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_620),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_620),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_605),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_554),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_550),
.B(n_512),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_605),
.Y(n_721)
);

AND2x6_ASAP7_75t_L g722 ( 
.A(n_550),
.B(n_286),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_578),
.A2(n_397),
.B1(n_403),
.B2(n_392),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_616),
.B(n_479),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_613),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_589),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_612),
.A2(n_352),
.B1(n_323),
.B2(n_267),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_541),
.B(n_493),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_554),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_616),
.B(n_502),
.C(n_499),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_600),
.A2(n_403),
.B1(n_405),
.B2(n_397),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_620),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_590),
.Y(n_733)
);

BUFx4f_ASAP7_75t_L g734 ( 
.A(n_551),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_557),
.Y(n_735)
);

INVxp33_ASAP7_75t_L g736 ( 
.A(n_544),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_561),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_613),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_598),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_620),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_612),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_541),
.B(n_522),
.Y(n_742)
);

BUFx4f_ASAP7_75t_L g743 ( 
.A(n_551),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_612),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_624),
.B(n_498),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_618),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_541),
.B(n_525),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_624),
.B(n_529),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_598),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_598),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_576),
.A2(n_528),
.B1(n_539),
.B2(n_527),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_590),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_620),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_557),
.B(n_531),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_SL g755 ( 
.A(n_618),
.B(n_284),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_590),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_598),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_598),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_620),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_557),
.B(n_532),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_557),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_618),
.A2(n_504),
.B1(n_524),
.B2(n_576),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_562),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_629),
.A2(n_374),
.B1(n_291),
.B2(n_293),
.Y(n_764)
);

AOI21x1_ASAP7_75t_L g765 ( 
.A1(n_549),
.A2(n_233),
.B(n_231),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_562),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_620),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_626),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_591),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_547),
.B(n_533),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_568),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_602),
.B(n_534),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_550),
.B(n_514),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_626),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_591),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_571),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_626),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_591),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_571),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_557),
.Y(n_780)
);

CKINVDCx14_ASAP7_75t_R g781 ( 
.A(n_589),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_626),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_626),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_563),
.B(n_246),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_662),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_706),
.B(n_770),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_691),
.B(n_563),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_662),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_763),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_662),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_660),
.B(n_563),
.Y(n_791)
);

NAND2x1p5_ASAP7_75t_L g792 ( 
.A(n_661),
.B(n_551),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_675),
.B(n_563),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_751),
.B(n_432),
.Y(n_794)
);

OAI221xp5_ASAP7_75t_L g795 ( 
.A1(n_644),
.A2(n_537),
.B1(n_523),
.B2(n_490),
.C(n_287),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_663),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_763),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_684),
.B(n_563),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_722),
.B(n_365),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_663),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_766),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_SL g802 ( 
.A(n_636),
.B(n_433),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_638),
.A2(n_440),
.B1(n_446),
.B2(n_439),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_766),
.Y(n_804)
);

INVx8_ASAP7_75t_L g805 ( 
.A(n_638),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_699),
.B(n_626),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_685),
.B(n_570),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_722),
.B(n_366),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_776),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_761),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_709),
.A2(n_417),
.B1(n_405),
.B2(n_600),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_694),
.B(n_299),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_707),
.B(n_626),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_640),
.A2(n_549),
.B(n_575),
.C(n_573),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_724),
.B(n_626),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_659),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_694),
.B(n_734),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_663),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_651),
.A2(n_517),
.B1(n_500),
.B2(n_322),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_633),
.B(n_504),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_748),
.B(n_568),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_659),
.B(n_524),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_664),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_664),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_776),
.B(n_568),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_779),
.B(n_568),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_779),
.B(n_709),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_673),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_694),
.B(n_299),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_645),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_720),
.B(n_602),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_694),
.B(n_299),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_645),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_730),
.B(n_573),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_734),
.B(n_299),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_754),
.A2(n_559),
.B(n_600),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_703),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_639),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_734),
.B(n_361),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_709),
.B(n_568),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_760),
.B(n_559),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_720),
.B(n_602),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_664),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_633),
.B(n_227),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_734),
.B(n_361),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_773),
.B(n_631),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_743),
.B(n_361),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_773),
.B(n_559),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_631),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_634),
.B(n_559),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_639),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_743),
.B(n_361),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_673),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_743),
.B(n_361),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_743),
.B(n_566),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_685),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_690),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_638),
.A2(n_313),
.B1(n_290),
.B2(n_343),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_703),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_661),
.A2(n_417),
.B1(n_604),
.B2(n_600),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_718),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_690),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_703),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_762),
.B(n_687),
.C(n_669),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_SL g865 ( 
.A(n_746),
.B(n_726),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_634),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_711),
.B(n_575),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_655),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_655),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_745),
.B(n_566),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_658),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_638),
.A2(n_233),
.B1(n_238),
.B2(n_231),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_658),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_670),
.B(n_559),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_745),
.B(n_566),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_670),
.B(n_566),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_661),
.B(n_566),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_772),
.A2(n_604),
.B(n_600),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_746),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_696),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_667),
.B(n_566),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_667),
.A2(n_733),
.B(n_756),
.C(n_752),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_674),
.B(n_566),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_761),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_674),
.B(n_566),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_667),
.A2(n_579),
.B(n_582),
.C(n_580),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_703),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_677),
.B(n_604),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_726),
.B(n_294),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_SL g890 ( 
.A(n_733),
.B(n_752),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_733),
.B(n_286),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_677),
.B(n_604),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_752),
.B(n_322),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_756),
.B(n_399),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_712),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_638),
.A2(n_420),
.B1(n_422),
.B2(n_369),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_639),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_712),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_697),
.B(n_570),
.C(n_608),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_712),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_649),
.B(n_472),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_682),
.B(n_604),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_756),
.B(n_399),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_761),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_722),
.A2(n_627),
.B1(n_621),
.B2(n_348),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_682),
.B(n_621),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_649),
.B(n_608),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_656),
.A2(n_370),
.B1(n_415),
.B2(n_378),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_712),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_715),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_SL g911 ( 
.A(n_700),
.B(n_701),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_656),
.A2(n_383),
.B1(n_402),
.B2(n_411),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_718),
.B(n_570),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_715),
.B(n_621),
.Y(n_914)
);

AOI221xp5_ASAP7_75t_L g915 ( 
.A1(n_736),
.A2(n_530),
.B1(n_288),
.B2(n_349),
.C(n_316),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_715),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_715),
.B(n_621),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_719),
.B(n_729),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_719),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_686),
.B(n_692),
.Y(n_920)
);

BUFx5_ASAP7_75t_L g921 ( 
.A(n_722),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_630),
.B(n_643),
.Y(n_922)
);

INVxp33_ASAP7_75t_L g923 ( 
.A(n_637),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_L g924 ( 
.A(n_722),
.B(n_385),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_722),
.A2(n_401),
.B1(n_396),
.B2(n_394),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_719),
.Y(n_926)
);

OAI22xp33_ASAP7_75t_L g927 ( 
.A1(n_727),
.A2(n_238),
.B1(n_244),
.B2(n_425),
.Y(n_927)
);

O2A1O1Ixp5_ASAP7_75t_L g928 ( 
.A1(n_739),
.A2(n_621),
.B(n_627),
.C(n_276),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_719),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_780),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_722),
.A2(n_627),
.B1(n_244),
.B2(n_245),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_686),
.B(n_627),
.Y(n_932)
);

INVx8_ASAP7_75t_L g933 ( 
.A(n_784),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_729),
.B(n_627),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_741),
.B(n_608),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_784),
.A2(n_308),
.B1(n_425),
.B2(n_421),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_741),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_780),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_729),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_729),
.B(n_577),
.Y(n_940)
);

OAI21xp33_ASAP7_75t_L g941 ( 
.A1(n_666),
.A2(n_515),
.B(n_514),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_735),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_735),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_692),
.B(n_591),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_704),
.A2(n_307),
.B1(n_421),
.B2(n_418),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_693),
.B(n_591),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_696),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_735),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_710),
.A2(n_731),
.B1(n_723),
.B2(n_695),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_693),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_735),
.B(n_577),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_698),
.B(n_591),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_698),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_780),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_714),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_714),
.B(n_591),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_849),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_855),
.A2(n_749),
.B(n_739),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_812),
.A2(n_750),
.B(n_749),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_937),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_849),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_810),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_866),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_840),
.A2(n_689),
.B(n_680),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_786),
.B(n_744),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_817),
.A2(n_689),
.B(n_680),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_817),
.A2(n_855),
.B(n_821),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_787),
.B(n_737),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_791),
.B(n_737),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_812),
.A2(n_757),
.B(n_750),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_806),
.A2(n_689),
.B(n_680),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_829),
.A2(n_758),
.B(n_757),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_829),
.A2(n_758),
.B(n_652),
.Y(n_973)
);

AOI21x1_ASAP7_75t_L g974 ( 
.A1(n_877),
.A2(n_652),
.B(n_650),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_813),
.A2(n_689),
.B(n_680),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_793),
.A2(n_798),
.B1(n_922),
.B2(n_875),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_832),
.A2(n_653),
.B(n_650),
.Y(n_977)
);

AOI21x1_ASAP7_75t_L g978 ( 
.A1(n_877),
.A2(n_657),
.B(n_653),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_846),
.B(n_784),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_844),
.B(n_784),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_816),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_815),
.A2(n_771),
.B(n_635),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_868),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_913),
.B(n_744),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_868),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_921),
.B(n_632),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_869),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_844),
.B(n_784),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_921),
.B(n_632),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_869),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_881),
.A2(n_771),
.B(n_635),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_L g992 ( 
.A(n_819),
.B(n_676),
.C(n_668),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_881),
.A2(n_771),
.B(n_635),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_841),
.A2(n_771),
.B(n_635),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_811),
.B(n_632),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_811),
.B(n_632),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_832),
.A2(n_725),
.B(n_657),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_871),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_921),
.B(n_641),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_827),
.A2(n_742),
.B(n_747),
.C(n_728),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_835),
.A2(n_845),
.B(n_839),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_871),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_901),
.B(n_822),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_835),
.A2(n_845),
.B(n_839),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_847),
.A2(n_738),
.B(n_725),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_873),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_789),
.B(n_641),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_847),
.A2(n_702),
.B(n_738),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_873),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_852),
.A2(n_671),
.B(n_665),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_852),
.A2(n_702),
.B(n_753),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_820),
.B(n_828),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_922),
.A2(n_654),
.B1(n_755),
.B2(n_683),
.Y(n_1013)
);

OAI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_901),
.A2(n_727),
.B(n_764),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_854),
.A2(n_702),
.B(n_753),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_797),
.B(n_641),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_801),
.B(n_641),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_820),
.A2(n_721),
.B(n_764),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_814),
.A2(n_882),
.B(n_886),
.C(n_899),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_854),
.A2(n_702),
.B(n_753),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_807),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_860),
.A2(n_249),
.B1(n_255),
.B2(n_245),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_804),
.B(n_642),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_915),
.A2(n_255),
.B(n_259),
.C(n_249),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_809),
.B(n_642),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_955),
.B(n_642),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_838),
.A2(n_702),
.B(n_753),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_807),
.B(n_726),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_L g1029 ( 
.A(n_803),
.B(n_765),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_853),
.Y(n_1030)
);

OAI321xp33_ASAP7_75t_L g1031 ( 
.A1(n_927),
.A2(n_350),
.A3(n_368),
.B1(n_345),
.B2(n_356),
.C(n_259),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_807),
.B(n_726),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_891),
.A2(n_671),
.B(n_665),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_950),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_935),
.Y(n_1035)
);

INVxp33_ASAP7_75t_SL g1036 ( 
.A(n_802),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_891),
.A2(n_671),
.B(n_665),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_838),
.A2(n_702),
.B(n_753),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_950),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_953),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_831),
.B(n_579),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_810),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_851),
.A2(n_759),
.B(n_753),
.Y(n_1043)
);

NOR2xp67_ASAP7_75t_SL g1044 ( 
.A(n_884),
.B(n_262),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_953),
.Y(n_1045)
);

OAI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_794),
.A2(n_335),
.B1(n_332),
.B2(n_418),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_851),
.A2(n_774),
.B(n_759),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_831),
.B(n_842),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_861),
.B(n_781),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_920),
.B(n_642),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_785),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_893),
.A2(n_679),
.B(n_678),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_897),
.A2(n_774),
.B(n_759),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_785),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_860),
.B(n_648),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_842),
.B(n_907),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_949),
.A2(n_356),
.B(n_273),
.C(n_274),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_837),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_859),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_945),
.A2(n_308),
.B1(n_408),
.B2(n_409),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_893),
.A2(n_679),
.B(n_678),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_863),
.Y(n_1062)
);

INVx8_ASAP7_75t_L g1063 ( 
.A(n_805),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_907),
.B(n_648),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_796),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_894),
.A2(n_273),
.B(n_262),
.C(n_274),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_810),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_830),
.B(n_647),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_870),
.B(n_648),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_870),
.B(n_648),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_875),
.B(n_678),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_848),
.B(n_679),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_894),
.A2(n_688),
.B(n_681),
.Y(n_1073)
);

BUFx4f_ASAP7_75t_L g1074 ( 
.A(n_833),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_921),
.B(n_639),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_949),
.B(n_681),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_895),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_856),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_884),
.B(n_681),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_890),
.B(n_639),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_810),
.Y(n_1081)
);

BUFx4f_ASAP7_75t_L g1082 ( 
.A(n_805),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_954),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_930),
.B(n_639),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_898),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_904),
.B(n_688),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_904),
.B(n_688),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_938),
.B(n_705),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_805),
.B(n_276),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_945),
.A2(n_864),
.B(n_941),
.C(n_858),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_938),
.B(n_705),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_921),
.B(n_672),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_954),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_954),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_834),
.B(n_705),
.Y(n_1095)
);

BUFx4f_ASAP7_75t_L g1096 ( 
.A(n_857),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_897),
.A2(n_774),
.B(n_759),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_880),
.A2(n_350),
.B(n_292),
.C(n_302),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_888),
.B(n_708),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_921),
.B(n_672),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_862),
.B(n_647),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_892),
.B(n_708),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_903),
.A2(n_713),
.B(n_708),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_947),
.B(n_580),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_903),
.A2(n_774),
.B(n_759),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_L g1106 ( 
.A(n_930),
.B(n_713),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_911),
.A2(n_345),
.B(n_292),
.C(n_302),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_902),
.B(n_713),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_879),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_914),
.A2(n_777),
.B(n_774),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_906),
.B(n_716),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_792),
.A2(n_717),
.B(n_716),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_932),
.B(n_878),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_923),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_917),
.A2(n_777),
.B(n_775),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_896),
.B(n_765),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_917),
.A2(n_777),
.B(n_775),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_905),
.B(n_672),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_934),
.A2(n_777),
.B(n_769),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_792),
.A2(n_717),
.B(n_716),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_934),
.A2(n_918),
.B(n_836),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_900),
.B(n_717),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_905),
.B(n_672),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_867),
.A2(n_283),
.B(n_307),
.C(n_315),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_918),
.A2(n_783),
.B1(n_782),
.B2(n_767),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_865),
.B(n_305),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_940),
.A2(n_740),
.B(n_732),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_936),
.A2(n_283),
.B(n_315),
.C(n_332),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_799),
.A2(n_777),
.B(n_769),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_909),
.A2(n_783),
.B1(n_782),
.B2(n_732),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_872),
.A2(n_409),
.B(n_335),
.C(n_368),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_954),
.B(n_672),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_910),
.B(n_732),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_808),
.A2(n_777),
.B(n_778),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_924),
.A2(n_778),
.B(n_767),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_850),
.A2(n_783),
.B(n_767),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_795),
.A2(n_408),
.B(n_588),
.C(n_582),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_874),
.A2(n_782),
.B(n_768),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_916),
.B(n_740),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_887),
.A2(n_768),
.B(n_740),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_908),
.B(n_912),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_919),
.A2(n_768),
.B(n_672),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_939),
.A2(n_646),
.B(n_594),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_931),
.A2(n_583),
.B1(n_628),
.B2(n_584),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_926),
.A2(n_597),
.B(n_628),
.C(n_584),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_929),
.A2(n_593),
.B1(n_625),
.B2(n_594),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_942),
.B(n_943),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_948),
.B(n_593),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1113),
.A2(n_931),
.B(n_933),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_SL g1150 ( 
.A1(n_965),
.A2(n_889),
.B(n_925),
.C(n_788),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_960),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_R g1152 ( 
.A(n_1109),
.B(n_933),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1135),
.A2(n_883),
.B(n_876),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_992),
.A2(n_933),
.B1(n_951),
.B2(n_940),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1051),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1014),
.A2(n_928),
.B(n_825),
.C(n_826),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_963),
.Y(n_1157)
);

AND2x2_ASAP7_75t_SL g1158 ( 
.A(n_992),
.B(n_885),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_976),
.A2(n_956),
.B1(n_952),
.B2(n_946),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_965),
.A2(n_944),
.B1(n_951),
.B2(n_843),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1036),
.B(n_796),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1013),
.B(n_312),
.C(n_310),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_990),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1067),
.B(n_818),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1004),
.A2(n_843),
.B1(n_824),
.B2(n_823),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_L g1166 ( 
.A(n_980),
.B(n_818),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1012),
.B(n_823),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1003),
.B(n_824),
.Y(n_1168)
);

OAI22x1_ASAP7_75t_L g1169 ( 
.A1(n_1012),
.A2(n_412),
.B1(n_339),
.B2(n_346),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1001),
.A2(n_800),
.B(n_790),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_998),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1019),
.A2(n_597),
.B(n_588),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_988),
.B(n_583),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1126),
.B(n_1018),
.C(n_1101),
.Y(n_1174)
);

OAI21xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1118),
.A2(n_592),
.B(n_623),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1068),
.A2(n_377),
.B1(n_426),
.B2(n_424),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_995),
.A2(n_592),
.B1(n_595),
.B2(n_623),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1054),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1141),
.B(n_595),
.Y(n_1179)
);

NOR3xp33_ASAP7_75t_L g1180 ( 
.A(n_1126),
.B(n_1068),
.C(n_1046),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_968),
.B(n_593),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_984),
.B(n_610),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1034),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1057),
.A2(n_617),
.B(n_619),
.C(n_610),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1057),
.A2(n_617),
.B(n_619),
.C(n_625),
.Y(n_1185)
);

AO22x1_ASAP7_75t_L g1186 ( 
.A1(n_1101),
.A2(n_395),
.B1(n_393),
.B2(n_388),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1114),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_967),
.A2(n_646),
.B(n_625),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1039),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_969),
.B(n_594),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1065),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_SL g1192 ( 
.A(n_1046),
.B(n_1024),
.C(n_1031),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1048),
.B(n_515),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1041),
.B(n_516),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_R g1195 ( 
.A(n_1096),
.B(n_341),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_957),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1090),
.B(n_603),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1090),
.B(n_603),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1049),
.B(n_294),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1056),
.B(n_603),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1041),
.B(n_516),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1063),
.B(n_518),
.Y(n_1202)
);

AOI21x1_ASAP7_75t_L g1203 ( 
.A1(n_958),
.A2(n_581),
.B(n_572),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_996),
.A2(n_419),
.B1(n_355),
.B2(n_357),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_961),
.Y(n_1205)
);

NAND2xp33_ASAP7_75t_R g1206 ( 
.A(n_1028),
.B(n_87),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1024),
.A2(n_622),
.B(n_614),
.C(n_611),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_R g1208 ( 
.A(n_1096),
.B(n_344),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1035),
.A2(n_376),
.B(n_375),
.Y(n_1209)
);

AOI33xp33_ASAP7_75t_L g1210 ( 
.A1(n_1060),
.A2(n_518),
.A3(n_520),
.B1(n_526),
.B2(n_538),
.B3(n_540),
.Y(n_1210)
);

NOR3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1098),
.B(n_400),
.C(n_362),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1000),
.A2(n_371),
.B(n_364),
.C(n_423),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1029),
.A2(n_622),
.B1(n_614),
.B2(n_611),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1114),
.B(n_520),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1035),
.B(n_367),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_979),
.A2(n_382),
.B(n_380),
.C(n_416),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1022),
.A2(n_1124),
.B(n_1145),
.C(n_1107),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1030),
.B(n_294),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_983),
.B(n_609),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1078),
.B(n_386),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_985),
.B(n_609),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1055),
.A2(n_622),
.B(n_614),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_964),
.A2(n_646),
.B(n_611),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1074),
.B(n_609),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_987),
.B(n_572),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1002),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1074),
.B(n_407),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1080),
.A2(n_410),
.B1(n_414),
.B2(n_585),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_981),
.B(n_572),
.Y(n_1229)
);

OR2x2_ASAP7_75t_SL g1230 ( 
.A(n_1021),
.B(n_1078),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1021),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1006),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_1104),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1112),
.A2(n_646),
.B(n_586),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1049),
.B(n_294),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1032),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1120),
.A2(n_646),
.B(n_586),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1104),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1009),
.Y(n_1239)
);

AO21x1_ASAP7_75t_L g1240 ( 
.A1(n_1121),
.A2(n_540),
.B(n_538),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1040),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1045),
.B(n_574),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1063),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1107),
.A2(n_586),
.B(n_585),
.C(n_581),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1089),
.B(n_379),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1058),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1064),
.B(n_379),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_962),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_962),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1080),
.A2(n_585),
.B1(n_581),
.B2(n_574),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1063),
.Y(n_1251)
);

OAI21xp33_ASAP7_75t_L g1252 ( 
.A1(n_1060),
.A2(n_1098),
.B(n_1128),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1050),
.B(n_574),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_962),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_SL g1255 ( 
.A1(n_1089),
.A2(n_526),
.B1(n_379),
.B2(n_10),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1072),
.B(n_577),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1075),
.A2(n_1100),
.B(n_1092),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_R g1258 ( 
.A(n_1082),
.B(n_94),
.Y(n_1258)
);

O2A1O1Ixp5_ASAP7_75t_SL g1259 ( 
.A1(n_1132),
.A2(n_379),
.B(n_8),
.C(n_10),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1144),
.A2(n_577),
.B(n_12),
.C(n_13),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1092),
.A2(n_577),
.B(n_200),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1082),
.A2(n_1118),
.B1(n_1123),
.B2(n_1076),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1042),
.B(n_577),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_962),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1059),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1067),
.B(n_577),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1062),
.B(n_7),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1100),
.A2(n_189),
.B(n_181),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1077),
.B(n_14),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1089),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1085),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1099),
.B(n_17),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1148),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1116),
.A2(n_178),
.B1(n_177),
.B2(n_174),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1007),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1102),
.B(n_17),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1122),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1067),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1123),
.A2(n_157),
.B1(n_153),
.B2(n_148),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1067),
.B(n_145),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1042),
.B(n_135),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1133),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1083),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1095),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_982),
.A2(n_132),
.B(n_130),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1139),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1083),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1071),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_1288)
);

BUFx2_ASAP7_75t_R g1289 ( 
.A(n_1132),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_971),
.A2(n_975),
.B(n_994),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1081),
.B(n_127),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1081),
.B(n_125),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_R g1293 ( 
.A(n_1093),
.B(n_123),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1108),
.B(n_25),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1093),
.A2(n_112),
.B1(n_111),
.B2(n_110),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1111),
.A2(n_106),
.B(n_104),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1094),
.B(n_25),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1084),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1094),
.B(n_103),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_959),
.A2(n_101),
.B1(n_100),
.B2(n_28),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1147),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1069),
.B(n_26),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1127),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1070),
.B(n_32),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1044),
.A2(n_1106),
.B1(n_1147),
.B2(n_1017),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_966),
.A2(n_32),
.B(n_36),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1084),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1128),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1016),
.Y(n_1309)
);

NAND2xp33_ASAP7_75t_R g1310 ( 
.A(n_1079),
.B(n_40),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1023),
.B(n_40),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_970),
.A2(n_41),
.B(n_43),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_991),
.A2(n_79),
.B(n_45),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_993),
.A2(n_41),
.B(n_45),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1149),
.A2(n_1129),
.B(n_1134),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1174),
.B(n_1137),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1203),
.A2(n_978),
.B(n_974),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1180),
.B(n_1025),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1167),
.B(n_1026),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_SL g1320 ( 
.A1(n_1312),
.A2(n_972),
.B(n_973),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1290),
.A2(n_1020),
.B(n_1011),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1155),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1180),
.A2(n_1131),
.B(n_1066),
.C(n_986),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1193),
.B(n_1088),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1240),
.A2(n_1262),
.A3(n_1159),
.B(n_1212),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1235),
.A2(n_1138),
.B(n_1136),
.C(n_1008),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1188),
.A2(n_1153),
.B(n_1170),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1263),
.A2(n_1015),
.B(n_999),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1156),
.A2(n_1105),
.A3(n_1110),
.B(n_1027),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1192),
.A2(n_1117),
.B(n_1115),
.C(n_1119),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1187),
.B(n_1066),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_SL g1332 ( 
.A1(n_1150),
.A2(n_986),
.B(n_989),
.C(n_999),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1300),
.A2(n_1038),
.A3(n_1043),
.B(n_1053),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1193),
.B(n_1086),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1162),
.A2(n_989),
.B(n_997),
.C(n_977),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1187),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1278),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1181),
.A2(n_1047),
.B(n_1097),
.Y(n_1338)
);

AO32x2_ASAP7_75t_L g1339 ( 
.A1(n_1177),
.A2(n_1010),
.A3(n_1005),
.B1(n_1073),
.B2(n_1061),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1223),
.A2(n_1103),
.B(n_1037),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1190),
.A2(n_1087),
.B(n_1091),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1166),
.A2(n_1033),
.B(n_1052),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1165),
.A2(n_1142),
.B(n_1140),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_L g1344 ( 
.A(n_1238),
.B(n_1125),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1151),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1246),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1243),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1233),
.B(n_1146),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1265),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_51),
.C(n_52),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1231),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1178),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1214),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1158),
.A2(n_1198),
.B(n_1197),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1256),
.A2(n_1130),
.B(n_53),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1192),
.A2(n_1217),
.B(n_1247),
.C(n_1252),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1191),
.Y(n_1357)
);

AND2x4_ASAP7_75t_SL g1358 ( 
.A(n_1251),
.B(n_46),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1253),
.A2(n_46),
.B(n_54),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1217),
.A2(n_54),
.B(n_55),
.C(n_60),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1277),
.B(n_60),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1303),
.A2(n_1160),
.A3(n_1237),
.B(n_1234),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1257),
.A2(n_62),
.B(n_65),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1173),
.A2(n_65),
.B(n_66),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_SL g1365 ( 
.A(n_1278),
.B(n_67),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1306),
.A2(n_68),
.A3(n_70),
.B(n_71),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1282),
.B(n_68),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1286),
.B(n_71),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1284),
.B(n_1233),
.Y(n_1369)
);

AOI221x1_ASAP7_75t_L g1370 ( 
.A1(n_1313),
.A2(n_72),
.B1(n_73),
.B2(n_1314),
.C(n_1279),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1172),
.A2(n_1158),
.B(n_1222),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1152),
.Y(n_1372)
);

NOR2xp67_ASAP7_75t_L g1373 ( 
.A(n_1220),
.B(n_1284),
.Y(n_1373)
);

BUFx2_ASAP7_75t_SL g1374 ( 
.A(n_1278),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1175),
.A2(n_1304),
.B(n_1302),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1168),
.B(n_1273),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1194),
.B(n_1201),
.Y(n_1377)
);

AOI221x1_ASAP7_75t_L g1378 ( 
.A1(n_1169),
.A2(n_1285),
.B1(n_1294),
.B2(n_1276),
.C(n_1272),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1261),
.A2(n_1219),
.B(n_1221),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1231),
.Y(n_1380)
);

BUFx12f_ASAP7_75t_L g1381 ( 
.A(n_1270),
.Y(n_1381)
);

CKINVDCx11_ASAP7_75t_R g1382 ( 
.A(n_1202),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1179),
.A2(n_1200),
.B(n_1225),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1250),
.A2(n_1216),
.A3(n_1297),
.B(n_1309),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1275),
.A2(n_1154),
.B(n_1305),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1271),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_SL g1387 ( 
.A(n_1289),
.B(n_1260),
.Y(n_1387)
);

INVx5_ASAP7_75t_L g1388 ( 
.A(n_1254),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1296),
.A2(n_1213),
.B(n_1291),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1242),
.A2(n_1244),
.B(n_1164),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_SL g1391 ( 
.A1(n_1299),
.A2(n_1280),
.B(n_1281),
.C(n_1292),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1259),
.A2(n_1185),
.B(n_1207),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1268),
.A2(n_1266),
.B(n_1161),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1267),
.A2(n_1269),
.A3(n_1228),
.B(n_1163),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1288),
.A2(n_1260),
.B1(n_1301),
.B2(n_1171),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1157),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1287),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1185),
.A2(n_1207),
.B(n_1184),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1288),
.A2(n_1183),
.B1(n_1189),
.B2(n_1274),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1194),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1164),
.A2(n_1298),
.B(n_1182),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1196),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1298),
.A2(n_1264),
.B(n_1241),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1298),
.A2(n_1264),
.B(n_1239),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1201),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1215),
.B(n_1218),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1298),
.A2(n_1226),
.B(n_1232),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1311),
.Y(n_1408)
);

BUFx2_ASAP7_75t_SL g1409 ( 
.A(n_1254),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1236),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1206),
.A2(n_1310),
.B1(n_1255),
.B2(n_1311),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1199),
.A2(n_1211),
.B(n_1308),
.C(n_1209),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1308),
.A2(n_1184),
.B(n_1210),
.C(n_1295),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1230),
.A2(n_1202),
.B1(n_1307),
.B2(n_1254),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1204),
.A2(n_1244),
.A3(n_1224),
.B(n_1293),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1229),
.A2(n_1283),
.B(n_1202),
.Y(n_1416)
);

OA22x2_ASAP7_75t_L g1417 ( 
.A1(n_1176),
.A2(n_1245),
.B1(n_1227),
.B2(n_1186),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1254),
.A2(n_1248),
.B(n_1249),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1249),
.A2(n_1258),
.B(n_1195),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1208),
.A2(n_786),
.B(n_1113),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1290),
.Y(n_1421)
);

AO32x2_ASAP7_75t_L g1422 ( 
.A1(n_1262),
.A2(n_1300),
.A3(n_1022),
.B1(n_1177),
.B2(n_1159),
.Y(n_1422)
);

AO32x2_ASAP7_75t_L g1423 ( 
.A1(n_1262),
.A2(n_1300),
.A3(n_1022),
.B1(n_1177),
.B2(n_1159),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1290),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1180),
.B(n_984),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1180),
.A2(n_786),
.B(n_1174),
.C(n_636),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1149),
.A2(n_786),
.B(n_1113),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1246),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1149),
.A2(n_786),
.B(n_1113),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1246),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1187),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1180),
.A2(n_786),
.B(n_1174),
.C(n_636),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1187),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_SL g1434 ( 
.A1(n_1235),
.A2(n_911),
.B(n_786),
.C(n_636),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1187),
.B(n_935),
.Y(n_1435)
);

INVx8_ASAP7_75t_L g1436 ( 
.A(n_1278),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1180),
.A2(n_786),
.B(n_1174),
.C(n_636),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1149),
.A2(n_786),
.B(n_1113),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1290),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1240),
.A2(n_1153),
.B(n_1290),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1187),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1290),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1246),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1174),
.B(n_786),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_SL g1445 ( 
.A1(n_1150),
.A2(n_1057),
.B(n_1090),
.C(n_786),
.Y(n_1445)
);

AOI211x1_ASAP7_75t_L g1446 ( 
.A1(n_1174),
.A2(n_1014),
.B(n_927),
.C(n_786),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1243),
.Y(n_1447)
);

AO31x2_ASAP7_75t_L g1448 ( 
.A1(n_1240),
.A2(n_1312),
.A3(n_1262),
.B(n_1107),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1233),
.B(n_1048),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1246),
.Y(n_1450)
);

NOR2xp67_ASAP7_75t_SL g1451 ( 
.A(n_1278),
.B(n_960),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1246),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1187),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1246),
.Y(n_1454)
);

CKINVDCx11_ASAP7_75t_R g1455 ( 
.A(n_1270),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1290),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1155),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1149),
.A2(n_786),
.B(n_1113),
.Y(n_1458)
);

AOI221xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1260),
.A2(n_1046),
.B1(n_1024),
.B2(n_1014),
.C(n_1022),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1155),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1156),
.A2(n_786),
.B(n_1019),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1246),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1180),
.B(n_984),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1180),
.B(n_984),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1151),
.Y(n_1465)
);

A2O1A1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1180),
.A2(n_786),
.B(n_1174),
.C(n_636),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1149),
.A2(n_786),
.B(n_1113),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1180),
.A2(n_786),
.B1(n_1174),
.B2(n_992),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1187),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1290),
.Y(n_1470)
);

O2A1O1Ixp5_ASAP7_75t_L g1471 ( 
.A1(n_1240),
.A2(n_786),
.B(n_911),
.C(n_548),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1155),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_R g1473 ( 
.A(n_1243),
.B(n_781),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1233),
.B(n_1048),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1149),
.A2(n_786),
.B(n_1113),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1156),
.A2(n_786),
.B(n_1019),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1246),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1246),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1246),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1180),
.B(n_786),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1180),
.B(n_786),
.C(n_1174),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1278),
.Y(n_1482)
);

AO31x2_ASAP7_75t_L g1483 ( 
.A1(n_1240),
.A2(n_1312),
.A3(n_1262),
.B(n_1107),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1290),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_SL g1485 ( 
.A1(n_1150),
.A2(n_1057),
.B(n_1090),
.C(n_786),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1187),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1174),
.B(n_786),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1346),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1396),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1427),
.A2(n_1438),
.B(n_1429),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1433),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1444),
.A2(n_1487),
.B1(n_1406),
.B2(n_1411),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1349),
.Y(n_1493)
);

NAND2x1p5_ASAP7_75t_L g1494 ( 
.A(n_1388),
.B(n_1441),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1410),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1322),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1481),
.A2(n_1468),
.B1(n_1480),
.B2(n_1387),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1481),
.A2(n_1387),
.B1(n_1463),
.B2(n_1425),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1426),
.B(n_1432),
.Y(n_1499)
);

BUFx8_ASAP7_75t_L g1500 ( 
.A(n_1381),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1437),
.B(n_1466),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1386),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1356),
.A2(n_1411),
.B1(n_1395),
.B2(n_1461),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1464),
.A2(n_1316),
.B1(n_1417),
.B2(n_1395),
.Y(n_1504)
);

BUFx4f_ASAP7_75t_SL g1505 ( 
.A(n_1447),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1373),
.A2(n_1476),
.B1(n_1449),
.B2(n_1474),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1377),
.A2(n_1449),
.B1(n_1474),
.B2(n_1414),
.Y(n_1507)
);

INVx6_ASAP7_75t_L g1508 ( 
.A(n_1436),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1476),
.A2(n_1365),
.B1(n_1371),
.B2(n_1399),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1318),
.A2(n_1408),
.B1(n_1364),
.B2(n_1348),
.Y(n_1510)
);

BUFx4_ASAP7_75t_R g1511 ( 
.A(n_1473),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1397),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1352),
.Y(n_1513)
);

INVx8_ASAP7_75t_L g1514 ( 
.A(n_1388),
.Y(n_1514)
);

BUFx8_ASAP7_75t_SL g1515 ( 
.A(n_1345),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1360),
.A2(n_1446),
.B1(n_1413),
.B2(n_1319),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1408),
.A2(n_1399),
.B1(n_1353),
.B2(n_1419),
.Y(n_1517)
);

INVx4_ASAP7_75t_SL g1518 ( 
.A(n_1366),
.Y(n_1518)
);

CKINVDCx6p67_ASAP7_75t_R g1519 ( 
.A(n_1382),
.Y(n_1519)
);

INVx6_ASAP7_75t_L g1520 ( 
.A(n_1388),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1465),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1319),
.A2(n_1412),
.B1(n_1376),
.B2(n_1479),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1354),
.B(n_1385),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1410),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1414),
.A2(n_1400),
.B1(n_1405),
.B2(n_1459),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1431),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1469),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1331),
.A2(n_1420),
.B1(n_1354),
.B2(n_1367),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1368),
.A2(n_1324),
.B1(n_1334),
.B2(n_1361),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1428),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1430),
.A2(n_1443),
.B1(n_1478),
.B2(n_1477),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1357),
.Y(n_1532)
);

OAI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1370),
.A2(n_1369),
.B1(n_1361),
.B2(n_1435),
.Y(n_1533)
);

CKINVDCx11_ASAP7_75t_R g1534 ( 
.A(n_1441),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1358),
.A2(n_1459),
.B1(n_1359),
.B2(n_1363),
.Y(n_1535)
);

INVx6_ASAP7_75t_L g1536 ( 
.A(n_1337),
.Y(n_1536)
);

BUFx12f_ASAP7_75t_L g1537 ( 
.A(n_1347),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1434),
.B(n_1458),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1344),
.A2(n_1375),
.B1(n_1380),
.B2(n_1486),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1450),
.A2(n_1452),
.B1(n_1462),
.B2(n_1454),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1402),
.Y(n_1541)
);

CKINVDCx11_ASAP7_75t_R g1542 ( 
.A(n_1380),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1375),
.A2(n_1336),
.B1(n_1472),
.B2(n_1457),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1451),
.B(n_1337),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1460),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1372),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1366),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1398),
.A2(n_1320),
.B1(n_1416),
.B2(n_1392),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_L g1549 ( 
.A(n_1374),
.Y(n_1549)
);

CKINVDCx11_ASAP7_75t_R g1550 ( 
.A(n_1482),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1366),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1351),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1398),
.A2(n_1475),
.B1(n_1467),
.B2(n_1392),
.Y(n_1553)
);

CKINVDCx11_ASAP7_75t_R g1554 ( 
.A(n_1409),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1383),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1394),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1330),
.A2(n_1355),
.B1(n_1323),
.B2(n_1350),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1422),
.A2(n_1423),
.B1(n_1389),
.B2(n_1485),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1403),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1401),
.A2(n_1404),
.B1(n_1342),
.B2(n_1335),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1393),
.A2(n_1407),
.B1(n_1326),
.B2(n_1341),
.Y(n_1561)
);

INVx3_ASAP7_75t_SL g1562 ( 
.A(n_1440),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1394),
.Y(n_1563)
);

CKINVDCx11_ASAP7_75t_R g1564 ( 
.A(n_1391),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1384),
.B(n_1471),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1390),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1384),
.Y(n_1567)
);

BUFx8_ASAP7_75t_L g1568 ( 
.A(n_1422),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1418),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1445),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1384),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1422),
.A2(n_1423),
.B1(n_1328),
.B2(n_1315),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1423),
.A2(n_1378),
.B1(n_1340),
.B2(n_1325),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1415),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1321),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1415),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1415),
.B(n_1325),
.Y(n_1577)
);

CKINVDCx6p67_ASAP7_75t_R g1578 ( 
.A(n_1332),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1338),
.A2(n_1339),
.B1(n_1448),
.B2(n_1483),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1379),
.A2(n_1343),
.B1(n_1484),
.B2(n_1424),
.Y(n_1580)
);

INVx4_ASAP7_75t_L g1581 ( 
.A(n_1329),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1325),
.A2(n_1339),
.B1(n_1448),
.B2(n_1483),
.Y(n_1582)
);

BUFx8_ASAP7_75t_L g1583 ( 
.A(n_1339),
.Y(n_1583)
);

OAI22x1_ASAP7_75t_L g1584 ( 
.A1(n_1448),
.A2(n_1483),
.B1(n_1362),
.B2(n_1333),
.Y(n_1584)
);

BUFx5_ASAP7_75t_L g1585 ( 
.A(n_1329),
.Y(n_1585)
);

NAND2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1317),
.B(n_1439),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1362),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1362),
.A2(n_1333),
.B1(n_1421),
.B2(n_1442),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1333),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1327),
.A2(n_786),
.B1(n_1411),
.B2(n_802),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1456),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1470),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1427),
.A2(n_1438),
.B(n_1429),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1436),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1433),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1387),
.A2(n_802),
.B1(n_794),
.B2(n_786),
.Y(n_1599)
);

BUFx12f_ASAP7_75t_L g1600 ( 
.A(n_1455),
.Y(n_1600)
);

INVx6_ASAP7_75t_L g1601 ( 
.A(n_1436),
.Y(n_1601)
);

INVx6_ASAP7_75t_L g1602 ( 
.A(n_1436),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1397),
.Y(n_1605)
);

INVx6_ASAP7_75t_L g1606 ( 
.A(n_1436),
.Y(n_1606)
);

INVx6_ASAP7_75t_L g1607 ( 
.A(n_1436),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1356),
.A2(n_786),
.B1(n_1411),
.B2(n_1288),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1388),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1436),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1453),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1480),
.B(n_1444),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1396),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1433),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1396),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1356),
.A2(n_786),
.B1(n_1411),
.B2(n_1288),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1388),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_SL g1623 ( 
.A(n_1447),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1388),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1433),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1455),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1356),
.A2(n_786),
.B1(n_1411),
.B2(n_1288),
.Y(n_1627)
);

BUFx12f_ASAP7_75t_L g1628 ( 
.A(n_1455),
.Y(n_1628)
);

CKINVDCx11_ASAP7_75t_R g1629 ( 
.A(n_1455),
.Y(n_1629)
);

BUFx8_ASAP7_75t_SL g1630 ( 
.A(n_1345),
.Y(n_1630)
);

BUFx8_ASAP7_75t_SL g1631 ( 
.A(n_1345),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1353),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1346),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1481),
.A2(n_1180),
.B1(n_786),
.B2(n_1174),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1396),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1396),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1356),
.A2(n_786),
.B1(n_1411),
.B2(n_1288),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1480),
.B(n_1444),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1444),
.A2(n_802),
.B1(n_1180),
.B2(n_786),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1388),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1480),
.B(n_1444),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1411),
.A2(n_786),
.B1(n_802),
.B2(n_794),
.Y(n_1643)
);

OAI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1411),
.A2(n_786),
.B1(n_802),
.B2(n_794),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1547),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1564),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1488),
.Y(n_1647)
);

INVx5_ASAP7_75t_L g1648 ( 
.A(n_1574),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1587),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1555),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1551),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1563),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1556),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1492),
.B(n_1613),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1490),
.A2(n_1594),
.B(n_1588),
.Y(n_1655)
);

BUFx2_ASAP7_75t_SL g1656 ( 
.A(n_1623),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1493),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1502),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1494),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1523),
.B(n_1613),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1632),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1571),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1530),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1518),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1491),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1639),
.B(n_1642),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1518),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1548),
.B(n_1518),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1639),
.B(n_1642),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1567),
.Y(n_1670)
);

AOI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1538),
.A2(n_1553),
.B(n_1557),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1640),
.B(n_1593),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1576),
.Y(n_1673)
);

OAI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1608),
.A2(n_1627),
.B1(n_1638),
.B2(n_1619),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1584),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1565),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1548),
.B(n_1589),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1581),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1595),
.B(n_1598),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1514),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1554),
.Y(n_1681)
);

AND2x2_ASAP7_75t_SL g1682 ( 
.A(n_1568),
.B(n_1497),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1577),
.Y(n_1683)
);

AND2x2_ASAP7_75t_SL g1684 ( 
.A(n_1504),
.B(n_1603),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1577),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1585),
.Y(n_1686)
);

AO21x1_ASAP7_75t_L g1687 ( 
.A1(n_1503),
.A2(n_1557),
.B(n_1608),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1604),
.A2(n_1615),
.B(n_1611),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1585),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1585),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1634),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1541),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1514),
.Y(n_1693)
);

NOR3xp33_ASAP7_75t_L g1694 ( 
.A(n_1643),
.B(n_1644),
.C(n_1599),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1597),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1531),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1494),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1575),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1559),
.B(n_1507),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1503),
.A2(n_1627),
.B1(n_1638),
.B2(n_1619),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1531),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1540),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1612),
.Y(n_1703)
);

AO21x1_ASAP7_75t_SL g1704 ( 
.A1(n_1499),
.A2(n_1501),
.B(n_1517),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1540),
.Y(n_1705)
);

INVxp33_ASAP7_75t_L g1706 ( 
.A(n_1534),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1489),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1614),
.Y(n_1708)
);

AOI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1538),
.A2(n_1560),
.B(n_1588),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1569),
.B(n_1617),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1586),
.A2(n_1561),
.B(n_1580),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1583),
.Y(n_1712)
);

AO21x2_ASAP7_75t_L g1713 ( 
.A1(n_1561),
.A2(n_1560),
.B(n_1566),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1542),
.Y(n_1714)
);

AOI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1591),
.A2(n_1501),
.B(n_1499),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1579),
.B(n_1498),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1612),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1509),
.B(n_1582),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1583),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1509),
.B(n_1582),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1616),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1636),
.B(n_1637),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1525),
.B(n_1610),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1586),
.A2(n_1579),
.B(n_1570),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1592),
.B(n_1514),
.Y(n_1725)
);

AO21x1_ASAP7_75t_L g1726 ( 
.A1(n_1516),
.A2(n_1590),
.B(n_1522),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1496),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1513),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1532),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1605),
.B(n_1512),
.Y(n_1730)
);

OR2x6_ASAP7_75t_L g1731 ( 
.A(n_1544),
.B(n_1516),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1545),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1618),
.A2(n_1620),
.B(n_1635),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1599),
.A2(n_1622),
.B1(n_1633),
.B2(n_1535),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1528),
.A2(n_1510),
.B(n_1539),
.Y(n_1735)
);

AOI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1522),
.A2(n_1552),
.B(n_1578),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1562),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1526),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1526),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1526),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1529),
.B(n_1524),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1573),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1573),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1572),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1572),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1558),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1558),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1544),
.B(n_1520),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1625),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_SL g1750 ( 
.A1(n_1543),
.A2(n_1506),
.B(n_1596),
.Y(n_1750)
);

AO21x2_ASAP7_75t_L g1751 ( 
.A1(n_1533),
.A2(n_1535),
.B(n_1520),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1520),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1527),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1515),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1609),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1621),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1495),
.B(n_1641),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1621),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1624),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1624),
.Y(n_1760)
);

NAND2x1p5_ASAP7_75t_L g1761 ( 
.A(n_1549),
.B(n_1641),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1624),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1623),
.A2(n_1505),
.B1(n_1519),
.B2(n_1537),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1536),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1508),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1601),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1549),
.B(n_1602),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1521),
.B(n_1550),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1601),
.B(n_1606),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1546),
.B(n_1607),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1721),
.Y(n_1771)
);

OR2x6_ASAP7_75t_L g1772 ( 
.A(n_1731),
.B(n_1600),
.Y(n_1772)
);

NAND2x1p5_ASAP7_75t_L g1773 ( 
.A(n_1648),
.B(n_1511),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1700),
.A2(n_1626),
.B(n_1602),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1660),
.B(n_1606),
.Y(n_1775)
);

O2A1O1Ixp33_ASAP7_75t_SL g1776 ( 
.A1(n_1674),
.A2(n_1629),
.B(n_1500),
.C(n_1628),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1734),
.A2(n_1606),
.B1(n_1607),
.B2(n_1500),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1757),
.B(n_1630),
.Y(n_1778)
);

A2O1A1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1694),
.A2(n_1631),
.B(n_1733),
.C(n_1688),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1687),
.A2(n_1654),
.B1(n_1726),
.B2(n_1679),
.C(n_1672),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1677),
.B(n_1712),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1677),
.B(n_1712),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1660),
.B(n_1666),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1684),
.A2(n_1682),
.B(n_1698),
.C(n_1716),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1684),
.A2(n_1682),
.B1(n_1666),
.B2(n_1669),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1719),
.B(n_1698),
.Y(n_1786)
);

AO32x2_ASAP7_75t_L g1787 ( 
.A1(n_1659),
.A2(n_1697),
.A3(n_1676),
.B1(n_1742),
.B2(n_1743),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1665),
.B(n_1695),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1696),
.B(n_1701),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1702),
.B(n_1705),
.Y(n_1790)
);

A2O1A1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1716),
.A2(n_1720),
.B(n_1718),
.C(n_1668),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1687),
.A2(n_1726),
.B1(n_1699),
.B2(n_1731),
.Y(n_1792)
);

O2A1O1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1741),
.A2(n_1750),
.B(n_1731),
.C(n_1703),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1736),
.A2(n_1671),
.B(n_1735),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1648),
.B(n_1725),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1735),
.A2(n_1699),
.B(n_1655),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1731),
.B(n_1725),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1718),
.A2(n_1720),
.B(n_1699),
.C(n_1730),
.Y(n_1798)
);

NOR2x1_ASAP7_75t_SL g1799 ( 
.A(n_1748),
.B(n_1725),
.Y(n_1799)
);

AND2x2_ASAP7_75t_SL g1800 ( 
.A(n_1646),
.B(n_1735),
.Y(n_1800)
);

AOI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1715),
.A2(n_1709),
.B(n_1667),
.Y(n_1801)
);

AO32x2_ASAP7_75t_L g1802 ( 
.A1(n_1659),
.A2(n_1697),
.A3(n_1742),
.B1(n_1743),
.B2(n_1745),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1648),
.B(n_1725),
.Y(n_1803)
);

O2A1O1Ixp33_ASAP7_75t_SL g1804 ( 
.A1(n_1714),
.A2(n_1768),
.B(n_1706),
.C(n_1769),
.Y(n_1804)
);

OR2x6_ASAP7_75t_L g1805 ( 
.A(n_1748),
.B(n_1711),
.Y(n_1805)
);

A2O1A1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1744),
.A2(n_1745),
.B(n_1656),
.C(n_1723),
.Y(n_1806)
);

AO32x2_ASAP7_75t_L g1807 ( 
.A1(n_1744),
.A2(n_1675),
.A3(n_1746),
.B1(n_1747),
.B2(n_1673),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1717),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1646),
.A2(n_1747),
.B1(n_1746),
.B2(n_1661),
.Y(n_1809)
);

AO32x2_ASAP7_75t_L g1810 ( 
.A1(n_1675),
.A2(n_1673),
.A3(n_1652),
.B1(n_1704),
.B2(n_1685),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_R g1811 ( 
.A(n_1754),
.B(n_1646),
.Y(n_1811)
);

AOI21xp33_ASAP7_75t_L g1812 ( 
.A1(n_1751),
.A2(n_1750),
.B(n_1713),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1723),
.A2(n_1656),
.B1(n_1751),
.B2(n_1748),
.Y(n_1813)
);

AO32x2_ASAP7_75t_L g1814 ( 
.A1(n_1652),
.A2(n_1704),
.A3(n_1685),
.B1(n_1683),
.B2(n_1645),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1723),
.A2(n_1751),
.B1(n_1748),
.B2(n_1749),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1711),
.A2(n_1646),
.B(n_1753),
.C(n_1648),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1710),
.A2(n_1724),
.B(n_1722),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1646),
.A2(n_1753),
.B1(n_1681),
.B2(n_1692),
.Y(n_1818)
);

OA21x2_ASAP7_75t_L g1819 ( 
.A1(n_1686),
.A2(n_1690),
.B(n_1689),
.Y(n_1819)
);

OAI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1647),
.A2(n_1691),
.B(n_1663),
.C(n_1658),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1662),
.A2(n_1681),
.B(n_1739),
.C(n_1740),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1657),
.B(n_1650),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1650),
.B(n_1710),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1770),
.B(n_1754),
.Y(n_1824)
);

O2A1O1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1738),
.A2(n_1740),
.B(n_1761),
.C(n_1752),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1651),
.B(n_1737),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1770),
.B(n_1766),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1651),
.Y(n_1828)
);

NAND2x1_ASAP7_75t_L g1829 ( 
.A(n_1653),
.B(n_1678),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1670),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1727),
.B(n_1729),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1819),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1828),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1805),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1829),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1783),
.B(n_1713),
.Y(n_1836)
);

INVxp67_ASAP7_75t_SL g1837 ( 
.A(n_1826),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1780),
.A2(n_1752),
.B1(n_1764),
.B2(n_1765),
.Y(n_1838)
);

INVx4_ASAP7_75t_L g1839 ( 
.A(n_1772),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1785),
.A2(n_1680),
.B1(n_1693),
.B2(n_1708),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1830),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1805),
.Y(n_1842)
);

AOI222xp33_ASAP7_75t_L g1843 ( 
.A1(n_1780),
.A2(n_1763),
.B1(n_1707),
.B2(n_1732),
.C1(n_1728),
.C2(n_1729),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1831),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1814),
.B(n_1664),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1814),
.B(n_1807),
.Y(n_1846)
);

AO22x1_ASAP7_75t_L g1847 ( 
.A1(n_1818),
.A2(n_1680),
.B1(n_1693),
.B2(n_1758),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1822),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1807),
.B(n_1649),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1822),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1796),
.B(n_1760),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1826),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1779),
.B(n_1680),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1796),
.B(n_1759),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1787),
.B(n_1759),
.Y(n_1855)
);

OAI221xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1784),
.A2(n_1792),
.B1(n_1791),
.B2(n_1798),
.C(n_1813),
.Y(n_1856)
);

NOR2xp67_ASAP7_75t_L g1857 ( 
.A(n_1820),
.B(n_1762),
.Y(n_1857)
);

INVx4_ASAP7_75t_R g1858 ( 
.A(n_1786),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1787),
.B(n_1756),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1787),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1802),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1802),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1810),
.B(n_1755),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1789),
.B(n_1755),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1810),
.B(n_1781),
.Y(n_1865)
);

NOR2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1795),
.B(n_1803),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1802),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1808),
.Y(n_1868)
);

OAI33xp33_ASAP7_75t_L g1869 ( 
.A1(n_1861),
.A2(n_1809),
.A3(n_1862),
.B1(n_1867),
.B2(n_1818),
.B3(n_1864),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1833),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1834),
.Y(n_1871)
);

OAI21xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1857),
.A2(n_1800),
.B(n_1815),
.Y(n_1872)
);

BUFx8_ASAP7_75t_L g1873 ( 
.A(n_1834),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1833),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1834),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1841),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1841),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1860),
.B(n_1836),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1837),
.B(n_1794),
.Y(n_1879)
);

NAND2xp67_ASAP7_75t_L g1880 ( 
.A(n_1851),
.B(n_1778),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1832),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1832),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1837),
.B(n_1790),
.Y(n_1883)
);

O2A1O1Ixp5_ASAP7_75t_L g1884 ( 
.A1(n_1856),
.A2(n_1812),
.B(n_1816),
.C(n_1809),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1846),
.B(n_1805),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1846),
.B(n_1817),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1857),
.B(n_1793),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1845),
.B(n_1865),
.Y(n_1888)
);

INVxp67_ASAP7_75t_SL g1889 ( 
.A(n_1849),
.Y(n_1889)
);

OAI33xp33_ASAP7_75t_L g1890 ( 
.A1(n_1861),
.A2(n_1771),
.A3(n_1777),
.B1(n_1775),
.B2(n_1825),
.B3(n_1823),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1852),
.B(n_1788),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1845),
.B(n_1801),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1865),
.B(n_1797),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1866),
.B(n_1799),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1855),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1836),
.B(n_1775),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1834),
.B(n_1797),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1855),
.Y(n_1898)
);

OAI221xp5_ASAP7_75t_L g1899 ( 
.A1(n_1856),
.A2(n_1774),
.B1(n_1777),
.B2(n_1776),
.C(n_1806),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1855),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1835),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1838),
.A2(n_1774),
.B1(n_1804),
.B2(n_1782),
.C(n_1827),
.Y(n_1902)
);

NOR3xp33_ASAP7_75t_SL g1903 ( 
.A(n_1899),
.B(n_1853),
.C(n_1824),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1887),
.B(n_1839),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1870),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1887),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1895),
.B(n_1898),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1870),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1894),
.B(n_1834),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1874),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1874),
.Y(n_1911)
);

NOR4xp25_ASAP7_75t_SL g1912 ( 
.A(n_1899),
.B(n_1821),
.C(n_1867),
.D(n_1847),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1895),
.B(n_1859),
.Y(n_1913)
);

NAND4xp25_ASAP7_75t_L g1914 ( 
.A(n_1884),
.B(n_1843),
.C(n_1840),
.D(n_1839),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1900),
.B(n_1863),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1879),
.B(n_1844),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1876),
.Y(n_1917)
);

NAND2x1_ASAP7_75t_L g1918 ( 
.A(n_1894),
.B(n_1858),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1881),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1896),
.B(n_1883),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1896),
.B(n_1848),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1876),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1877),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1883),
.B(n_1848),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1879),
.B(n_1850),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1873),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1889),
.B(n_1863),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1881),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1894),
.B(n_1842),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1901),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1886),
.B(n_1851),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1886),
.B(n_1851),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1886),
.B(n_1854),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1894),
.B(n_1842),
.Y(n_1934)
);

XOR2x2_ASAP7_75t_L g1935 ( 
.A(n_1902),
.B(n_1847),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1909),
.B(n_1885),
.Y(n_1936)
);

NAND2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1904),
.B(n_1871),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1906),
.B(n_1880),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1909),
.B(n_1929),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1909),
.B(n_1885),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1909),
.B(n_1885),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1906),
.B(n_1880),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1904),
.B(n_1880),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1920),
.B(n_1878),
.Y(n_1944)
);

OR2x6_ASAP7_75t_L g1945 ( 
.A(n_1926),
.B(n_1772),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1926),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1920),
.B(n_1925),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1909),
.B(n_1894),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1925),
.B(n_1892),
.Y(n_1949)
);

INVx3_ASAP7_75t_L g1950 ( 
.A(n_1918),
.Y(n_1950)
);

O2A1O1Ixp33_ASAP7_75t_SL g1951 ( 
.A1(n_1918),
.A2(n_1902),
.B(n_1901),
.C(n_1868),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1905),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1924),
.B(n_1892),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1929),
.B(n_1888),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1907),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1905),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1919),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1908),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1929),
.B(n_1897),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1919),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1908),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1929),
.B(n_1888),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1935),
.B(n_1868),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1929),
.B(n_1888),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1934),
.B(n_1893),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1910),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1924),
.B(n_1892),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1935),
.B(n_1891),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1910),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1907),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1934),
.B(n_1893),
.Y(n_1971)
);

NOR2xp67_ASAP7_75t_SL g1972 ( 
.A(n_1914),
.B(n_1839),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1934),
.B(n_1893),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1921),
.B(n_1882),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1935),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1911),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1935),
.B(n_1891),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1911),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1934),
.B(n_1931),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1917),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1917),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1907),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1946),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1947),
.B(n_1916),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1950),
.B(n_1934),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1954),
.B(n_1931),
.Y(n_1986)
);

INVx2_ASAP7_75t_SL g1987 ( 
.A(n_1950),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1954),
.B(n_1931),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1962),
.B(n_1932),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1975),
.B(n_1921),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1968),
.B(n_1977),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1962),
.B(n_1932),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1964),
.B(n_1932),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1963),
.B(n_1927),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1964),
.B(n_1933),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1965),
.B(n_1933),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1957),
.B(n_1960),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1946),
.B(n_1927),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1938),
.B(n_1927),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1952),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1952),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1955),
.B(n_1933),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1956),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1965),
.B(n_1918),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1955),
.B(n_1915),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1937),
.B(n_1913),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1971),
.B(n_1915),
.Y(n_2007)
);

INVx2_ASAP7_75t_SL g2008 ( 
.A(n_1950),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1937),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1971),
.B(n_1915),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1972),
.B(n_1926),
.Y(n_2011)
);

AND2x4_ASAP7_75t_SL g2012 ( 
.A(n_1945),
.B(n_1903),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1973),
.B(n_1913),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1955),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1970),
.B(n_1928),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1970),
.B(n_1928),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1956),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1973),
.B(n_1913),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1970),
.B(n_1922),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1982),
.B(n_1922),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1982),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1982),
.B(n_1923),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1947),
.B(n_1923),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1987),
.Y(n_2024)
);

OAI21xp5_ASAP7_75t_SL g2025 ( 
.A1(n_1991),
.A2(n_1914),
.B(n_1937),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2004),
.B(n_1939),
.Y(n_2026)
);

AOI21xp33_ASAP7_75t_SL g2027 ( 
.A1(n_2011),
.A2(n_1943),
.B(n_1972),
.Y(n_2027)
);

OAI221xp5_ASAP7_75t_L g2028 ( 
.A1(n_1990),
.A2(n_1903),
.B1(n_1951),
.B2(n_1945),
.C(n_1884),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1983),
.B(n_1942),
.Y(n_2029)
);

AOI31xp33_ASAP7_75t_L g2030 ( 
.A1(n_1983),
.A2(n_1773),
.A3(n_1890),
.B(n_1872),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2000),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_2012),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_2012),
.B(n_1959),
.Y(n_2033)
);

INVxp67_ASAP7_75t_L g2034 ( 
.A(n_1997),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1987),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1990),
.B(n_1979),
.Y(n_2036)
);

AOI33xp33_ASAP7_75t_L g2037 ( 
.A1(n_2012),
.A2(n_1912),
.A3(n_1979),
.B1(n_1939),
.B2(n_1959),
.B3(n_1969),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2004),
.B(n_1936),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1997),
.B(n_1936),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2000),
.Y(n_2040)
);

INVxp33_ASAP7_75t_L g2041 ( 
.A(n_1994),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1985),
.B(n_1940),
.Y(n_2042)
);

NOR3xp33_ASAP7_75t_L g2043 ( 
.A(n_1999),
.B(n_1994),
.C(n_1998),
.Y(n_2043)
);

NOR4xp25_ASAP7_75t_L g2044 ( 
.A(n_2009),
.B(n_1872),
.C(n_1949),
.D(n_1974),
.Y(n_2044)
);

INVxp67_ASAP7_75t_L g2045 ( 
.A(n_1998),
.Y(n_2045)
);

XNOR2xp5_ASAP7_75t_L g2046 ( 
.A(n_1999),
.B(n_1773),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1985),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1996),
.B(n_1940),
.Y(n_2048)
);

AOI21xp33_ASAP7_75t_SL g2049 ( 
.A1(n_1987),
.A2(n_1945),
.B(n_1912),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1996),
.B(n_1941),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_2014),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2001),
.Y(n_2052)
);

OAI322xp33_ASAP7_75t_L g2053 ( 
.A1(n_2034),
.A2(n_2045),
.A3(n_2028),
.B1(n_2049),
.B2(n_2029),
.C1(n_2027),
.C2(n_2039),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_2043),
.A2(n_1890),
.B1(n_2009),
.B2(n_1945),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2042),
.B(n_2038),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_2025),
.A2(n_1945),
.B(n_2015),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2051),
.Y(n_2057)
);

O2A1O1Ixp33_ASAP7_75t_SL g2058 ( 
.A1(n_2049),
.A2(n_2008),
.B(n_2014),
.C(n_1950),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2025),
.A2(n_2032),
.B1(n_2033),
.B2(n_2042),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2038),
.B(n_1941),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_2032),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2026),
.B(n_1985),
.Y(n_2062)
);

AOI322xp5_ASAP7_75t_L g2063 ( 
.A1(n_2036),
.A2(n_2006),
.A3(n_2010),
.B1(n_2007),
.B2(n_2013),
.C1(n_2018),
.C2(n_1988),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_SL g2064 ( 
.A(n_2037),
.B(n_2006),
.C(n_2002),
.D(n_1988),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2031),
.Y(n_2065)
);

AND2x2_ASAP7_75t_SL g2066 ( 
.A(n_2044),
.B(n_1985),
.Y(n_2066)
);

A2O1A1Ixp33_ASAP7_75t_SL g2067 ( 
.A1(n_2024),
.A2(n_2001),
.B(n_2017),
.C(n_2003),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2031),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2026),
.B(n_1959),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_2030),
.A2(n_2016),
.B(n_2015),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2041),
.B(n_1959),
.Y(n_2071)
);

O2A1O1Ixp33_ASAP7_75t_L g2072 ( 
.A1(n_2027),
.A2(n_2008),
.B(n_2016),
.C(n_2006),
.Y(n_2072)
);

AOI21xp33_ASAP7_75t_L g2073 ( 
.A1(n_2030),
.A2(n_2008),
.B(n_1984),
.Y(n_2073)
);

OAI32xp33_ASAP7_75t_L g2074 ( 
.A1(n_2044),
.A2(n_2005),
.A3(n_2002),
.B1(n_1984),
.B2(n_2023),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2047),
.Y(n_2075)
);

OAI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_2059),
.A2(n_2047),
.B1(n_2050),
.B2(n_2048),
.Y(n_2076)
);

XNOR2x2_ASAP7_75t_L g2077 ( 
.A(n_2061),
.B(n_2040),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2062),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2066),
.B(n_2046),
.Y(n_2079)
);

XNOR2xp5_ASAP7_75t_L g2080 ( 
.A(n_2055),
.B(n_2046),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2066),
.B(n_2075),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_2075),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2064),
.A2(n_1869),
.B1(n_1948),
.B2(n_2007),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2057),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_2053),
.A2(n_2052),
.B1(n_2040),
.B2(n_1869),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2062),
.B(n_2024),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2065),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2068),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2060),
.B(n_2010),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2071),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2054),
.A2(n_2018),
.B1(n_2013),
.B2(n_1992),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_2056),
.Y(n_2092)
);

NAND3xp33_ASAP7_75t_SL g2093 ( 
.A(n_2079),
.B(n_2072),
.C(n_2054),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2081),
.B(n_2071),
.Y(n_2094)
);

O2A1O1Ixp33_ASAP7_75t_L g2095 ( 
.A1(n_2076),
.A2(n_2067),
.B(n_2058),
.C(n_2073),
.Y(n_2095)
);

NOR3xp33_ASAP7_75t_L g2096 ( 
.A(n_2092),
.B(n_2067),
.C(n_2058),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2082),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2085),
.A2(n_2070),
.B1(n_2052),
.B2(n_2035),
.Y(n_2098)
);

AOI211xp5_ASAP7_75t_L g2099 ( 
.A1(n_2091),
.A2(n_2074),
.B(n_2069),
.C(n_2035),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2077),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2078),
.B(n_2063),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2086),
.B(n_1988),
.Y(n_2102)
);

NAND3xp33_ASAP7_75t_L g2103 ( 
.A(n_2085),
.B(n_2017),
.C(n_2003),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2086),
.B(n_1992),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_2092),
.B(n_2080),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2078),
.B(n_1992),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2090),
.B(n_1986),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2102),
.Y(n_2108)
);

AOI21xp33_ASAP7_75t_L g2109 ( 
.A1(n_2095),
.A2(n_2084),
.B(n_2087),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2097),
.B(n_2089),
.Y(n_2110)
);

OAI211xp5_ASAP7_75t_L g2111 ( 
.A1(n_2100),
.A2(n_2077),
.B(n_2083),
.C(n_2088),
.Y(n_2111)
);

OAI211xp5_ASAP7_75t_SL g2112 ( 
.A1(n_2105),
.A2(n_2021),
.B(n_2005),
.C(n_2023),
.Y(n_2112)
);

OAI21xp33_ASAP7_75t_SL g2113 ( 
.A1(n_2098),
.A2(n_1989),
.B(n_1986),
.Y(n_2113)
);

A2O1A1Ixp33_ASAP7_75t_L g2114 ( 
.A1(n_2096),
.A2(n_2021),
.B(n_1948),
.C(n_1989),
.Y(n_2114)
);

NAND4xp25_ASAP7_75t_L g2115 ( 
.A(n_2101),
.B(n_2021),
.C(n_1993),
.D(n_1995),
.Y(n_2115)
);

AOI221xp5_ASAP7_75t_L g2116 ( 
.A1(n_2111),
.A2(n_2098),
.B1(n_2093),
.B2(n_2103),
.C(n_2099),
.Y(n_2116)
);

OAI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2114),
.A2(n_2094),
.B1(n_2104),
.B2(n_2106),
.Y(n_2117)
);

AOI221xp5_ASAP7_75t_L g2118 ( 
.A1(n_2109),
.A2(n_2107),
.B1(n_1995),
.B2(n_1993),
.C(n_2019),
.Y(n_2118)
);

BUFx6f_ASAP7_75t_L g2119 ( 
.A(n_2110),
.Y(n_2119)
);

AOI22x1_ASAP7_75t_L g2120 ( 
.A1(n_2108),
.A2(n_1930),
.B1(n_1944),
.B2(n_1761),
.Y(n_2120)
);

OAI221xp5_ASAP7_75t_SL g2121 ( 
.A1(n_2113),
.A2(n_2022),
.B1(n_2020),
.B2(n_2019),
.C(n_1944),
.Y(n_2121)
);

AOI211xp5_ASAP7_75t_L g2122 ( 
.A1(n_2112),
.A2(n_1811),
.B(n_2020),
.C(n_2022),
.Y(n_2122)
);

INVxp33_ASAP7_75t_SL g2123 ( 
.A(n_2115),
.Y(n_2123)
);

NAND4xp25_ASAP7_75t_L g2124 ( 
.A(n_2111),
.B(n_1839),
.C(n_1843),
.D(n_1875),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2119),
.Y(n_2125)
);

NAND2x1p5_ASAP7_75t_SL g2126 ( 
.A(n_2120),
.B(n_2123),
.Y(n_2126)
);

OAI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2116),
.A2(n_1949),
.B(n_1953),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_2117),
.B(n_2119),
.Y(n_2128)
);

XNOR2x1_ASAP7_75t_L g2129 ( 
.A(n_2118),
.B(n_1772),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_2122),
.A2(n_1967),
.B1(n_1953),
.B2(n_1978),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2124),
.Y(n_2131)
);

OAI221xp5_ASAP7_75t_L g2132 ( 
.A1(n_2127),
.A2(n_2121),
.B1(n_1967),
.B2(n_1974),
.C(n_1875),
.Y(n_2132)
);

NOR2x1_ASAP7_75t_L g2133 ( 
.A(n_2128),
.B(n_1958),
.Y(n_2133)
);

AOI22x1_ASAP7_75t_L g2134 ( 
.A1(n_2125),
.A2(n_1930),
.B1(n_1980),
.B2(n_1978),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2134),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2135),
.A2(n_2132),
.B1(n_2131),
.B2(n_2129),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_2136),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2136),
.Y(n_2138)
);

AOI22x1_ASAP7_75t_L g2139 ( 
.A1(n_2137),
.A2(n_2135),
.B1(n_2126),
.B2(n_2133),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2137),
.B(n_2130),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2139),
.Y(n_2141)
);

OAI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_2140),
.A2(n_2138),
.B(n_2137),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2142),
.Y(n_2143)
);

OAI21xp5_ASAP7_75t_SL g2144 ( 
.A1(n_2143),
.A2(n_2141),
.B(n_1761),
.Y(n_2144)
);

XNOR2xp5_ASAP7_75t_L g2145 ( 
.A(n_2144),
.B(n_1767),
.Y(n_2145)
);

OAI221xp5_ASAP7_75t_L g2146 ( 
.A1(n_2145),
.A2(n_1981),
.B1(n_1958),
.B2(n_1961),
.C(n_1980),
.Y(n_2146)
);

AOI211xp5_ASAP7_75t_L g2147 ( 
.A1(n_2146),
.A2(n_1981),
.B(n_1966),
.C(n_1976),
.Y(n_2147)
);


endmodule