module fake_jpeg_4108_n_177 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_20),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_2),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_21),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_49),
.B1(n_17),
.B2(n_16),
.Y(n_63)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_52),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_14),
.B(n_18),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_51),
.B(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_15),
.B1(n_19),
.B2(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_27),
.A2(n_15),
.B1(n_19),
.B2(n_17),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_21),
.B(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_57),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_21),
.B(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_65),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_35),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_33),
.B1(n_15),
.B2(n_16),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_16),
.B1(n_24),
.B2(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_67),
.B1(n_68),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_44),
.B1(n_38),
.B2(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_64),
.B1(n_62),
.B2(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_81),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_84),
.B(n_81),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_30),
.B(n_35),
.C(n_40),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_53),
.B1(n_66),
.B2(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_36),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_28),
.B(n_29),
.C(n_23),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_94),
.Y(n_115)
);

AO221x1_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_66),
.B1(n_64),
.B2(n_30),
.C(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_95),
.B1(n_78),
.B2(n_83),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_68),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_97),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_99),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_35),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_79),
.B(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_82),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_105),
.B(n_39),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_77),
.B(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_80),
.B1(n_82),
.B2(n_73),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_113),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_80),
.B1(n_85),
.B2(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_80),
.C(n_71),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_117),
.C(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_39),
.C(n_30),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_119),
.C(n_122),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_112),
.C(n_109),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_93),
.C(n_98),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_97),
.C(n_95),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_117),
.C(n_103),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_72),
.Y(n_138)
);

OA21x2_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_86),
.B(n_100),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_128),
.A3(n_113),
.B1(n_106),
.B2(n_116),
.C(n_108),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_89),
.C(n_92),
.Y(n_128)
);

OAI21x1_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_30),
.B(n_72),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_72),
.B(n_108),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_131),
.A2(n_25),
.B(n_22),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_139),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_30),
.C(n_70),
.Y(n_139)
);

OA21x2_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_110),
.B(n_70),
.Y(n_140)
);

AOI31xp67_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_25),
.A3(n_22),
.B(n_4),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_110),
.C(n_25),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_143),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_124),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_25),
.C(n_22),
.Y(n_143)
);

OAI21x1_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_120),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_148),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_120),
.B1(n_125),
.B2(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_2),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_160),
.B(n_8),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_3),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_159),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_7),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_5),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_9),
.B(n_11),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_145),
.B1(n_146),
.B2(n_10),
.C(n_11),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_159),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_166),
.B(n_157),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_170),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_12),
.CON(n_171),
.SN(n_171)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_167),
.C(n_171),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);


endmodule