module fake_jpeg_1936_n_535 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_535);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_417;
wire n_362;
wire n_142;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_45),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_48),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_49),
.Y(n_145)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_50),
.Y(n_109)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_52),
.Y(n_112)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_58),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_13),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_61),
.Y(n_116)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_82),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_69),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_13),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_94),
.B(n_31),
.C(n_58),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_41),
.B(n_30),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

BUFx2_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_95),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_21),
.B(n_0),
.CON(n_94),
.SN(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_97),
.Y(n_130)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_99),
.Y(n_157)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_43),
.B1(n_31),
.B2(n_30),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_101),
.A2(n_35),
.B1(n_25),
.B2(n_16),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_19),
.B1(n_18),
.B2(n_42),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_106),
.A2(n_89),
.B1(n_113),
.B2(n_117),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_111),
.B(n_114),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_51),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_123),
.B(n_159),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_17),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_126),
.B(n_153),
.Y(n_209)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_37),
.B1(n_23),
.B2(n_25),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_131),
.A2(n_42),
.B1(n_23),
.B2(n_37),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_34),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_54),
.B(n_34),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_29),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_158),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_53),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_65),
.B(n_42),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_35),
.C(n_95),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_48),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_67),
.B(n_29),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_107),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_176),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_101),
.A2(n_74),
.B1(n_76),
.B2(n_93),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_106),
.B1(n_125),
.B2(n_148),
.Y(n_215)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_165),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_127),
.A2(n_79),
.B1(n_92),
.B2(n_77),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_166),
.A2(n_182),
.B1(n_107),
.B2(n_128),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_SL g227 ( 
.A1(n_173),
.A2(n_181),
.B(n_189),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_183),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_127),
.A2(n_19),
.B1(n_42),
.B2(n_18),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_129),
.A2(n_81),
.B1(n_84),
.B2(n_46),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_185),
.Y(n_223)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_191),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_19),
.B1(n_18),
.B2(n_42),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_157),
.Y(n_234)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_197),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_152),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_204),
.B(n_208),
.Y(n_236)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx6p67_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_200),
.A2(n_173),
.B1(n_189),
.B2(n_164),
.Y(n_216)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_129),
.B(n_126),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_157),
.B1(n_140),
.B2(n_160),
.Y(n_217)
);

BUFx12_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_215),
.A2(n_221),
.B1(n_226),
.B2(n_178),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_216),
.A2(n_166),
.B1(n_182),
.B2(n_190),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_154),
.C(n_115),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_209),
.C(n_167),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_149),
.B1(n_147),
.B2(n_136),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_151),
.B1(n_150),
.B2(n_128),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_231),
.B1(n_203),
.B2(n_177),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_172),
.A2(n_155),
.B1(n_146),
.B2(n_133),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_208),
.B(n_131),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_181),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_88),
.B(n_59),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_199),
.B(n_162),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_245),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_124),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_215),
.A2(n_196),
.B1(n_174),
.B2(n_171),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_246),
.A2(n_255),
.B(n_260),
.Y(n_297)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_242),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_253),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_220),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_258),
.C(n_267),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_190),
.B(n_196),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_211),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_230),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_262),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_168),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_259),
.B(n_263),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_138),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_231),
.B1(n_229),
.B2(n_218),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_198),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_133),
.B1(n_121),
.B2(n_179),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_269),
.B1(n_228),
.B2(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_134),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_230),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_210),
.A2(n_232),
.B(n_222),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_226),
.B(n_218),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_275),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_276),
.A2(n_278),
.B1(n_304),
.B2(n_305),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_281),
.A2(n_302),
.B(n_263),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_294),
.Y(n_309)
);

XOR2x2_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_221),
.Y(n_290)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_256),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_229),
.B1(n_223),
.B2(n_244),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_291),
.A2(n_295),
.B1(n_248),
.B2(n_254),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_250),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_249),
.A2(n_218),
.B1(n_223),
.B2(n_238),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_244),
.C(n_235),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_301),
.C(n_257),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_243),
.C(n_224),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_274),
.A2(n_218),
.B(n_224),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_255),
.A2(n_155),
.B1(n_186),
.B2(n_121),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_246),
.A2(n_237),
.B1(n_238),
.B2(n_219),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_260),
.B(n_252),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_306),
.A2(n_319),
.B(n_328),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_290),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_286),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_336),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_260),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_310),
.A2(n_322),
.B(n_329),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_253),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_270),
.C(n_257),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_315),
.C(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_293),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_326),
.B1(n_333),
.B2(n_288),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_257),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_280),
.B(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_260),
.B(n_268),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_258),
.C(n_256),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_337),
.Y(n_346)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_286),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_271),
.Y(n_327)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_284),
.A2(n_252),
.B(n_263),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_264),
.B(n_273),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_302),
.A2(n_259),
.B(n_247),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_218),
.B(n_266),
.Y(n_369)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_287),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_336),
.B1(n_296),
.B2(n_318),
.Y(n_339)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_335),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_285),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_275),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_349),
.B1(n_352),
.B2(n_356),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_331),
.A2(n_291),
.B1(n_292),
.B2(n_294),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_309),
.B1(n_320),
.B2(n_328),
.Y(n_372)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_334),
.A2(n_276),
.B1(n_304),
.B2(n_296),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_326),
.B(n_285),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_350),
.B(n_355),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_308),
.A2(n_305),
.B1(n_289),
.B2(n_292),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_301),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_358),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g355 ( 
.A(n_312),
.B(n_300),
.CI(n_301),
.CON(n_355),
.SN(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_314),
.A2(n_289),
.B1(n_297),
.B2(n_278),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_300),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_364),
.C(n_368),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_306),
.A2(n_287),
.B1(n_290),
.B2(n_295),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_362),
.A2(n_356),
.B1(n_349),
.B2(n_340),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_315),
.B(n_225),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_316),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_366),
.B(n_311),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_266),
.C(n_243),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_367),
.B(n_309),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_371),
.B(n_388),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_372),
.A2(n_374),
.B1(n_330),
.B2(n_310),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_339),
.B1(n_351),
.B2(n_340),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_327),
.Y(n_375)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_344),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_378),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_338),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_369),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_380),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_381),
.A2(n_393),
.B1(n_379),
.B2(n_390),
.Y(n_415)
);

NOR4xp25_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_335),
.C(n_332),
.D(n_337),
.Y(n_383)
);

AOI21xp33_ASAP7_75t_L g405 ( 
.A1(n_383),
.A2(n_389),
.B(n_319),
.Y(n_405)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_307),
.C(n_312),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_359),
.C(n_364),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_357),
.B(n_324),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_306),
.B(n_322),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_352),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_390),
.B(n_392),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_342),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_362),
.A2(n_331),
.B1(n_310),
.B2(n_330),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_341),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_310),
.Y(n_395)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_396),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_353),
.B(n_266),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_397),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_324),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_399),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_423),
.C(n_384),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_368),
.C(n_307),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_410),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_329),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_372),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_376),
.C(n_395),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_355),
.C(n_346),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_411),
.B(n_416),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_415),
.A2(n_417),
.B1(n_425),
.B2(n_396),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_355),
.C(n_313),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_381),
.A2(n_365),
.B1(n_363),
.B2(n_361),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_374),
.B(n_325),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_393),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_321),
.C(n_317),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_382),
.A2(n_238),
.B1(n_219),
.B2(n_240),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_425),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_373),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_431),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_373),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_407),
.A2(n_377),
.B1(n_382),
.B2(n_378),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_434),
.A2(n_449),
.B1(n_184),
.B2(n_207),
.Y(n_470)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_422),
.Y(n_435)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_437),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_385),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_446),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_380),
.C(n_387),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_443),
.C(n_414),
.Y(n_451)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_375),
.B1(n_389),
.B2(n_387),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_444),
.B1(n_402),
.B2(n_412),
.Y(n_461)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_423),
.C(n_408),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_394),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_419),
.B(n_398),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_448),
.Y(n_459)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_451),
.B(n_457),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_428),
.A2(n_404),
.B(n_409),
.Y(n_453)
);

AOI21x1_ASAP7_75t_SL g474 ( 
.A1(n_453),
.A2(n_437),
.B(n_427),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_438),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_466),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_418),
.C(n_400),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_433),
.A2(n_432),
.B(n_414),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_463),
.B(n_465),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_443),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_432),
.A2(n_413),
.B(n_426),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_441),
.A2(n_424),
.B1(n_237),
.B2(n_219),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_467),
.A2(n_468),
.B1(n_436),
.B2(n_446),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_431),
.A2(n_237),
.B1(n_240),
.B2(n_225),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_240),
.C(n_180),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_213),
.C(n_142),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_13),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_453),
.A2(n_213),
.B(n_214),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_476),
.A2(n_477),
.B(n_483),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_461),
.A2(n_452),
.B(n_451),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_478),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_214),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_482),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_214),
.C(n_213),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_450),
.A2(n_156),
.B(n_194),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_464),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_485),
.Y(n_490)
);

NAND2x1_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_194),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_25),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_487),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_161),
.C(n_156),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_161),
.C(n_156),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_469),
.C(n_99),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_472),
.A2(n_467),
.B1(n_459),
.B2(n_456),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_494),
.A2(n_501),
.B1(n_0),
.B2(n_1),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_471),
.A2(n_462),
.B1(n_466),
.B2(n_468),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_497),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_502),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_45),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_499),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_9),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_9),
.B1(n_14),
.B2(n_2),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_14),
.C(n_1),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_491),
.A2(n_485),
.B(n_475),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_503),
.A2(n_504),
.B(n_507),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_474),
.B(n_480),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_482),
.C(n_487),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_510),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_500),
.A2(n_488),
.B(n_478),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_14),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_511),
.B(n_2),
.Y(n_521)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_494),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_493),
.A2(n_14),
.B(n_9),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_496),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_493),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_514),
.B(n_515),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_492),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_505),
.A2(n_489),
.B(n_502),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_517),
.A2(n_521),
.B(n_2),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_519),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_0),
.C(n_1),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_523),
.A2(n_524),
.B(n_526),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_3),
.C(n_4),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_519),
.C(n_4),
.Y(n_526)
);

OAI311xp33_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.C1(n_6),
.Y(n_527)
);

AOI322xp5_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_333),
.C1(n_316),
.C2(n_311),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_522),
.A2(n_3),
.B(n_5),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_6),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_530),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_529),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_531),
.B(n_7),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_6),
.C(n_7),
.Y(n_535)
);


endmodule