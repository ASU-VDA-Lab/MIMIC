module fake_jpeg_19805_n_318 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_62),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_34),
.B1(n_29),
.B2(n_23),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_59),
.B1(n_38),
.B2(n_25),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_34),
.B1(n_18),
.B2(n_21),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_35),
.B1(n_27),
.B2(n_23),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_34),
.B1(n_29),
.B2(n_23),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_25),
.B1(n_20),
.B2(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_35),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_53),
.B1(n_49),
.B2(n_64),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_35),
.B(n_32),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_72),
.A2(n_78),
.B1(n_87),
.B2(n_90),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_45),
.C(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_42),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_89),
.Y(n_103)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_31),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_24),
.B1(n_30),
.B2(n_33),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_25),
.B(n_24),
.C(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_47),
.B(n_22),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_30),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_24),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_92),
.B(n_88),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_56),
.C(n_65),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_78),
.C(n_48),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

BUFx16f_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_19),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_93),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_65),
.B1(n_20),
.B2(n_26),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_77),
.B1(n_84),
.B2(n_79),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_17),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_79),
.B(n_67),
.C(n_89),
.D(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_72),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_70),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_129),
.B(n_130),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_72),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_133),
.A2(n_140),
.B(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_143),
.B1(n_151),
.B2(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_76),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_144),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_88),
.B(n_95),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_111),
.B(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_68),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_150),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_68),
.B1(n_85),
.B2(n_94),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_73),
.C(n_85),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_102),
.A2(n_96),
.B(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_109),
.B(n_73),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_100),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_71),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_73),
.B1(n_71),
.B2(n_80),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_80),
.C(n_26),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_120),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_17),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_111),
.B(n_113),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_171),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_159),
.A2(n_118),
.B1(n_16),
.B2(n_15),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_168),
.B1(n_170),
.B2(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_188),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_169),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_130),
.B(n_137),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_165),
.A2(n_183),
.B(n_1),
.C(n_2),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_127),
.A2(n_121),
.B1(n_123),
.B2(n_97),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_121),
.B1(n_97),
.B2(n_117),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_122),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_132),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_139),
.C(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_105),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_108),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_101),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_101),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_126),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_115),
.B(n_116),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_116),
.B(n_17),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_182),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_104),
.B1(n_112),
.B2(n_107),
.C(n_10),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_143),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_210),
.Y(n_220)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_133),
.B(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_131),
.Y(n_195)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_199),
.B(n_207),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_216),
.C(n_184),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_154),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_152),
.B1(n_125),
.B2(n_134),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_208),
.A2(n_160),
.B1(n_189),
.B2(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_177),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_160),
.A2(n_125),
.B1(n_118),
.B2(n_3),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_162),
.B1(n_188),
.B2(n_186),
.Y(n_234)
);

NOR4xp25_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_125),
.C(n_9),
.D(n_10),
.Y(n_213)
);

AOI321xp33_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_187),
.A3(n_182),
.B1(n_181),
.B2(n_183),
.C(n_11),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_186),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_16),
.C(n_14),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_163),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_238),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_163),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_234),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_233),
.B1(n_212),
.B2(n_208),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_235),
.C(n_237),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_171),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_193),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_232),
.B(n_197),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_189),
.A2(n_167),
.B1(n_165),
.B2(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_175),
.C(n_180),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_191),
.B(n_170),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_236),
.A2(n_191),
.B(n_197),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_175),
.C(n_167),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_168),
.B1(n_166),
.B2(n_158),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_166),
.C(n_179),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_196),
.C(n_216),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_215),
.C(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_238),
.B(n_225),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_193),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_255),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_194),
.B(n_207),
.C(n_215),
.D(n_196),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_220),
.B(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_203),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_157),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_233),
.B1(n_227),
.B2(n_218),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_267),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_230),
.C(n_217),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_274),
.C(n_243),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_258),
.B1(n_247),
.B2(n_225),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_247),
.B(n_246),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_221),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_229),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_283),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_279),
.B(n_276),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_252),
.B(n_249),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_266),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_241),
.C(n_255),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_287),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_253),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_261),
.B(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_249),
.C(n_237),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_271),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_288),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

OAI321xp33_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_215),
.A3(n_263),
.B1(n_256),
.B2(n_270),
.C(n_267),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_292),
.B(n_295),
.Y(n_305)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_231),
.B(n_235),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_299),
.A2(n_215),
.B1(n_206),
.B2(n_209),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_306),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_294),
.A2(n_271),
.B1(n_277),
.B2(n_204),
.Y(n_303)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_303),
.Y(n_311)
);

OAI221xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_262),
.B1(n_204),
.B2(n_206),
.C(n_14),
.Y(n_306)
);

AO221x1_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_14),
.B1(n_13),
.B2(n_3),
.C(n_4),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_2),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_309),
.A3(n_310),
.B1(n_312),
.B2(n_301),
.C1(n_6),
.C2(n_7),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_298),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_296),
.A3(n_13),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_5),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_305),
.A3(n_302),
.B1(n_13),
.B2(n_8),
.C1(n_7),
.C2(n_6),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_5),
.C(n_8),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_315),
.B(n_314),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule