module fake_jpeg_14933_n_348 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_0),
.Y(n_72)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_43),
.CON(n_59),
.SN(n_59)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_33),
.B1(n_20),
.B2(n_25),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_60),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_33),
.B1(n_20),
.B2(n_25),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_40),
.B1(n_45),
.B2(n_2),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_33),
.B1(n_24),
.B2(n_19),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_28),
.B1(n_26),
.B2(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_72),
.Y(n_97)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_46),
.B1(n_39),
.B2(n_42),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_79),
.B1(n_43),
.B2(n_59),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_46),
.B1(n_42),
.B2(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_81),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_100),
.B1(n_67),
.B2(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_43),
.B1(n_28),
.B2(n_26),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_93),
.B1(n_30),
.B2(n_29),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_43),
.B1(n_21),
.B2(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_103),
.Y(n_138)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_72),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_105),
.B1(n_125),
.B2(n_83),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_51),
.B1(n_62),
.B2(n_53),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_108),
.A2(n_128),
.B1(n_18),
.B2(n_29),
.Y(n_157)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_45),
.C(n_44),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_35),
.C(n_44),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_72),
.B1(n_73),
.B2(n_70),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_98),
.B1(n_77),
.B2(n_95),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_68),
.B1(n_53),
.B2(n_51),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_117),
.B1(n_90),
.B2(n_94),
.Y(n_145)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_50),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_50),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_35),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_31),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_57),
.B1(n_52),
.B2(n_50),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_90),
.B1(n_52),
.B2(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_147),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_150),
.B1(n_125),
.B2(n_102),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_137),
.C(n_156),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_0),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_136),
.B(n_154),
.Y(n_164)
);

AO22x2_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_48),
.B1(n_61),
.B2(n_91),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_148),
.B1(n_111),
.B2(n_123),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_101),
.C(n_113),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_112),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_157),
.B1(n_118),
.B2(n_123),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_107),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_83),
.B1(n_77),
.B2(n_48),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_153),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_37),
.B(n_66),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_37),
.C(n_27),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_158),
.A2(n_172),
.B1(n_173),
.B2(n_176),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_150),
.B1(n_134),
.B2(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_175),
.B1(n_176),
.B2(n_179),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_111),
.B1(n_126),
.B2(n_106),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_131),
.B(n_66),
.Y(n_203)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_127),
.B1(n_122),
.B2(n_109),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_122),
.B1(n_118),
.B2(n_61),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_112),
.B1(n_48),
.B2(n_14),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_136),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_138),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_212),
.B1(n_179),
.B2(n_160),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_194),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_137),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_200),
.C(n_207),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_184),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_156),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_181),
.B1(n_180),
.B2(n_174),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_196),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_154),
.B(n_147),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_203),
.B(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_139),
.C(n_146),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_136),
.A3(n_145),
.B1(n_149),
.B2(n_18),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_203),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_23),
.B(n_29),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_27),
.C(n_11),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_170),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_37),
.C(n_27),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_160),
.C(n_163),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_1),
.B(n_2),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_158),
.A2(n_165),
.B(n_175),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_172),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_215),
.C(n_222),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_171),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_235),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_250)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_211),
.B1(n_204),
.B2(n_193),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_187),
.B1(n_205),
.B2(n_193),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_234),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_30),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_169),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_227),
.C(n_230),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_183),
.C(n_37),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_233),
.B1(n_219),
.B2(n_230),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_195),
.B1(n_204),
.B2(n_192),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_209),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_37),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_30),
.Y(n_253)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_238),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_241),
.B(n_244),
.Y(n_268)
);

FAx1_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_202),
.CI(n_210),
.CON(n_243),
.SN(n_243)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_1),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_224),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_31),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_254),
.B(n_23),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_215),
.B1(n_221),
.B2(n_231),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_255),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_226),
.B(n_15),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_261),
.Y(n_280)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_214),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_266),
.C(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_222),
.C(n_223),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_30),
.C(n_22),
.Y(n_270)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_248),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_22),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_278),
.C(n_281),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_22),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_255),
.C(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_239),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_241),
.C(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_297),
.C(n_264),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_265),
.A2(n_243),
.B(n_257),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_294),
.C(n_268),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_250),
.B1(n_256),
.B2(n_247),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_276),
.B1(n_295),
.B2(n_297),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_296),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_263),
.A2(n_252),
.B(n_254),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_253),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_244),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_1),
.C(n_3),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_268),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_13),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_310),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_304),
.B1(n_311),
.B2(n_5),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_296),
.B1(n_284),
.B2(n_271),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_302),
.B(n_309),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_283),
.C(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_266),
.C(n_270),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_262),
.C(n_4),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_312),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_316),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_300),
.A2(n_3),
.B(n_4),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_12),
.B(n_11),
.Y(n_317)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_4),
.B(n_5),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_324),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_319),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_299),
.B(n_5),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_6),
.B(n_7),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_10),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_6),
.Y(n_332)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

XOR2x2_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_303),
.Y(n_326)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_326),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_334),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_306),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_332),
.B(n_316),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_320),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_335),
.B(n_336),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_323),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_324),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_337),
.A2(n_340),
.B(n_329),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_343),
.C(n_333),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_342),
.C(n_338),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_345),
.A2(n_316),
.B(n_8),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_10),
.B(n_7),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_8),
.C(n_340),
.Y(n_348)
);


endmodule