module fake_jpeg_5733_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_16),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_27),
.B(n_12),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_11),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_7),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_38),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_14),
.B1(n_19),
.B2(n_26),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_14),
.B1(n_19),
.B2(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_21),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_47),
.Y(n_50)
);

CKINVDCx10_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_35),
.C(n_25),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_44),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_61),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI21x1_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_48),
.B(n_53),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_52),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_52),
.B(n_51),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_66),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_63),
.C(n_9),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_71),
.Y(n_73)
);


endmodule