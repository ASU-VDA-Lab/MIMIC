module fake_ibex_1553_n_963 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_963);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_963;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_506;
wire n_444;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

BUFx3_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_33),
.B(n_99),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_98),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_19),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_62),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_30),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_71),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_113),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_21),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_10),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_55),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_5),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_102),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_121),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_86),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_104),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_72),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_110),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_34),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_10),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_14),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_27),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_60),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_3),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_48),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_74),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_82),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_131),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_95),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_66),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_22),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_150),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_111),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_127),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_73),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_106),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_20),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_114),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_159),
.Y(n_234)
);

INVxp33_ASAP7_75t_SL g235 ( 
.A(n_42),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_87),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_142),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_88),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_148),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_97),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_143),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_56),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_94),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_31),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_22),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_65),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_44),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_164),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_40),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_118),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_84),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_79),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_76),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_167),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_128),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_132),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_8),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_37),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_124),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_52),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_108),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_123),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_101),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g270 ( 
.A(n_46),
.B(n_93),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_11),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_11),
.B(n_37),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_4),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_14),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_6),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_105),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_141),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_43),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_135),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_119),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_45),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_17),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_157),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_39),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_153),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_34),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_1),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_64),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_221),
.A2(n_231),
.B1(n_223),
.B2(n_224),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g291 ( 
.A(n_177),
.B(n_0),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_177),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_177),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_180),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_2),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_181),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_202),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_186),
.A2(n_91),
.B(n_168),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_181),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_228),
.B(n_7),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_7),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_208),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_202),
.B(n_8),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_186),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_207),
.Y(n_309)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_208),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_207),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_174),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_185),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_195),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_175),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_184),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_178),
.B(n_12),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_212),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_170),
.B(n_12),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_211),
.Y(n_325)
);

AOI22x1_ASAP7_75t_SL g326 ( 
.A1(n_275),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_170),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_229),
.B(n_13),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_188),
.B(n_16),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_225),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_234),
.B(n_17),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_225),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_189),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_242),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_190),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_236),
.B(n_247),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_282),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_249),
.Y(n_339)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_212),
.A2(n_243),
.B(n_239),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_192),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_240),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_240),
.B(n_23),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_262),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_239),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_172),
.Y(n_347)
);

BUFx8_ASAP7_75t_L g348 ( 
.A(n_243),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_194),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_232),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_232),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_253),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_197),
.B(n_25),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_204),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_265),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_272),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_265),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_248),
.Y(n_359)
);

CKINVDCx6p67_ASAP7_75t_R g360 ( 
.A(n_172),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_271),
.B(n_26),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_230),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_198),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_200),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_230),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_201),
.B(n_28),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_205),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_206),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_209),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_290),
.A2(n_235),
.B1(n_264),
.B2(n_280),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_295),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_176),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_291),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_203),
.Y(n_377)
);

NOR3xp33_ASAP7_75t_L g378 ( 
.A(n_294),
.B(n_273),
.C(n_199),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_291),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_313),
.B(n_176),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

BUFx6f_ASAP7_75t_SL g383 ( 
.A(n_313),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_353),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_305),
.B(n_210),
.Y(n_388)
);

NAND2xp33_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_179),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_297),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_179),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_305),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_319),
.B(n_254),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_348),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_324),
.B(n_213),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_320),
.A2(n_235),
.B1(n_214),
.B2(n_286),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_319),
.B(n_215),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_324),
.B(n_216),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_320),
.A2(n_279),
.B1(n_219),
.B2(n_220),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_297),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_292),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_355),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_324),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_339),
.B(n_182),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_293),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_317),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_339),
.B(n_182),
.Y(n_422)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_298),
.B(n_270),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_363),
.B(n_183),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_306),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_317),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_321),
.B(n_187),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_296),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_333),
.B(n_256),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_306),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

NOR2x1p5_ASAP7_75t_L g433 ( 
.A(n_360),
.B(n_256),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_L g434 ( 
.A(n_304),
.B(n_258),
.C(n_257),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_311),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_329),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_333),
.B(n_226),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_335),
.B(n_257),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_359),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_322),
.B(n_258),
.Y(n_441)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_352),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_336),
.B(n_241),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_336),
.B(n_260),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_322),
.B(n_260),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_310),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_347),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_310),
.Y(n_453)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_328),
.Y(n_455)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_366),
.B(n_328),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_310),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_341),
.B(n_263),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_310),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_310),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_SL g461 ( 
.A1(n_341),
.A2(n_250),
.B(n_244),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_301),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_311),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_301),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_369),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_349),
.B(n_251),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_337),
.B(n_288),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_301),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_314),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_314),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_314),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_369),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_369),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_330),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_362),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_331),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_303),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_303),
.Y(n_479)
);

NAND2xp33_ASAP7_75t_L g480 ( 
.A(n_364),
.B(n_266),
.Y(n_480)
);

AOI22x1_ASAP7_75t_L g481 ( 
.A1(n_364),
.A2(n_255),
.B1(n_259),
.B2(n_284),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_331),
.B(n_287),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_332),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_468),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_332),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_381),
.B(n_393),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_408),
.B(n_315),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_424),
.B(n_342),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_400),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_415),
.B(n_316),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_428),
.B(n_362),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_377),
.B(n_344),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_398),
.B(n_361),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_396),
.B(n_422),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_382),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_437),
.A2(n_368),
.B(n_367),
.C(n_354),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_439),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_455),
.B(n_440),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_441),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_390),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_462),
.Y(n_504)
);

O2A1O1Ixp5_ASAP7_75t_L g505 ( 
.A1(n_388),
.A2(n_367),
.B(n_368),
.C(n_346),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_450),
.B(n_346),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_371),
.B(n_173),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_434),
.B(n_318),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_405),
.B(n_325),
.Y(n_509)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_456),
.B(n_375),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_456),
.B(n_345),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_470),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_386),
.Y(n_513)
);

INVx8_ASAP7_75t_L g514 ( 
.A(n_383),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_418),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_389),
.A2(n_357),
.B1(n_338),
.B2(n_365),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_379),
.B(n_299),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_389),
.A2(n_365),
.B1(n_326),
.B2(n_350),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_299),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_380),
.A2(n_308),
.B1(n_350),
.B2(n_309),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_472),
.B(n_302),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_472),
.B(n_191),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_410),
.B(n_238),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_414),
.B(n_193),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_436),
.B(n_196),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_427),
.A2(n_326),
.B1(n_358),
.B2(n_323),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_383),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_402),
.B(n_217),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_430),
.B(n_218),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_376),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_307),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_376),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_401),
.B(n_406),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_372),
.A2(n_323),
.B1(n_312),
.B2(n_358),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_222),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_227),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_478),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_480),
.B(n_233),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_402),
.B(n_237),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_465),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_469),
.Y(n_542)
);

NOR3xp33_ASAP7_75t_L g543 ( 
.A(n_378),
.B(n_171),
.C(n_269),
.Y(n_543)
);

NOR3xp33_ASAP7_75t_L g544 ( 
.A(n_461),
.B(n_277),
.C(n_281),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_401),
.B(n_245),
.Y(n_545)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_416),
.Y(n_546)
);

O2A1O1Ixp5_ASAP7_75t_L g547 ( 
.A1(n_418),
.A2(n_420),
.B(n_419),
.C(n_373),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_442),
.A2(n_276),
.B1(n_246),
.B2(n_285),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_370),
.B(n_307),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_442),
.A2(n_283),
.B1(n_278),
.B2(n_268),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_395),
.B(n_252),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_395),
.B(n_300),
.Y(n_552)
);

O2A1O1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_423),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_419),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_412),
.B(n_32),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_447),
.B(n_35),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_454),
.B(n_38),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_447),
.B(n_36),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_476),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_433),
.B(n_36),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_454),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_467),
.B(n_54),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_496),
.A2(n_423),
.B(n_417),
.C(n_409),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_SL g565 ( 
.A(n_484),
.B(n_394),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_488),
.B(n_394),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_542),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_531),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_492),
.B(n_394),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_493),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_492),
.B(n_407),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_407),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_510),
.A2(n_423),
.B1(n_467),
.B2(n_452),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_510),
.B(n_475),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_552),
.A2(n_420),
.B(n_431),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_547),
.A2(n_435),
.B(n_425),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_515),
.A2(n_464),
.B1(n_479),
.B2(n_481),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_503),
.B(n_451),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_515),
.A2(n_463),
.B(n_474),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_501),
.B(n_476),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_503),
.B(n_451),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_547),
.A2(n_474),
.B(n_473),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_514),
.B(n_463),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_453),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_497),
.A2(n_466),
.B(n_374),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_495),
.B(n_453),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_509),
.B(n_457),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_486),
.A2(n_374),
.B(n_413),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_508),
.B(n_544),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_554),
.A2(n_460),
.B1(n_459),
.B2(n_457),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_546),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_486),
.A2(n_397),
.B(n_411),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_494),
.A2(n_397),
.B(n_411),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_514),
.B(n_459),
.Y(n_596)
);

OR2x6_ASAP7_75t_SL g597 ( 
.A(n_560),
.B(n_460),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_554),
.A2(n_385),
.B1(n_391),
.B2(n_392),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_522),
.B(n_525),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_508),
.B(n_392),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_502),
.B(n_57),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_500),
.B(n_399),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_506),
.B(n_403),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_499),
.A2(n_403),
.B1(n_404),
.B2(n_413),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_L g605 ( 
.A(n_549),
.B(n_404),
.C(n_448),
.Y(n_605)
);

CKINVDCx14_ASAP7_75t_R g606 ( 
.A(n_518),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_528),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_532),
.B(n_58),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_546),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_516),
.B(n_528),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_529),
.B(n_59),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g612 ( 
.A1(n_563),
.A2(n_446),
.B(n_445),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_523),
.B(n_61),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_533),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_520),
.A2(n_445),
.B1(n_444),
.B2(n_426),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_546),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_521),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_561),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_545),
.B(n_67),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_538),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_540),
.B(n_70),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_505),
.A2(n_438),
.B(n_432),
.C(n_429),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_520),
.A2(n_432),
.B1(n_429),
.B2(n_443),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_507),
.B(n_75),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_535),
.A2(n_443),
.B1(n_421),
.B2(n_387),
.Y(n_626)
);

AO21x1_ASAP7_75t_L g627 ( 
.A1(n_562),
.A2(n_80),
.B(n_81),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_545),
.B(n_83),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_505),
.A2(n_443),
.B(n_421),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_483),
.A2(n_485),
.B(n_490),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_524),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_535),
.A2(n_384),
.B1(n_387),
.B2(n_92),
.Y(n_632)
);

O2A1O1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_556),
.A2(n_169),
.B(n_100),
.C(n_103),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_517),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_548),
.B(n_109),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_541),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_558),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_559),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_555),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_559),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_551),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_526),
.A2(n_133),
.B1(n_134),
.B2(n_139),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_550),
.B(n_140),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_568),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_617),
.B(n_504),
.Y(n_645)
);

NAND2x1p5_ASAP7_75t_L g646 ( 
.A(n_617),
.B(n_489),
.Y(n_646)
);

AO31x2_ASAP7_75t_L g647 ( 
.A1(n_627),
.A2(n_557),
.A3(n_512),
.B(n_527),
.Y(n_647)
);

INVxp67_ASAP7_75t_SL g648 ( 
.A(n_613),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_577),
.B(n_553),
.Y(n_649)
);

AO31x2_ASAP7_75t_L g650 ( 
.A1(n_604),
.A2(n_487),
.A3(n_498),
.B(n_513),
.Y(n_650)
);

OA21x2_ASAP7_75t_L g651 ( 
.A1(n_578),
.A2(n_537),
.B(n_539),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_593),
.Y(n_652)
);

BUFx8_ASAP7_75t_L g653 ( 
.A(n_593),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_636),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_634),
.B(n_591),
.Y(n_655)
);

OA21x2_ASAP7_75t_L g656 ( 
.A1(n_578),
.A2(n_536),
.B(n_530),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_618),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_630),
.A2(n_145),
.B(n_146),
.C(n_147),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_571),
.B(n_155),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_593),
.B(n_156),
.Y(n_661)
);

AOI221xp5_ASAP7_75t_L g662 ( 
.A1(n_582),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.C(n_166),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_597),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_609),
.Y(n_664)
);

OAI22x1_ASAP7_75t_L g665 ( 
.A1(n_574),
.A2(n_625),
.B1(n_642),
.B2(n_610),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_599),
.A2(n_594),
.B(n_590),
.Y(n_666)
);

AO31x2_ASAP7_75t_L g667 ( 
.A1(n_598),
.A2(n_632),
.A3(n_579),
.B(n_592),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_573),
.B(n_608),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_641),
.B(n_564),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_607),
.B(n_631),
.Y(n_670)
);

O2A1O1Ixp5_ASAP7_75t_L g671 ( 
.A1(n_622),
.A2(n_620),
.B(n_628),
.C(n_611),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_609),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_605),
.A2(n_570),
.B1(n_606),
.B2(n_566),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_SL g674 ( 
.A(n_609),
.B(n_585),
.Y(n_674)
);

AO31x2_ASAP7_75t_L g675 ( 
.A1(n_598),
.A2(n_623),
.A3(n_616),
.B(n_600),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_619),
.B(n_575),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_581),
.A2(n_586),
.B(n_589),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_565),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_637),
.B(n_633),
.C(n_601),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_569),
.B(n_615),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_621),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_580),
.B(n_583),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_587),
.A2(n_603),
.B(n_595),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_602),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_639),
.A2(n_614),
.B1(n_643),
.B2(n_635),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_588),
.B(n_638),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_588),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_640),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_585),
.A2(n_627),
.A3(n_604),
.B(n_626),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_596),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_630),
.A2(n_486),
.B(n_492),
.C(n_572),
.Y(n_691)
);

AO31x2_ASAP7_75t_L g692 ( 
.A1(n_627),
.A2(n_604),
.A3(n_626),
.B(n_624),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_568),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_576),
.A2(n_547),
.B(n_630),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_568),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_629),
.A2(n_612),
.B(n_584),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_576),
.A2(n_552),
.B(n_515),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_630),
.A2(n_486),
.B(n_492),
.C(n_572),
.Y(n_698)
);

NAND3x1_ASAP7_75t_L g699 ( 
.A(n_582),
.B(n_518),
.C(n_334),
.Y(n_699)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_582),
.A2(n_428),
.B(n_484),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_636),
.Y(n_701)
);

OAI21xp33_ASAP7_75t_L g702 ( 
.A1(n_582),
.A2(n_428),
.B(n_484),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_568),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_568),
.B(n_484),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_636),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_577),
.B(n_514),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_572),
.A2(n_510),
.B1(n_634),
.B2(n_456),
.Y(n_707)
);

AND2x6_ASAP7_75t_L g708 ( 
.A(n_593),
.B(n_609),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_577),
.Y(n_709)
);

OAI21xp33_ASAP7_75t_L g710 ( 
.A1(n_582),
.A2(n_428),
.B(n_484),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_636),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_571),
.B(n_484),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_636),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_568),
.B(n_484),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_568),
.Y(n_715)
);

AO31x2_ASAP7_75t_L g716 ( 
.A1(n_627),
.A2(n_604),
.A3(n_626),
.B(n_624),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_568),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_582),
.B(n_493),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_SL g719 ( 
.A(n_617),
.B(n_362),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_613),
.B(n_484),
.Y(n_720)
);

NAND3xp33_ASAP7_75t_L g721 ( 
.A(n_582),
.B(n_543),
.C(n_544),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_627),
.A2(n_604),
.A3(n_626),
.B(n_624),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_617),
.B(n_577),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_629),
.A2(n_612),
.B(n_584),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_613),
.B(n_484),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_613),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_613),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_629),
.A2(n_612),
.B(n_584),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_652),
.B(n_663),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_658),
.B(n_652),
.Y(n_730)
);

OA21x2_ASAP7_75t_L g731 ( 
.A1(n_696),
.A2(n_728),
.B(n_724),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_694),
.A2(n_666),
.B(n_683),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_705),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_644),
.Y(n_734)
);

AOI21xp33_ASAP7_75t_SL g735 ( 
.A1(n_718),
.A2(n_700),
.B(n_710),
.Y(n_735)
);

NOR2x1_ASAP7_75t_R g736 ( 
.A(n_652),
.B(n_723),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_723),
.B(n_648),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_653),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_654),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_701),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_711),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_713),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_668),
.A2(n_655),
.B(n_721),
.C(n_685),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_677),
.A2(n_671),
.B(n_679),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_726),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_702),
.A2(n_727),
.B1(n_719),
.B2(n_720),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_651),
.A2(n_656),
.B(n_686),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_657),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_725),
.B(n_712),
.Y(n_750)
);

AOI21xp33_ASAP7_75t_SL g751 ( 
.A1(n_706),
.A2(n_704),
.B(n_714),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_665),
.A2(n_669),
.B1(n_673),
.B2(n_649),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_659),
.A2(n_681),
.B(n_682),
.Y(n_753)
);

OAI21x1_ASAP7_75t_L g754 ( 
.A1(n_664),
.A2(n_660),
.B(n_646),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_684),
.Y(n_755)
);

OA21x2_ASAP7_75t_L g756 ( 
.A1(n_662),
.A2(n_722),
.B(n_716),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_653),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_688),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_672),
.B(n_674),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_693),
.B(n_703),
.Y(n_760)
);

OAI21x1_ASAP7_75t_L g761 ( 
.A1(n_650),
.A2(n_675),
.B(n_689),
.Y(n_761)
);

AO31x2_ASAP7_75t_L g762 ( 
.A1(n_647),
.A2(n_675),
.A3(n_722),
.B(n_716),
.Y(n_762)
);

OA21x2_ASAP7_75t_L g763 ( 
.A1(n_692),
.A2(n_722),
.B(n_716),
.Y(n_763)
);

INVx3_ASAP7_75t_SL g764 ( 
.A(n_706),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_647),
.A2(n_692),
.B(n_689),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_667),
.B(n_676),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_667),
.B(n_699),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_717),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_690),
.A2(n_647),
.B(n_678),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_661),
.A2(n_645),
.B(n_670),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_709),
.Y(n_771)
);

NAND2x1p5_ASAP7_75t_L g772 ( 
.A(n_645),
.B(n_661),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_650),
.A2(n_675),
.B(n_689),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_687),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_692),
.B(n_708),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_715),
.B(n_695),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_708),
.A2(n_698),
.B(n_691),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_691),
.A2(n_698),
.B(n_697),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_691),
.A2(n_698),
.B(n_694),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_658),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_691),
.A2(n_698),
.B(n_694),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_655),
.B(n_658),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_691),
.A2(n_698),
.B(n_697),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_691),
.A2(n_698),
.B(n_668),
.C(n_707),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_718),
.A2(n_510),
.B1(n_702),
.B2(n_700),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_655),
.B(n_658),
.Y(n_786)
);

INVx6_ASAP7_75t_L g787 ( 
.A(n_653),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_705),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_691),
.A2(n_698),
.B(n_697),
.Y(n_789)
);

INVx4_ASAP7_75t_SL g790 ( 
.A(n_708),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_648),
.B(n_726),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_691),
.A2(n_698),
.B(n_697),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_648),
.B(n_726),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_658),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_655),
.B(n_658),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_691),
.A2(n_698),
.B(n_668),
.C(n_707),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_733),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_791),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_793),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_731),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_748),
.B(n_750),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_788),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_782),
.B(n_786),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_737),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_795),
.B(n_780),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_795),
.B(n_794),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_752),
.A2(n_785),
.B1(n_767),
.B2(n_755),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_737),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_790),
.B(n_777),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_739),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_787),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_740),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_772),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_741),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_767),
.B(n_766),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_742),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_766),
.B(n_743),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_735),
.B(n_755),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_730),
.B(n_754),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_749),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_770),
.B(n_796),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_759),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_770),
.B(n_784),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_745),
.B(n_763),
.Y(n_824)
);

AO21x2_ASAP7_75t_L g825 ( 
.A1(n_744),
.A2(n_792),
.B(n_789),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_775),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_759),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_776),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_SL g829 ( 
.A1(n_787),
.A2(n_768),
.B1(n_738),
.B2(n_734),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_778),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_778),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_763),
.B(n_746),
.Y(n_832)
);

OA21x2_ASAP7_75t_L g833 ( 
.A1(n_744),
.A2(n_732),
.B(n_781),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_736),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_734),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_765),
.B(n_762),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_760),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_758),
.B(n_771),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_729),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_787),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_824),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_824),
.B(n_765),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_800),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_803),
.B(n_779),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_803),
.B(n_761),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_819),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_836),
.B(n_773),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_836),
.B(n_762),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_826),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_805),
.B(n_762),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_801),
.B(n_738),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_815),
.B(n_798),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_819),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_809),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_817),
.B(n_779),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_818),
.B(n_751),
.C(n_783),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_822),
.Y(n_857)
);

AND2x4_ASAP7_75t_SL g858 ( 
.A(n_804),
.B(n_790),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_817),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_806),
.B(n_756),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_835),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_797),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_806),
.B(n_825),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_822),
.Y(n_864)
);

AOI221xp5_ASAP7_75t_L g865 ( 
.A1(n_821),
.A2(n_753),
.B1(n_769),
.B2(n_764),
.C(n_757),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_823),
.B(n_747),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_863),
.B(n_848),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_852),
.B(n_810),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_862),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_854),
.B(n_809),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_863),
.B(n_832),
.Y(n_871)
);

INVxp67_ASAP7_75t_SL g872 ( 
.A(n_849),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_852),
.B(n_831),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_850),
.B(n_812),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_859),
.B(n_841),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_843),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_846),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_848),
.B(n_845),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_850),
.B(n_812),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_845),
.B(n_832),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_861),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_860),
.B(n_833),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_844),
.B(n_830),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_860),
.B(n_833),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_881),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_876),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_867),
.B(n_861),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_869),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_878),
.B(n_847),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_869),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_878),
.B(n_847),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_867),
.B(n_868),
.Y(n_892)
);

INVxp33_ASAP7_75t_L g893 ( 
.A(n_874),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_871),
.B(n_842),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_871),
.B(n_842),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_877),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_879),
.B(n_873),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_880),
.B(n_866),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_873),
.B(n_844),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_880),
.B(n_855),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_875),
.B(n_855),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_882),
.B(n_866),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_894),
.B(n_895),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_896),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_885),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_889),
.B(n_882),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_896),
.A2(n_872),
.B(n_853),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_888),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_887),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_892),
.B(n_884),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_902),
.B(n_870),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_888),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_889),
.B(n_884),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_890),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_886),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_906),
.B(n_913),
.Y(n_916)
);

OAI31xp33_ASAP7_75t_L g917 ( 
.A1(n_907),
.A2(n_904),
.A3(n_834),
.B(n_893),
.Y(n_917)
);

OAI21xp33_ASAP7_75t_L g918 ( 
.A1(n_904),
.A2(n_891),
.B(n_902),
.Y(n_918)
);

OAI322xp33_ASAP7_75t_L g919 ( 
.A1(n_910),
.A2(n_900),
.A3(n_897),
.B1(n_901),
.B2(n_899),
.C1(n_875),
.C2(n_883),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_908),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_911),
.B(n_877),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_912),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_914),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_906),
.B(n_891),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_L g925 ( 
.A(n_905),
.B(n_829),
.C(n_856),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_909),
.Y(n_926)
);

OAI32xp33_ASAP7_75t_L g927 ( 
.A1(n_909),
.A2(n_900),
.A3(n_901),
.B1(n_857),
.B2(n_898),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_917),
.A2(n_926),
.B(n_918),
.Y(n_928)
);

AOI221xp5_ASAP7_75t_L g929 ( 
.A1(n_919),
.A2(n_903),
.B1(n_913),
.B2(n_911),
.C(n_856),
.Y(n_929)
);

AOI221xp5_ASAP7_75t_SL g930 ( 
.A1(n_927),
.A2(n_840),
.B1(n_910),
.B2(n_851),
.C(n_898),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_925),
.A2(n_911),
.B1(n_894),
.B2(n_895),
.Y(n_931)
);

AOI21xp33_ASAP7_75t_SL g932 ( 
.A1(n_921),
.A2(n_834),
.B(n_811),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_916),
.B(n_915),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_929),
.B(n_931),
.Y(n_934)
);

AOI221xp5_ASAP7_75t_L g935 ( 
.A1(n_928),
.A2(n_923),
.B1(n_922),
.B2(n_920),
.C(n_916),
.Y(n_935)
);

AOI221xp5_ASAP7_75t_L g936 ( 
.A1(n_930),
.A2(n_924),
.B1(n_921),
.B2(n_828),
.C(n_865),
.Y(n_936)
);

NOR2x1_ASAP7_75t_L g937 ( 
.A(n_934),
.B(n_857),
.Y(n_937)
);

NAND4xp75_ASAP7_75t_L g938 ( 
.A(n_935),
.B(n_811),
.C(n_823),
.D(n_865),
.Y(n_938)
);

AND5x1_ASAP7_75t_L g939 ( 
.A(n_938),
.B(n_936),
.C(n_932),
.D(n_769),
.E(n_753),
.Y(n_939)
);

NOR2x1_ASAP7_75t_L g940 ( 
.A(n_937),
.B(n_857),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_940),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_939),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_941),
.B(n_933),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_942),
.B(n_924),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_944),
.A2(n_839),
.B1(n_921),
.B2(n_837),
.Y(n_945)
);

OA22x2_ASAP7_75t_L g946 ( 
.A1(n_943),
.A2(n_838),
.B1(n_799),
.B2(n_858),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_943),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_947),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_945),
.B(n_810),
.Y(n_949)
);

NOR2xp67_ASAP7_75t_L g950 ( 
.A(n_946),
.B(n_857),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_947),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_948),
.B(n_915),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_951),
.A2(n_774),
.B(n_816),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_949),
.A2(n_816),
.B(n_814),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_950),
.B(n_814),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_951),
.B(n_820),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_948),
.A2(n_807),
.B1(n_864),
.B2(n_858),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_952),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_956),
.A2(n_820),
.B(n_802),
.Y(n_959)
);

OA21x2_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_953),
.B(n_955),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_959),
.A2(n_957),
.B(n_954),
.Y(n_961)
);

OA22x2_ASAP7_75t_L g962 ( 
.A1(n_961),
.A2(n_858),
.B1(n_808),
.B2(n_813),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_962),
.A2(n_960),
.B1(n_864),
.B2(n_827),
.Y(n_963)
);


endmodule