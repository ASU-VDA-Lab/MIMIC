module real_jpeg_6778_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_1),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_1),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_1),
.A2(n_187),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_1),
.A2(n_187),
.B1(n_404),
.B2(n_406),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_1),
.A2(n_187),
.B1(n_459),
.B2(n_464),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_2),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_40),
.B1(n_86),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_3),
.A2(n_40),
.B1(n_46),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_3),
.A2(n_40),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_4),
.B(n_268),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_4),
.A2(n_267),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_4),
.B(n_192),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_4),
.B(n_37),
.C(n_377),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_L g380 ( 
.A1(n_4),
.A2(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_4),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_4),
.B(n_138),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_4),
.A2(n_26),
.B1(n_425),
.B2(n_428),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_5),
.A2(n_258),
.B1(n_284),
.B2(n_286),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_5),
.A2(n_286),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_5),
.A2(n_286),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_5),
.A2(n_286),
.B1(n_409),
.B2(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_6),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_6),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_6),
.A2(n_291),
.B1(n_322),
.B2(n_326),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_6),
.A2(n_291),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_6),
.A2(n_160),
.B1(n_291),
.B2(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_7),
.Y(n_514)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_9),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_9),
.Y(n_307)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_9),
.Y(n_342)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_9),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_10),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_77),
.B1(n_105),
.B2(n_108),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_77),
.B1(n_160),
.B2(n_165),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_10),
.A2(n_77),
.B1(n_118),
.B2(n_197),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_11),
.Y(n_262)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_13),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_13),
.Y(n_190)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_13),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_14),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_15),
.A2(n_44),
.B1(n_140),
.B2(n_144),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_15),
.A2(n_44),
.B1(n_237),
.B2(n_239),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_15),
.A2(n_44),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_17),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_17),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_17),
.A2(n_117),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_17),
.A2(n_117),
.B1(n_189),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_17),
.A2(n_117),
.B1(n_161),
.B2(n_273),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_508),
.B(n_511),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_496),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_216),
.A3(n_241),
.B(n_493),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_198),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_22),
.B(n_198),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_111),
.C(n_154),
.Y(n_22)
);

FAx1_ASAP7_75t_L g367 ( 
.A(n_23),
.B(n_111),
.CI(n_154),
.CON(n_367),
.SN(n_367)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_80),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_24),
.A2(n_25),
.B(n_82),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_25),
.A2(n_81),
.B1(n_82),
.B2(n_110),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_25),
.A2(n_41),
.B1(n_81),
.B2(n_359),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_34),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_26),
.B(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_26),
.A2(n_271),
.B1(n_276),
.B2(n_277),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_26),
.A2(n_277),
.B(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_26),
.A2(n_168),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_26),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_26),
.A2(n_414),
.B1(n_425),
.B2(n_428),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_26),
.A2(n_34),
.B(n_306),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_31),
.Y(n_419)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_34),
.Y(n_169)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_41),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_54),
.B(n_70),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_43),
.A2(n_55),
.B1(n_71),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_48),
.Y(n_390)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_48),
.Y(n_447)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_49),
.Y(n_463)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_50),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_50),
.Y(n_383)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_50),
.Y(n_386)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_53),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_120)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_53),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_54),
.B(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_54),
.A2(n_72),
.B(n_148),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_54),
.A2(n_72),
.B1(n_152),
.B2(n_176),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_54),
.A2(n_70),
.B(n_148),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_54),
.A2(n_477),
.B(n_478),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_55),
.A2(n_71),
.B1(n_380),
.B2(n_387),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_55),
.A2(n_71),
.B1(n_387),
.B2(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_55),
.A2(n_71),
.B1(n_398),
.B2(n_458),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_64),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_56)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_57),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_63),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_67),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_67),
.Y(n_405)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_67),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_69),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_72),
.B(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_76),
.Y(n_399)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_101),
.B(n_103),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_83),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_83),
.A2(n_192),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_83),
.A2(n_192),
.B1(n_283),
.B2(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_84),
.A2(n_184),
.B(n_191),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_84),
.A2(n_109),
.B1(n_184),
.B2(n_288),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_84),
.A2(n_109),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_84),
.A2(n_503),
.B(n_504),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_94),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_85)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_93),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_96),
.Y(n_257)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_97),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_97),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_101),
.B(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_103),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_104),
.Y(n_213)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_106),
.Y(n_290)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_108),
.Y(n_293)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_109),
.A2(n_209),
.B(n_212),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_146),
.B(n_153),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_112),
.B(n_146),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_119),
.B1(n_138),
.B2(n_139),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_114),
.A2(n_120),
.B(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_115),
.Y(n_249)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_119),
.B(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_119),
.A2(n_139),
.B(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_119),
.A2(n_227),
.B(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_119),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_119),
.A2(n_138),
.B1(n_347),
.B2(n_456),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_119),
.A2(n_138),
.B(n_501),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_128),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_120),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_120),
.A2(n_301),
.B1(n_321),
.B2(n_329),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_120),
.A2(n_301),
.B1(n_321),
.B2(n_346),
.Y(n_345)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g448 ( 
.A(n_123),
.Y(n_448)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_125),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_131),
.B1(n_134),
.B2(n_137),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_136),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_138),
.B(n_196),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g456 ( 
.A1(n_140),
.A2(n_381),
.B(n_449),
.Y(n_456)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_142),
.Y(n_348)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_147),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_153),
.B(n_199),
.CI(n_215),
.CON(n_198),
.SN(n_198)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_182),
.C(n_193),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_155),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_173),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_156),
.A2(n_173),
.B1(n_174),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_156),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_168),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_158),
.A2(n_272),
.B(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_159),
.Y(n_308)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_162),
.Y(n_427)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_163),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_164),
.Y(n_280)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_166),
.B(n_434),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_172),
.Y(n_276)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_182),
.A2(n_183),
.B1(n_193),
.B2(n_194),
.Y(n_361)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_198),
.B(n_218),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_208),
.B2(n_214),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_207),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_202),
.B(n_224),
.C(n_234),
.Y(n_505)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_205),
.A2(n_228),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_208),
.B(n_219),
.C(n_222),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_210),
.Y(n_258)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_211),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_217),
.A2(n_494),
.B(n_495),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_228),
.Y(n_501)
);

INVx8_ASAP7_75t_L g444 ( 
.A(n_229),
.Y(n_444)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_233),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_236),
.Y(n_503)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_368),
.B(n_487),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_353),
.C(n_365),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_331),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_244),
.A2(n_489),
.B(n_490),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_310),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_245),
.B(n_310),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_294),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_246),
.B(n_295),
.C(n_297),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_253),
.C(n_282),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx6_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_270),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_254),
.B(n_270),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_258),
.A3(n_259),
.B1(n_263),
.B2(n_266),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g350 ( 
.A(n_257),
.Y(n_350)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_275),
.Y(n_415)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_304),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_299),
.B(n_303),
.C(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_309),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.C(n_330),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_330),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.C(n_320),
.Y(n_313)
);

FAx1_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_315),
.CI(n_320),
.CON(n_333),
.SN(n_333)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_326),
.B(n_381),
.Y(n_449)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_351),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_332),
.B(n_351),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.C(n_335),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_333),
.B(n_485),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_333),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_334),
.B(n_335),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_343),
.C(n_345),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_336),
.A2(n_337),
.B1(n_343),
.B2(n_344),
.Y(n_472)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_381),
.Y(n_434)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_345),
.B(n_472),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

A2O1A1O1Ixp25_ASAP7_75t_L g487 ( 
.A1(n_353),
.A2(n_365),
.B(n_488),
.C(n_491),
.D(n_492),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_364),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_354),
.B(n_364),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_358),
.C(n_363),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_360),
.B1(n_362),
.B2(n_363),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_358),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_360),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_366),
.B(n_367),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_367),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_482),
.B(n_486),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_467),
.B(n_481),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_438),
.B(n_466),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_410),
.B(n_437),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_393),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_373),
.B(n_393),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_379),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_379),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_402),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_397),
.B2(n_401),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_401),
.C(n_402),
.Y(n_439)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_397),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_451),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_403),
.Y(n_417)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_421),
.B(n_436),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_420),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_420),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_422),
.A2(n_431),
.B(n_435),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_423),
.B(n_424),
.Y(n_435)
);

INVx4_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_440),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_454),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_455),
.C(n_457),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_453),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_453),
.Y(n_475)
);

OAI32xp33_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_445),
.A3(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx6_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_458),
.Y(n_477)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_468),
.B(n_469),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_473),
.B2(n_474),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_476),
.C(n_479),
.Y(n_483)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_475),
.A2(n_476),
.B1(n_479),
.B2(n_480),
.Y(n_474)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_475),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_476),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_483),
.B(n_484),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_506),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_499),
.Y(n_507)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_499),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_502),
.CI(n_505),
.CON(n_499),
.SN(n_499)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

BUFx4f_ASAP7_75t_SL g508 ( 
.A(n_509),
.Y(n_508)
);

INVx13_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_510),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.Y(n_511)
);

BUFx12f_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);


endmodule