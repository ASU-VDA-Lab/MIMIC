module fake_netlist_5_2056_n_1749 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1749);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1749;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx5_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_28),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_84),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_74),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_78),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_43),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_96),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_105),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_28),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_69),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_23),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_63),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_26),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_46),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_35),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_68),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_73),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_60),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_116),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_0),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_91),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_30),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_85),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_75),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_21),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_121),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_104),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_30),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_36),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_77),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_56),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_21),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_50),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_26),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_0),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_31),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_61),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_19),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_54),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_22),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_122),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_81),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_22),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_31),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_79),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_29),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_2),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_47),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_58),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_72),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_55),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_7),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_51),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_134),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_27),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_71),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_115),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_14),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_34),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_111),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_34),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_106),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_50),
.Y(n_243)
);

INVx4_ASAP7_75t_R g244 ( 
.A(n_46),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_17),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_45),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_94),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_7),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_109),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_67),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_59),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_76),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_124),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_103),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_40),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_19),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_38),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_53),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_47),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_70),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_80),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_25),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_20),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_90),
.Y(n_271)
);

CKINVDCx12_ASAP7_75t_R g272 ( 
.A(n_36),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_12),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_16),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_33),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_5),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_137),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_87),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_38),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_133),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_17),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_23),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_5),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_42),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_83),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_12),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_52),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_151),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_95),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_129),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_27),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_1),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_118),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_98),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_33),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_107),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_49),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_120),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_82),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_18),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_1),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_48),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_298),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_190),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_191),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_193),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_153),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_153),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_153),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_154),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_235),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_290),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_194),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_153),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_153),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_200),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_199),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_241),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_207),
.Y(n_322)
);

BUFx6f_ASAP7_75t_SL g323 ( 
.A(n_163),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_177),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_211),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_213),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_214),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_187),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_215),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_153),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_236),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_153),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_153),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_2),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_242),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_222),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_236),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_222),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_216),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_178),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_222),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_222),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_219),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_227),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_203),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_305),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_233),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_253),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_254),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_223),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_248),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_223),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_248),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_277),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_155),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_278),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_285),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_288),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_162),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_294),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_173),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_164),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_186),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_203),
.B(n_3),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_255),
.B(n_3),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_192),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_204),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_218),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_289),
.B(n_4),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_188),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_232),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_196),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_157),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_237),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_202),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_238),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_205),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_206),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_178),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_365),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_336),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_157),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_165),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_178),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_339),
.B(n_178),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_343),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_312),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_331),
.A2(n_184),
.B(n_182),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

OR2x6_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_178),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_198),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_335),
.B(n_201),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_337),
.B(n_158),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_362),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_368),
.B(n_158),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_364),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_367),
.B(n_208),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_366),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_372),
.B(n_163),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_306),
.A2(n_250),
.B1(n_303),
.B2(n_302),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_338),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_371),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_329),
.A2(n_243),
.B1(n_221),
.B2(n_279),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_354),
.B(n_356),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_313),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_356),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_315),
.B(n_210),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_307),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_409),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_308),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_309),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_409),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_426),
.B(n_316),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_426),
.A2(n_320),
.B1(n_350),
.B2(n_347),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_383),
.Y(n_463)
);

BUFx4f_ASAP7_75t_L g464 ( 
.A(n_417),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_382),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_319),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_408),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_413),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_408),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_382),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_384),
.B(n_322),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_389),
.B(n_415),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_411),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_411),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

BUFx4f_ASAP7_75t_L g481 ( 
.A(n_417),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_384),
.B(n_325),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_L g484 ( 
.A(n_418),
.B(n_326),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_437),
.A2(n_329),
.B1(n_197),
.B2(n_217),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_415),
.B(n_226),
.C(n_224),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_417),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_423),
.A2(n_265),
.B1(n_282),
.B2(n_281),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_SL g491 ( 
.A(n_428),
.B(n_376),
.Y(n_491)
);

BUFx8_ASAP7_75t_SL g492 ( 
.A(n_441),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_387),
.B(n_327),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_437),
.A2(n_225),
.B1(n_189),
.B2(n_262),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_390),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_450),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_390),
.Y(n_499)
);

AOI21x1_ASAP7_75t_L g500 ( 
.A1(n_391),
.A2(n_239),
.B(n_228),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_391),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_387),
.B(n_330),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_385),
.Y(n_505)
);

INVx4_ASAP7_75t_SL g506 ( 
.A(n_417),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_423),
.A2(n_450),
.B1(n_412),
.B2(n_421),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_389),
.B(n_378),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_385),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_415),
.B(n_249),
.C(n_245),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_391),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_385),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_394),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_392),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_392),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_382),
.B(n_342),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_389),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_415),
.B(n_380),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_394),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_421),
.B(n_346),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_406),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_393),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_396),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_L g529 ( 
.A(n_430),
.B(n_349),
.C(n_353),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_440),
.B(n_423),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_394),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_394),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_412),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_442),
.B(n_257),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_414),
.B(n_267),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_442),
.B(n_351),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_406),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_394),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_431),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_396),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_442),
.B(n_352),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_398),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_394),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_406),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_398),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_398),
.Y(n_547)
);

BUFx4f_ASAP7_75t_L g548 ( 
.A(n_417),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_444),
.B(n_349),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_398),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_412),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_414),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_382),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_382),
.B(n_357),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_382),
.B(n_448),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_414),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_402),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_399),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_449),
.B(n_359),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_444),
.B(n_355),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_449),
.B(n_363),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_440),
.B(n_448),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_402),
.B(n_381),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_396),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_402),
.B(n_360),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_417),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_412),
.A2(n_402),
.B1(n_417),
.B2(n_440),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_414),
.B(n_280),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_430),
.B(n_361),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_431),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_399),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_399),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_399),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_448),
.B(n_332),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_448),
.B(n_295),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_441),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_414),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_402),
.B(n_300),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_400),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_400),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_406),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_400),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_412),
.A2(n_261),
.B1(n_264),
.B2(n_275),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_400),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_430),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_396),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_412),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_404),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_402),
.B(n_159),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_412),
.B(n_324),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_412),
.B(n_328),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_404),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_406),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_417),
.B(n_159),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_419),
.B(n_259),
.C(n_195),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_396),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_404),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_482),
.B(n_314),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_525),
.B(n_507),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_457),
.A2(n_321),
.B1(n_291),
.B2(n_273),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_563),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_472),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_563),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_472),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_489),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_520),
.B(n_417),
.Y(n_608)
);

BUFx6f_ASAP7_75t_SL g609 ( 
.A(n_535),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_473),
.B(n_323),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_452),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_489),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_520),
.B(n_422),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_501),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_452),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_474),
.B(n_422),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_501),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_474),
.B(n_531),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_531),
.B(n_422),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_576),
.B(n_523),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_455),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_589),
.A2(n_551),
.B1(n_534),
.B2(n_465),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_528),
.B(n_422),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_566),
.A2(n_169),
.B1(n_168),
.B2(n_166),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_455),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_459),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_480),
.B(n_323),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_496),
.A2(n_410),
.B(n_446),
.C(n_445),
.Y(n_629)
);

AND2x4_ASAP7_75t_SL g630 ( 
.A(n_498),
.B(n_535),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_458),
.B(n_323),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_498),
.B(n_406),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_422),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_498),
.B(n_553),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_459),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_467),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_460),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_528),
.B(n_541),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_576),
.B(n_422),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_541),
.B(n_439),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_541),
.B(n_439),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_323),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_R g643 ( 
.A(n_491),
.B(n_453),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_523),
.B(n_439),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_565),
.B(n_439),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_572),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_498),
.B(n_406),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_553),
.Y(n_648)
);

O2A1O1Ixp5_ASAP7_75t_L g649 ( 
.A1(n_502),
.A2(n_511),
.B(n_513),
.C(n_504),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_553),
.B(n_406),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_565),
.B(n_439),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_460),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_565),
.B(n_439),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_504),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_588),
.B(n_598),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_588),
.B(n_416),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_542),
.B(n_559),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_468),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_468),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_495),
.B(n_160),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_588),
.B(n_416),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_467),
.B(n_469),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_560),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_598),
.B(n_552),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_598),
.B(n_416),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_553),
.B(n_416),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_511),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_513),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_534),
.B(n_419),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_567),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_519),
.B(n_416),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_487),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_487),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_554),
.B(n_416),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_555),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_524),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_564),
.B(n_524),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_503),
.B(n_160),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_469),
.B(n_161),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_555),
.A2(n_410),
.B1(n_404),
.B2(n_420),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_532),
.B(n_416),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_555),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_532),
.Y(n_683)
);

BUFx6f_ASAP7_75t_SL g684 ( 
.A(n_535),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_475),
.B(n_161),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_533),
.B(n_416),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_555),
.A2(n_410),
.B1(n_424),
.B2(n_420),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_533),
.B(n_416),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_475),
.B(n_166),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_539),
.B(n_396),
.Y(n_690)
);

BUFx5_ASAP7_75t_L g691 ( 
.A(n_567),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_539),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_544),
.B(n_556),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_544),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_556),
.B(n_420),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_514),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_514),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_570),
.B(n_420),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_570),
.B(n_420),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_579),
.B(n_420),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_464),
.B(n_410),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_464),
.B(n_420),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_L g703 ( 
.A(n_568),
.B(n_168),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_479),
.B(n_169),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_420),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_464),
.B(n_420),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_479),
.B(n_171),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_551),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_591),
.B(n_424),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_508),
.B(n_424),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_508),
.B(n_424),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_585),
.A2(n_424),
.B1(n_433),
.B2(n_427),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_562),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_515),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_454),
.B(n_424),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_515),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_481),
.B(n_424),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_461),
.B(n_171),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_454),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_562),
.B(n_419),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_560),
.B(n_172),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_454),
.B(n_424),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_481),
.B(n_424),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_572),
.B(n_163),
.Y(n_724)
);

O2A1O1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_484),
.A2(n_447),
.B(n_446),
.C(n_445),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_536),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_476),
.B(n_386),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_476),
.B(n_386),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_481),
.B(n_172),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_548),
.B(n_174),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_535),
.A2(n_304),
.B1(n_170),
.B2(n_175),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_483),
.B(n_386),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_483),
.B(n_557),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_483),
.B(n_388),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_557),
.B(n_388),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_516),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_557),
.B(n_388),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_549),
.B(n_174),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_577),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_581),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_516),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_517),
.Y(n_742)
);

AND2x6_ASAP7_75t_SL g743 ( 
.A(n_535),
.B(n_223),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_490),
.B(n_425),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_549),
.B(n_176),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_548),
.B(n_176),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_462),
.B(n_181),
.Y(n_747)
);

OAI22x1_ASAP7_75t_SL g748 ( 
.A1(n_587),
.A2(n_156),
.B1(n_304),
.B2(n_301),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_577),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_557),
.B(n_401),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_577),
.A2(n_427),
.B1(n_429),
.B2(n_433),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_537),
.B(n_181),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_548),
.B(n_183),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_540),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_577),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_505),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_580),
.B(n_401),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_589),
.B(n_401),
.Y(n_758)
);

NOR2xp67_ASAP7_75t_L g759 ( 
.A(n_486),
.B(n_425),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_571),
.B(n_447),
.C(n_446),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_L g761 ( 
.A1(n_496),
.A2(n_269),
.B1(n_170),
.B2(n_175),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_505),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_581),
.B(n_582),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_582),
.B(n_590),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_561),
.B(n_183),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_517),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_492),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_596),
.A2(n_405),
.B(n_407),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_590),
.B(n_403),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_592),
.B(n_185),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_594),
.B(n_403),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_670),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_601),
.B(n_603),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_670),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_603),
.B(n_594),
.Y(n_775)
);

NOR2xp67_ASAP7_75t_L g776 ( 
.A(n_767),
.B(n_486),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_646),
.B(n_593),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_713),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_657),
.B(n_529),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_600),
.B(n_578),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_605),
.B(n_521),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_747),
.A2(n_510),
.B(n_485),
.C(n_597),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_638),
.A2(n_488),
.B(n_451),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_754),
.B(n_578),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_605),
.B(n_521),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_682),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_644),
.A2(n_510),
.B1(n_536),
.B2(n_569),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_655),
.A2(n_488),
.B(n_451),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_644),
.A2(n_618),
.B1(n_621),
.B2(n_770),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_660),
.A2(n_485),
.B(n_597),
.C(n_512),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_675),
.A2(n_299),
.B1(n_185),
.B2(n_229),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_639),
.B(n_522),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_733),
.A2(n_664),
.B(n_671),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_639),
.B(n_522),
.Y(n_794)
);

OAI21xp5_ASAP7_75t_L g795 ( 
.A1(n_649),
.A2(n_530),
.B(n_527),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_674),
.A2(n_488),
.B(n_451),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_663),
.B(n_595),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_616),
.A2(n_530),
.B(n_527),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_656),
.A2(n_488),
.B(n_451),
.Y(n_799)
);

AND2x2_ASAP7_75t_SL g800 ( 
.A(n_724),
.B(n_244),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_703),
.A2(n_599),
.B(n_586),
.C(n_584),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_682),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_620),
.A2(n_546),
.B(n_543),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_661),
.A2(n_488),
.B(n_451),
.Y(n_804)
);

BUFx4f_ASAP7_75t_L g805 ( 
.A(n_621),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_669),
.B(n_543),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_648),
.B(n_451),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_713),
.B(n_425),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_665),
.A2(n_666),
.B(n_650),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_694),
.B(n_506),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_SL g811 ( 
.A(n_609),
.B(n_167),
.Y(n_811)
);

NOR3xp33_ASAP7_75t_L g812 ( 
.A(n_752),
.B(n_434),
.C(n_432),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_650),
.A2(n_494),
.B(n_488),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_669),
.B(n_546),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_662),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_669),
.B(n_547),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_662),
.B(n_270),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_708),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_666),
.A2(n_494),
.B(n_518),
.Y(n_819)
);

AO21x1_ASAP7_75t_L g820 ( 
.A1(n_623),
.A2(n_500),
.B(n_558),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_636),
.B(n_595),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_636),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_679),
.B(n_685),
.Y(n_823)
);

BUFx8_ASAP7_75t_SL g824 ( 
.A(n_609),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_547),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_632),
.A2(n_494),
.B(n_518),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_721),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_677),
.B(n_550),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_670),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_608),
.A2(n_599),
.B(n_558),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_611),
.B(n_550),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_624),
.A2(n_586),
.B(n_584),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_648),
.B(n_494),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_703),
.A2(n_573),
.B(n_575),
.C(n_574),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_632),
.A2(n_494),
.B(n_518),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_611),
.B(n_573),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_647),
.A2(n_494),
.B(n_518),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_720),
.B(n_432),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_617),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_648),
.B(n_518),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_615),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_622),
.B(n_574),
.Y(n_842)
);

AO21x1_ASAP7_75t_L g843 ( 
.A1(n_711),
.A2(n_500),
.B(n_575),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_622),
.B(n_456),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_647),
.A2(n_518),
.B(n_595),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_633),
.A2(n_583),
.B(n_493),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_648),
.B(n_691),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_668),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_694),
.B(n_506),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_720),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_626),
.B(n_627),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_640),
.A2(n_477),
.B(n_470),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_629),
.A2(n_447),
.B(n_432),
.C(n_434),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_641),
.A2(n_583),
.B(n_493),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_626),
.B(n_456),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_645),
.A2(n_583),
.B(n_493),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_675),
.A2(n_536),
.B1(n_569),
.B2(n_509),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_708),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_651),
.A2(n_583),
.B(n_493),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_653),
.A2(n_583),
.B(n_493),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_627),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_643),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_709),
.A2(n_545),
.B(n_538),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_607),
.B(n_463),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_668),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_629),
.A2(n_701),
.B(n_680),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_701),
.A2(n_477),
.B(n_463),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_612),
.B(n_470),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_634),
.A2(n_737),
.B(n_735),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_635),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_708),
.Y(n_871)
);

NOR2x1_ASAP7_75t_L g872 ( 
.A(n_758),
.B(n_675),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_635),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_637),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_634),
.A2(n_750),
.B(n_687),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_637),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_614),
.B(n_471),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_690),
.A2(n_545),
.B(n_538),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_670),
.A2(n_229),
.B1(n_297),
.B2(n_271),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_648),
.B(n_506),
.Y(n_880)
);

AOI21x1_ASAP7_75t_L g881 ( 
.A1(n_702),
.A2(n_471),
.B(n_478),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_652),
.B(n_478),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_738),
.B(n_434),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_744),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_619),
.A2(n_438),
.B(n_435),
.C(n_436),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_689),
.B(n_256),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_658),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_658),
.B(n_497),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_659),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_659),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_670),
.A2(n_256),
.B1(n_297),
.B2(n_271),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_702),
.A2(n_545),
.B(n_538),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_708),
.Y(n_893)
);

NOR2x1_ASAP7_75t_L g894 ( 
.A(n_610),
.B(n_435),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_745),
.B(n_270),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_654),
.A2(n_438),
.B(n_435),
.C(n_436),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_706),
.A2(n_545),
.B(n_538),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_672),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_706),
.A2(n_545),
.B(n_538),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_704),
.B(n_258),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_672),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_707),
.B(n_765),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_673),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_673),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_691),
.B(n_497),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_678),
.B(n_270),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_691),
.B(n_499),
.Y(n_907)
);

AO21x2_ASAP7_75t_L g908 ( 
.A1(n_768),
.A2(n_403),
.B(n_405),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_691),
.B(n_506),
.Y(n_909)
);

OAI21xp33_ASAP7_75t_L g910 ( 
.A1(n_718),
.A2(n_179),
.B(n_156),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_667),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_602),
.B(n_445),
.C(n_438),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_717),
.A2(n_526),
.B(n_509),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_691),
.B(n_499),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_717),
.A2(n_526),
.B(n_512),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_723),
.A2(n_526),
.B(n_427),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_723),
.A2(n_526),
.B(n_427),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_676),
.B(n_526),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_604),
.B(n_436),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_681),
.A2(n_433),
.B(n_429),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_683),
.B(n_536),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_708),
.A2(n_630),
.B1(n_692),
.B2(n_755),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_630),
.A2(n_258),
.B1(n_263),
.B2(n_266),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_686),
.A2(n_433),
.B(n_429),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_628),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_744),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_760),
.B(n_443),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_748),
.Y(n_928)
);

BUFx12f_ASAP7_75t_L g929 ( 
.A(n_743),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_691),
.B(n_536),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_691),
.B(n_536),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_613),
.A2(n_569),
.B(n_536),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_740),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_739),
.A2(n_749),
.B1(n_606),
.B2(n_693),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_740),
.B(n_569),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_757),
.B(n_569),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_729),
.A2(n_443),
.B(n_407),
.C(n_405),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_759),
.B(n_569),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_631),
.B(n_569),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_688),
.A2(n_429),
.B(n_395),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_715),
.A2(n_397),
.B(n_395),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_722),
.A2(n_397),
.B(n_395),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_729),
.A2(n_397),
.B(n_395),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_726),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_642),
.B(n_263),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_731),
.B(n_266),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_719),
.A2(n_299),
.B1(n_443),
.B2(n_209),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_625),
.B(n_167),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_763),
.A2(n_764),
.B(n_727),
.Y(n_949)
);

AO21x1_ASAP7_75t_L g950 ( 
.A1(n_730),
.A2(n_407),
.B(n_167),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_609),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_696),
.B(n_395),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_730),
.A2(n_397),
.B(n_395),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_697),
.B(n_397),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_746),
.A2(n_397),
.B(n_212),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_769),
.A2(n_119),
.B(n_144),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_746),
.A2(n_753),
.B(n_761),
.C(n_725),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_784),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_951),
.B(n_726),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_773),
.B(n_697),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_823),
.A2(n_684),
.B1(n_753),
.B2(n_762),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_850),
.B(n_756),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_902),
.A2(n_684),
.B1(n_728),
.B2(n_732),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_778),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_926),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_817),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_793),
.A2(n_751),
.B(n_734),
.Y(n_967)
);

OAI22x1_ASAP7_75t_L g968 ( 
.A1(n_780),
.A2(n_268),
.B1(n_260),
.B2(n_301),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_777),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_951),
.B(n_714),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_841),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_861),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_829),
.B(n_714),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_926),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_818),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_L g976 ( 
.A(n_886),
.B(n_286),
.C(n_220),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_805),
.B(n_716),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_R g978 ( 
.A(n_810),
.B(n_849),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_870),
.Y(n_979)
);

AOI221xp5_ASAP7_75t_L g980 ( 
.A1(n_946),
.A2(n_179),
.B1(n_180),
.B2(n_260),
.C(n_268),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_773),
.B(n_716),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_805),
.B(n_736),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_789),
.B(n_736),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_876),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_875),
.A2(n_712),
.B(n_695),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_827),
.B(n_815),
.Y(n_986)
);

INVx3_ASAP7_75t_SL g987 ( 
.A(n_862),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_930),
.A2(n_705),
.B(n_698),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_866),
.A2(n_700),
.B(n_699),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_SL g990 ( 
.A1(n_945),
.A2(n_771),
.B(n_684),
.C(n_296),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_884),
.B(n_766),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_839),
.Y(n_992)
);

OR2x2_ASAP7_75t_SL g993 ( 
.A(n_838),
.B(n_269),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_SL g994 ( 
.A(n_800),
.B(n_180),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_883),
.B(n_766),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_930),
.A2(n_742),
.B(n_741),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_931),
.A2(n_742),
.B(n_741),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_779),
.B(n_293),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_900),
.B(n_292),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_911),
.B(n_287),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_810),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_782),
.A2(n_284),
.B(n_283),
.C(n_274),
.Y(n_1002)
);

AOI221xp5_ASAP7_75t_L g1003 ( 
.A1(n_910),
.A2(n_252),
.B1(n_251),
.B2(n_247),
.C(n_246),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_822),
.B(n_240),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_848),
.B(n_234),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_808),
.Y(n_1006)
);

AOI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_957),
.A2(n_231),
.B(n_230),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_929),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_SL g1009 ( 
.A(n_906),
.B(n_8),
.C(n_9),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_925),
.B(n_8),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_847),
.A2(n_62),
.B(n_145),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_928),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_865),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_933),
.B(n_57),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_895),
.B(n_11),
.Y(n_1015)
);

INVx3_ASAP7_75t_SL g1016 ( 
.A(n_919),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_792),
.B(n_150),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_849),
.B(n_142),
.Y(n_1018)
);

OAI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_948),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_790),
.A2(n_18),
.B(n_20),
.C(n_24),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_797),
.B(n_24),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_SL g1022 ( 
.A1(n_923),
.A2(n_927),
.B1(n_944),
.B2(n_802),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_905),
.A2(n_914),
.B(n_907),
.Y(n_1023)
);

NOR2xp67_ASAP7_75t_L g1024 ( 
.A(n_776),
.B(n_66),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_829),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_919),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_792),
.B(n_65),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_824),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_905),
.A2(n_88),
.B(n_138),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_907),
.A2(n_64),
.B(n_136),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_872),
.B(n_141),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_794),
.B(n_127),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_791),
.B(n_32),
.C(n_35),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_914),
.A2(n_126),
.B(n_113),
.Y(n_1034)
);

NOR2xp67_ASAP7_75t_SL g1035 ( 
.A(n_818),
.B(n_858),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_912),
.B(n_32),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_873),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_828),
.A2(n_112),
.B(n_100),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_934),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_818),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_881),
.A2(n_97),
.B(n_92),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_811),
.B(n_39),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_828),
.A2(n_89),
.B(n_42),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_879),
.B(n_41),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_794),
.B(n_41),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_949),
.A2(n_44),
.B(n_45),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_944),
.B(n_44),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_887),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_869),
.A2(n_49),
.B(n_51),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_786),
.A2(n_812),
.B1(n_950),
.B2(n_889),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_874),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_SL g1052 ( 
.A1(n_922),
.A2(n_901),
.B(n_903),
.C(n_904),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_891),
.B(n_821),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_809),
.A2(n_787),
.B(n_936),
.C(n_853),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_SL g1055 ( 
.A1(n_935),
.A2(n_939),
.B(n_936),
.C(n_938),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_947),
.A2(n_896),
.B(n_885),
.C(n_890),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_944),
.B(n_858),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_894),
.B(n_898),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_851),
.B(n_775),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_SL g1060 ( 
.A(n_955),
.B(n_880),
.C(n_775),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_921),
.A2(n_851),
.B(n_935),
.C(n_932),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_858),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_772),
.B(n_774),
.Y(n_1063)
);

CKINVDCx8_ASAP7_75t_R g1064 ( 
.A(n_871),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_825),
.A2(n_863),
.B(n_909),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_871),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_781),
.A2(n_785),
.B1(n_871),
.B2(n_814),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_781),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_772),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_785),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_774),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_937),
.A2(n_918),
.B(n_868),
.C(n_877),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_807),
.A2(n_878),
.B(n_816),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_SL g1074 ( 
.A(n_833),
.B(n_840),
.C(n_806),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_864),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_952),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_SL g1077 ( 
.A1(n_795),
.A2(n_867),
.B(n_893),
.C(n_803),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_893),
.B(n_857),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_956),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_820),
.A2(n_843),
.B1(n_831),
.B2(n_842),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_831),
.B(n_836),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_836),
.A2(n_842),
.B(n_801),
.C(n_834),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_R g1083 ( 
.A(n_844),
.B(n_882),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_952),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_844),
.B(n_888),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_908),
.B(n_882),
.Y(n_1086)
);

OAI22x1_ASAP7_75t_L g1087 ( 
.A1(n_855),
.A2(n_888),
.B1(n_954),
.B2(n_807),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_916),
.A2(n_917),
.B(n_913),
.C(n_915),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_845),
.B(n_892),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_846),
.A2(n_860),
.B(n_856),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_920),
.A2(n_924),
.B(n_897),
.C(n_899),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_854),
.A2(n_859),
.B(n_796),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_855),
.B(n_798),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_783),
.A2(n_788),
.B(n_830),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_908),
.B(n_954),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_SL g1096 ( 
.A(n_813),
.B(n_837),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_832),
.B(n_940),
.C(n_943),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_852),
.B(n_942),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_953),
.Y(n_1099)
);

OAI22x1_ASAP7_75t_L g1100 ( 
.A1(n_941),
.A2(n_819),
.B1(n_826),
.B2(n_835),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1006),
.B(n_799),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_992),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_1007),
.A2(n_804),
.B(n_999),
.Y(n_1103)
);

NOR2x1_ASAP7_75t_R g1104 ( 
.A(n_1028),
.B(n_1008),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1054),
.A2(n_1077),
.B(n_1061),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1059),
.A2(n_967),
.B(n_1093),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1059),
.A2(n_1098),
.B(n_1082),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_SL g1108 ( 
.A1(n_1020),
.A2(n_1002),
.B(n_1014),
.C(n_1031),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1015),
.A2(n_1009),
.B(n_969),
.C(n_958),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1044),
.A2(n_1036),
.B1(n_1022),
.B2(n_998),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_964),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1023),
.A2(n_1085),
.B(n_1094),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1065),
.A2(n_985),
.B(n_1073),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1013),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1037),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1092),
.A2(n_1090),
.B(n_996),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_SL g1117 ( 
.A(n_1064),
.B(n_1019),
.Y(n_1117)
);

INVxp33_ASAP7_75t_L g1118 ( 
.A(n_986),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_974),
.B(n_966),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_997),
.A2(n_1041),
.B(n_988),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1052),
.A2(n_1080),
.B(n_989),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1007),
.A2(n_968),
.B1(n_1042),
.B2(n_980),
.C(n_1039),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1055),
.A2(n_1081),
.B(n_1072),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_1087),
.A2(n_1091),
.A3(n_1088),
.B(n_1100),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_1035),
.B(n_1025),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1051),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1053),
.A2(n_1021),
.B(n_1046),
.C(n_976),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_989),
.A2(n_1095),
.B(n_1086),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1067),
.A2(n_1095),
.B(n_1027),
.Y(n_1130)
);

AOI221x1_ASAP7_75t_L g1131 ( 
.A1(n_1049),
.A2(n_1043),
.B1(n_1097),
.B2(n_1067),
.C(n_1045),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_1066),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1010),
.A2(n_994),
.B(n_1033),
.C(n_1005),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_SL g1134 ( 
.A1(n_1014),
.A2(n_1045),
.B(n_1027),
.C(n_1017),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_963),
.A2(n_965),
.B1(n_1016),
.B2(n_1012),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1017),
.A2(n_1032),
.B(n_983),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_962),
.B(n_1026),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_971),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_972),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1032),
.A2(n_983),
.B(n_982),
.C(n_977),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_979),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_984),
.Y(n_1142)
);

OA21x2_ASAP7_75t_L g1143 ( 
.A1(n_1050),
.A2(n_1060),
.B(n_960),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_994),
.B(n_961),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1069),
.Y(n_1145)
);

AO22x2_ASAP7_75t_L g1146 ( 
.A1(n_1078),
.A2(n_1075),
.B1(n_995),
.B2(n_1005),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_960),
.A2(n_981),
.B(n_973),
.Y(n_1147)
);

AND3x2_ASAP7_75t_L g1148 ( 
.A(n_1047),
.B(n_1018),
.C(n_959),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_1047),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_1062),
.Y(n_1150)
);

AO22x2_ASAP7_75t_L g1151 ( 
.A1(n_1078),
.A2(n_1018),
.B1(n_1004),
.B2(n_970),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1048),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_SL g1153 ( 
.A1(n_1076),
.A2(n_1057),
.B(n_1056),
.C(n_991),
.Y(n_1153)
);

INVx3_ASAP7_75t_SL g1154 ( 
.A(n_987),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_978),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1089),
.A2(n_1096),
.B(n_1099),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1069),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_990),
.A2(n_1011),
.B(n_1029),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_1066),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_959),
.B(n_1001),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1084),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1058),
.A2(n_1038),
.A3(n_1030),
.B(n_1034),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_970),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1066),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1071),
.A2(n_1025),
.B(n_1001),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1083),
.B(n_1063),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1069),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1089),
.A2(n_1096),
.B(n_1079),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1063),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_975),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1074),
.A2(n_1089),
.B(n_1024),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1000),
.A2(n_1003),
.B1(n_1040),
.B2(n_993),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_SL g1173 ( 
.A(n_1040),
.B(n_600),
.C(n_823),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1079),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1079),
.B(n_1068),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1069),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1087),
.A2(n_820),
.A3(n_1054),
.B(n_950),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1059),
.A2(n_648),
.B(n_967),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_992),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1080),
.A2(n_1094),
.B(n_1090),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1039),
.A2(n_782),
.B1(n_1019),
.B2(n_1046),
.C(n_1020),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_992),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_1046),
.A2(n_823),
.B(n_601),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1069),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_SL g1187 ( 
.A1(n_1046),
.A2(n_1014),
.B(n_1056),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1015),
.A2(n_823),
.B1(n_747),
.B2(n_600),
.C(n_602),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_964),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_992),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1059),
.A2(n_648),
.B(n_967),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1073),
.A2(n_1092),
.B(n_1090),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1059),
.A2(n_648),
.B(n_967),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1073),
.A2(n_1092),
.B(n_1090),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1087),
.A2(n_820),
.A3(n_1054),
.B(n_950),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_987),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1062),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1069),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_998),
.Y(n_1199)
);

AOI21xp33_ASAP7_75t_L g1200 ( 
.A1(n_1007),
.A2(n_823),
.B(n_601),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1054),
.A2(n_1077),
.B(n_1061),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_992),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1006),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1087),
.A2(n_820),
.A3(n_1054),
.B(n_950),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1015),
.B(n_823),
.C(n_886),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1006),
.B(n_646),
.Y(n_1206)
);

BUFx8_ASAP7_75t_L g1207 ( 
.A(n_1008),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1059),
.A2(n_648),
.B(n_967),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1087),
.A2(n_820),
.A3(n_1054),
.B(n_950),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_992),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_964),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1015),
.A2(n_823),
.B(n_601),
.C(n_902),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_992),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1214)
);

BUFx8_ASAP7_75t_L g1215 ( 
.A(n_1008),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1015),
.A2(n_823),
.B(n_601),
.C(n_902),
.Y(n_1216)
);

AOI31xp67_ASAP7_75t_L g1217 ( 
.A1(n_1080),
.A2(n_1098),
.A3(n_963),
.B(n_1031),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1015),
.A2(n_823),
.B1(n_902),
.B2(n_900),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1015),
.A2(n_823),
.B(n_601),
.C(n_902),
.Y(n_1219)
);

BUFx8_ASAP7_75t_L g1220 ( 
.A(n_1008),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1062),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_969),
.B(n_958),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_969),
.B(n_958),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1059),
.A2(n_926),
.B1(n_601),
.B2(n_823),
.Y(n_1224)
);

BUFx12f_ASAP7_75t_L g1225 ( 
.A(n_1008),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_959),
.B(n_974),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_992),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1059),
.A2(n_648),
.B(n_967),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1059),
.A2(n_648),
.B(n_967),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1008),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1066),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1062),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_969),
.B(n_958),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1054),
.A2(n_1077),
.B(n_1061),
.Y(n_1235)
);

BUFx2_ASAP7_75t_R g1236 ( 
.A(n_1028),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1062),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1110),
.A2(n_1205),
.B1(n_1188),
.B2(n_1122),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1188),
.A2(n_1205),
.B1(n_1122),
.B2(n_1218),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1110),
.A2(n_1216),
.B1(n_1212),
.B2(n_1219),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1197),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1221),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1190),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1146),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1207),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1200),
.A2(n_1144),
.B1(n_1184),
.B2(n_1199),
.Y(n_1246)
);

BUFx12f_ASAP7_75t_L g1247 ( 
.A(n_1207),
.Y(n_1247)
);

CKINVDCx11_ASAP7_75t_R g1248 ( 
.A(n_1225),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1163),
.B(n_1165),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1137),
.B(n_1222),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1206),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1199),
.A2(n_1224),
.B1(n_1149),
.B2(n_1155),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1200),
.A2(n_1224),
.B1(n_1173),
.B2(n_1187),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1227),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1117),
.A2(n_1146),
.B1(n_1135),
.B2(n_1172),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1233),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1102),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1142),
.Y(n_1258)
);

INVx6_ASAP7_75t_L g1259 ( 
.A(n_1226),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1118),
.A2(n_1166),
.B1(n_1203),
.B2(n_1226),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1237),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1172),
.A2(n_1121),
.B1(n_1161),
.B2(n_1235),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_SL g1263 ( 
.A1(n_1151),
.A2(n_1143),
.B1(n_1235),
.B2(n_1201),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1114),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1151),
.A2(n_1101),
.B1(n_1203),
.B2(n_1223),
.Y(n_1265)
);

BUFx8_ASAP7_75t_L g1266 ( 
.A(n_1231),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1183),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1234),
.A2(n_1128),
.B1(n_1182),
.B2(n_1166),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1121),
.A2(n_1201),
.B1(n_1105),
.B2(n_1143),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1154),
.Y(n_1270)
);

INVx4_ASAP7_75t_L g1271 ( 
.A(n_1167),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1150),
.B(n_1111),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1105),
.A2(n_1107),
.B1(n_1148),
.B2(n_1180),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1112),
.A2(n_1156),
.B(n_1113),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1202),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1210),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1182),
.A2(n_1119),
.B1(n_1196),
.B2(n_1169),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1189),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1213),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1211),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1215),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1115),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1171),
.A2(n_1228),
.B1(n_1186),
.B2(n_1180),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1126),
.A2(n_1228),
.B1(n_1214),
.B2(n_1186),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1171),
.A2(n_1126),
.B1(n_1214),
.B2(n_1181),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1109),
.A2(n_1133),
.B1(n_1127),
.B2(n_1175),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1175),
.A2(n_1152),
.B1(n_1141),
.B2(n_1139),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1157),
.A2(n_1138),
.B1(n_1145),
.B2(n_1198),
.Y(n_1288)
);

INVx11_ASAP7_75t_L g1289 ( 
.A(n_1215),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1103),
.A2(n_1129),
.B1(n_1123),
.B2(n_1106),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1220),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1136),
.A2(n_1160),
.B1(n_1208),
.B2(n_1193),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1153),
.B(n_1160),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1131),
.A2(n_1160),
.B1(n_1125),
.B2(n_1191),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1145),
.B(n_1176),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1220),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1174),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1236),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1178),
.A2(n_1229),
.B1(n_1230),
.B2(n_1130),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1125),
.A2(n_1168),
.B1(n_1170),
.B2(n_1198),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1147),
.A2(n_1185),
.B1(n_1158),
.B2(n_1164),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1132),
.A2(n_1232),
.B1(n_1159),
.B2(n_1108),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1132),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1236),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1159),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1232),
.A2(n_1116),
.B1(n_1194),
.B2(n_1192),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1217),
.A2(n_1120),
.B1(n_1134),
.B2(n_1140),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1124),
.Y(n_1308)
);

INVx6_ASAP7_75t_L g1309 ( 
.A(n_1104),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1177),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1162),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1177),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1195),
.A2(n_1204),
.B1(n_1209),
.B2(n_1162),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1195),
.A2(n_1110),
.B1(n_1205),
.B2(n_601),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1204),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1209),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1137),
.B(n_1161),
.Y(n_1317)
);

OAI22x1_ASAP7_75t_L g1318 ( 
.A1(n_1110),
.A2(n_1205),
.B1(n_1144),
.B2(n_1172),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1207),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1179),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1179),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1188),
.A2(n_1205),
.B1(n_1122),
.B2(n_823),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_SL g1323 ( 
.A(n_1197),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1179),
.Y(n_1324)
);

BUFx2_ASAP7_75t_SL g1325 ( 
.A(n_1197),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1188),
.A2(n_600),
.B(n_1110),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1188),
.A2(n_1205),
.B1(n_1122),
.B2(n_823),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1110),
.A2(n_1205),
.B1(n_601),
.B2(n_1047),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1179),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1218),
.A2(n_1205),
.B1(n_600),
.B2(n_1110),
.Y(n_1330)
);

INVx8_ASAP7_75t_L g1331 ( 
.A(n_1160),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1161),
.B(n_1203),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1197),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1149),
.A2(n_1042),
.B1(n_600),
.B2(n_747),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1226),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1206),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1179),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1218),
.A2(n_1205),
.B1(n_600),
.B2(n_1110),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1179),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1218),
.A2(n_1205),
.B1(n_600),
.B2(n_1110),
.Y(n_1340)
);

BUFx2_ASAP7_75t_SL g1341 ( 
.A(n_1197),
.Y(n_1341)
);

BUFx5_ASAP7_75t_L g1342 ( 
.A(n_1174),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1218),
.A2(n_1205),
.B1(n_600),
.B2(n_1110),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1205),
.A2(n_600),
.B1(n_724),
.B2(n_1042),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1188),
.A2(n_1205),
.B1(n_1122),
.B2(n_823),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1188),
.A2(n_1205),
.B1(n_1122),
.B2(n_823),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1110),
.A2(n_1205),
.B1(n_601),
.B2(n_1047),
.Y(n_1347)
);

BUFx5_ASAP7_75t_L g1348 ( 
.A(n_1174),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1167),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1179),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1167),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1179),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1316),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1315),
.Y(n_1354)
);

AND2x4_ASAP7_75t_SL g1355 ( 
.A(n_1273),
.B(n_1244),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1310),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1326),
.A2(n_1334),
.B(n_1344),
.C(n_1327),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1274),
.A2(n_1299),
.B(n_1307),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1312),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1308),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1308),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1331),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1311),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1257),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1330),
.A2(n_1343),
.B1(n_1340),
.B2(n_1338),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1244),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1313),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1264),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1267),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1270),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1299),
.A2(n_1307),
.B(n_1306),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1275),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1306),
.A2(n_1292),
.B(n_1301),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1263),
.B(n_1262),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1292),
.A2(n_1301),
.B(n_1290),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1251),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1276),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1322),
.B(n_1345),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1279),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1332),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1336),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1331),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1283),
.B(n_1253),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1282),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1240),
.A2(n_1290),
.B(n_1294),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1345),
.B(n_1346),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1294),
.A2(n_1314),
.B(n_1238),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1283),
.B(n_1253),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1331),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1238),
.A2(n_1346),
.B(n_1347),
.C(n_1328),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1249),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1297),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1285),
.B(n_1268),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1293),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1317),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1344),
.B(n_1239),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1342),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1285),
.B(n_1246),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1287),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1246),
.B(n_1318),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1286),
.A2(n_1352),
.B(n_1350),
.Y(n_1403)
);

AND2x4_ASAP7_75t_SL g1404 ( 
.A(n_1273),
.B(n_1284),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1288),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1342),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1287),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1243),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1314),
.A2(n_1328),
.B(n_1347),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1325),
.B(n_1341),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1342),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1254),
.B(n_1329),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1265),
.B(n_1284),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1259),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1320),
.B(n_1324),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1321),
.Y(n_1416)
);

BUFx12f_ASAP7_75t_L g1417 ( 
.A(n_1296),
.Y(n_1417)
);

OAI211xp5_ASAP7_75t_L g1418 ( 
.A1(n_1239),
.A2(n_1255),
.B(n_1252),
.C(n_1277),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1255),
.A2(n_1337),
.B(n_1339),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1280),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1348),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1247),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1245),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1250),
.B(n_1252),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1258),
.B(n_1260),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1295),
.B(n_1303),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1281),
.Y(n_1427)
);

AOI21xp33_ASAP7_75t_L g1428 ( 
.A1(n_1300),
.A2(n_1302),
.B(n_1272),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1305),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1259),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1302),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1259),
.B(n_1335),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1374),
.B(n_1242),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1374),
.B(n_1261),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1365),
.A2(n_1241),
.B(n_1278),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1370),
.A2(n_1304),
.B1(n_1298),
.B2(n_1291),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1354),
.B(n_1396),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1382),
.B(n_1256),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1354),
.B(n_1351),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1364),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_SL g1441 ( 
.A(n_1410),
.B(n_1319),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1383),
.B(n_1333),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1392),
.A2(n_1387),
.B(n_1357),
.C(n_1404),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1394),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1425),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1404),
.A2(n_1398),
.B(n_1418),
.C(n_1385),
.Y(n_1446)
);

NAND2x1_ASAP7_75t_L g1447 ( 
.A(n_1410),
.B(n_1335),
.Y(n_1447)
);

AO32x2_ASAP7_75t_L g1448 ( 
.A1(n_1405),
.A2(n_1391),
.A3(n_1389),
.B1(n_1414),
.B2(n_1430),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1410),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1380),
.A2(n_1323),
.B(n_1309),
.C(n_1266),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1354),
.B(n_1349),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1354),
.B(n_1271),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1368),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1425),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1389),
.A2(n_1271),
.B(n_1323),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1397),
.B(n_1309),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1417),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1389),
.A2(n_1309),
.B(n_1266),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1396),
.B(n_1289),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1424),
.B(n_1248),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1395),
.B(n_1376),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1395),
.B(n_1376),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1388),
.A2(n_1428),
.B(n_1373),
.C(n_1385),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1364),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_SL g1465 ( 
.A(n_1378),
.B(n_1424),
.C(n_1402),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1369),
.B(n_1372),
.Y(n_1466)
);

O2A1O1Ixp5_ASAP7_75t_L g1467 ( 
.A1(n_1390),
.A2(n_1373),
.B(n_1403),
.C(n_1400),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1390),
.A2(n_1402),
.B(n_1377),
.Y(n_1468)
);

OAI21xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1400),
.A2(n_1405),
.B(n_1419),
.Y(n_1469)
);

AO32x2_ASAP7_75t_L g1470 ( 
.A1(n_1391),
.A2(n_1430),
.A3(n_1414),
.B1(n_1366),
.B2(n_1409),
.Y(n_1470)
);

NOR2x1_ASAP7_75t_SL g1471 ( 
.A(n_1403),
.B(n_1401),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1404),
.A2(n_1413),
.B1(n_1396),
.B2(n_1355),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1355),
.A2(n_1413),
.B(n_1377),
.C(n_1401),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1409),
.A2(n_1407),
.B1(n_1431),
.B2(n_1367),
.C(n_1355),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1366),
.B(n_1379),
.Y(n_1475)
);

AO32x2_ASAP7_75t_L g1476 ( 
.A1(n_1409),
.A2(n_1367),
.A3(n_1356),
.B1(n_1359),
.B2(n_1361),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1381),
.B(n_1372),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1407),
.B(n_1420),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_SL g1479 ( 
.A(n_1393),
.B(n_1360),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1358),
.A2(n_1411),
.B(n_1421),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1386),
.B(n_1399),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1444),
.B(n_1386),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1481),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1453),
.Y(n_1484)
);

INVx8_ASAP7_75t_L g1485 ( 
.A(n_1459),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1481),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1471),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1443),
.B(n_1426),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1449),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1465),
.A2(n_1415),
.B1(n_1412),
.B2(n_1417),
.Y(n_1490)
);

NOR2xp67_ASAP7_75t_L g1491 ( 
.A(n_1449),
.B(n_1429),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1475),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1440),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1470),
.B(n_1375),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1466),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1443),
.A2(n_1432),
.B1(n_1415),
.B2(n_1412),
.Y(n_1496)
);

NOR2x1_ASAP7_75t_SL g1497 ( 
.A(n_1472),
.B(n_1406),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1470),
.B(n_1375),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1464),
.Y(n_1499)
);

OAI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1446),
.A2(n_1384),
.B1(n_1362),
.B2(n_1416),
.C(n_1408),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1468),
.B(n_1353),
.Y(n_1501)
);

INVxp67_ASAP7_75t_SL g1502 ( 
.A(n_1479),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1470),
.B(n_1371),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_1478),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1470),
.B(n_1371),
.Y(n_1505)
);

NOR2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1447),
.B(n_1384),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1457),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1448),
.B(n_1363),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1448),
.B(n_1363),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1508),
.B(n_1445),
.Y(n_1511)
);

AND2x2_ASAP7_75t_SL g1512 ( 
.A(n_1494),
.B(n_1474),
.Y(n_1512)
);

NOR2xp67_ASAP7_75t_L g1513 ( 
.A(n_1500),
.B(n_1469),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1508),
.B(n_1448),
.Y(n_1514)
);

INVx5_ASAP7_75t_L g1515 ( 
.A(n_1503),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1508),
.B(n_1448),
.Y(n_1516)
);

OAI222xp33_ASAP7_75t_L g1517 ( 
.A1(n_1500),
.A2(n_1463),
.B1(n_1458),
.B2(n_1461),
.C1(n_1462),
.C2(n_1455),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1504),
.B(n_1461),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1496),
.B(n_1450),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1509),
.B(n_1454),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1509),
.B(n_1477),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1493),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1489),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1509),
.B(n_1476),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1497),
.A2(n_1473),
.A3(n_1480),
.B(n_1411),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1494),
.B(n_1476),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1507),
.B(n_1460),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1494),
.B(n_1498),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1498),
.B(n_1486),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1502),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1488),
.A2(n_1462),
.B1(n_1460),
.B2(n_1434),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1504),
.B(n_1478),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1502),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1488),
.B(n_1442),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1487),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1499),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1499),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1515),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1523),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1515),
.B(n_1523),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1512),
.B(n_1492),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1515),
.B(n_1528),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1512),
.B(n_1492),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1528),
.B(n_1515),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1528),
.B(n_1497),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1515),
.B(n_1486),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1515),
.B(n_1487),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1515),
.B(n_1514),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1522),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1537),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1503),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1514),
.B(n_1505),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1537),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1530),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1516),
.B(n_1524),
.Y(n_1557)
);

NOR3xp33_ASAP7_75t_SL g1558 ( 
.A(n_1517),
.B(n_1457),
.C(n_1427),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1511),
.B(n_1501),
.Y(n_1559)
);

NAND2x1_ASAP7_75t_L g1560 ( 
.A(n_1530),
.B(n_1491),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1532),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1510),
.B(n_1486),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1512),
.B(n_1495),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1524),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1538),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1511),
.B(n_1520),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1524),
.B(n_1505),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1523),
.B(n_1506),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1511),
.B(n_1501),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1510),
.B(n_1486),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1510),
.B(n_1483),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1526),
.B(n_1505),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1520),
.B(n_1521),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1535),
.B(n_1527),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1518),
.B(n_1495),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1568),
.B(n_1533),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1568),
.B(n_1533),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1518),
.Y(n_1579)
);

OAI21xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1542),
.A2(n_1513),
.B(n_1519),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1568),
.B(n_1546),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1550),
.Y(n_1582)
);

OAI33xp33_ASAP7_75t_L g1583 ( 
.A1(n_1561),
.A2(n_1532),
.A3(n_1482),
.B1(n_1520),
.B2(n_1438),
.B3(n_1484),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1550),
.Y(n_1584)
);

NAND2x1p5_ASAP7_75t_L g1585 ( 
.A(n_1540),
.B(n_1513),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1568),
.B(n_1536),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1544),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1572),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1572),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1546),
.B(n_1536),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1544),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1541),
.B(n_1523),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1541),
.B(n_1523),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1558),
.A2(n_1446),
.B1(n_1496),
.B2(n_1490),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1541),
.B(n_1523),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1541),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1561),
.B(n_1563),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1539),
.B(n_1525),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1574),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1555),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1523),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1540),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1540),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1558),
.A2(n_1517),
.B(n_1531),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1575),
.A2(n_1441),
.B(n_1531),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1556),
.B(n_1526),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1563),
.B(n_1521),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1559),
.B(n_1521),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1551),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1559),
.B(n_1529),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1576),
.B(n_1526),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1551),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1576),
.B(n_1534),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1555),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1554),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1556),
.B(n_1543),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1540),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1591),
.B(n_1571),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1579),
.B(n_1574),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1614),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1587),
.B(n_1571),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1585),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1609),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1616),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1609),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1601),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_SL g1628 ( 
.A(n_1580),
.B(n_1540),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1601),
.B(n_1557),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1600),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1580),
.B(n_1562),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1596),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1612),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1540),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1612),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1570),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1615),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1616),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1599),
.B(n_1570),
.Y(n_1641)
);

AND2x2_ASAP7_75t_SL g1642 ( 
.A(n_1594),
.B(n_1540),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1599),
.B(n_1433),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1579),
.B(n_1566),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1596),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1615),
.Y(n_1646)
);

AO21x2_ASAP7_75t_L g1647 ( 
.A1(n_1617),
.A2(n_1549),
.B(n_1548),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1602),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1592),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1604),
.A2(n_1467),
.B(n_1560),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1599),
.B(n_1433),
.Y(n_1651)
);

INVxp33_ASAP7_75t_L g1652 ( 
.A(n_1604),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1585),
.B(n_1434),
.Y(n_1653)
);

OAI211xp5_ASAP7_75t_L g1654 ( 
.A1(n_1630),
.A2(n_1650),
.B(n_1621),
.C(n_1637),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1624),
.Y(n_1655)
);

NAND4xp25_ASAP7_75t_L g1656 ( 
.A(n_1628),
.B(n_1594),
.C(n_1605),
.D(n_1595),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1652),
.B(n_1422),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1642),
.A2(n_1585),
.B(n_1592),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1631),
.A2(n_1595),
.B(n_1593),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1630),
.A2(n_1583),
.B1(n_1582),
.B2(n_1584),
.C(n_1589),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1629),
.B(n_1581),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1649),
.B(n_1607),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1649),
.B(n_1607),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1645),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1624),
.Y(n_1665)
);

AOI211x1_ASAP7_75t_L g1666 ( 
.A1(n_1653),
.A2(n_1581),
.B(n_1578),
.C(n_1586),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1642),
.B(n_1577),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1642),
.A2(n_1593),
.B1(n_1578),
.B2(n_1586),
.Y(n_1668)
);

AOI33xp33_ASAP7_75t_L g1669 ( 
.A1(n_1627),
.A2(n_1577),
.A3(n_1582),
.B1(n_1589),
.B2(n_1584),
.B3(n_1588),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1629),
.B(n_1590),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1627),
.B(n_1590),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1628),
.B(n_1588),
.C(n_1603),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1625),
.A2(n_1539),
.B1(n_1618),
.B2(n_1435),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1625),
.B(n_1606),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1632),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1632),
.Y(n_1676)
);

OAI322xp33_ASAP7_75t_L g1677 ( 
.A1(n_1644),
.A2(n_1588),
.A3(n_1610),
.B1(n_1608),
.B2(n_1618),
.C1(n_1613),
.C2(n_1611),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1640),
.A2(n_1548),
.B1(n_1560),
.B2(n_1539),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1656),
.A2(n_1623),
.B1(n_1640),
.B2(n_1634),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1655),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1664),
.B(n_1648),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1669),
.B(n_1648),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1654),
.A2(n_1636),
.B1(n_1651),
.B2(n_1643),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_SL g1684 ( 
.A(n_1654),
.B(n_1647),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1675),
.B(n_1644),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1657),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1665),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1662),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1660),
.A2(n_1620),
.B1(n_1622),
.B2(n_1619),
.C(n_1638),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1659),
.B(n_1423),
.Y(n_1690)
);

OAI21xp33_ASAP7_75t_L g1691 ( 
.A1(n_1668),
.A2(n_1641),
.B(n_1620),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1658),
.B(n_1634),
.Y(n_1692)
);

O2A1O1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1672),
.A2(n_1603),
.B(n_1646),
.C(n_1639),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1667),
.B(n_1436),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1661),
.B(n_1671),
.Y(n_1695)
);

AND3x1_ASAP7_75t_L g1696 ( 
.A(n_1660),
.B(n_1633),
.C(n_1626),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1670),
.A2(n_1548),
.B1(n_1647),
.B2(n_1639),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1684),
.Y(n_1698)
);

AOI222xp33_ASAP7_75t_L g1699 ( 
.A1(n_1682),
.A2(n_1673),
.B1(n_1675),
.B2(n_1676),
.C1(n_1674),
.C2(n_1646),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1685),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1695),
.B(n_1688),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1696),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1681),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1694),
.A2(n_1673),
.B1(n_1663),
.B2(n_1678),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1680),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1693),
.B(n_1666),
.C(n_1633),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1690),
.B(n_1606),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1687),
.Y(n_1708)
);

NOR2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1701),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1707),
.B(n_1694),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1703),
.Y(n_1712)
);

NAND4xp25_ASAP7_75t_L g1713 ( 
.A(n_1699),
.B(n_1691),
.C(n_1683),
.D(n_1692),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1702),
.A2(n_1689),
.B1(n_1679),
.B2(n_1697),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1702),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1707),
.B(n_1679),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1698),
.B(n_1626),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_R g1718 ( 
.A(n_1712),
.B(n_1710),
.Y(n_1718)
);

OAI211xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1714),
.A2(n_1698),
.B(n_1704),
.C(n_1706),
.Y(n_1719)
);

NAND4xp25_ASAP7_75t_L g1720 ( 
.A(n_1713),
.B(n_1708),
.C(n_1705),
.D(n_1635),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1716),
.A2(n_1647),
.B1(n_1635),
.B2(n_1548),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1715),
.B(n_1611),
.Y(n_1722)
);

O2A1O1Ixp5_ASAP7_75t_SL g1723 ( 
.A1(n_1722),
.A2(n_1717),
.B(n_1709),
.C(n_1711),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1719),
.A2(n_1677),
.B1(n_1598),
.B2(n_1506),
.Y(n_1724)
);

OAI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1718),
.A2(n_1613),
.B(n_1549),
.C(n_1490),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1721),
.A2(n_1598),
.B1(n_1549),
.B2(n_1608),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1720),
.A2(n_1598),
.B1(n_1552),
.B2(n_1543),
.C(n_1545),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1719),
.A2(n_1598),
.B1(n_1459),
.B2(n_1543),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1725),
.B(n_1610),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1728),
.B(n_1545),
.Y(n_1730)
);

AO22x2_ASAP7_75t_L g1731 ( 
.A1(n_1726),
.A2(n_1552),
.B1(n_1564),
.B2(n_1557),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1724),
.A2(n_1459),
.B1(n_1452),
.B2(n_1439),
.Y(n_1732)
);

NOR2x1_ASAP7_75t_L g1733 ( 
.A(n_1723),
.B(n_1552),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1729),
.A2(n_1727),
.B(n_1456),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1733),
.B(n_1554),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1730),
.B(n_1565),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1735),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1737),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1738),
.A2(n_1736),
.B(n_1734),
.C(n_1732),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1738),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1731),
.B1(n_1566),
.B2(n_1564),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1739),
.A2(n_1564),
.B1(n_1569),
.B2(n_1567),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1547),
.B1(n_1553),
.B2(n_1573),
.Y(n_1743)
);

OAI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1569),
.B1(n_1565),
.B2(n_1529),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1744),
.B(n_1553),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1743),
.B(n_1439),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1746),
.Y(n_1747)
);

OAI221xp5_ASAP7_75t_R g1748 ( 
.A1(n_1747),
.A2(n_1485),
.B1(n_1525),
.B2(n_1573),
.C(n_1567),
.Y(n_1748)
);

AOI211xp5_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1452),
.B(n_1451),
.C(n_1439),
.Y(n_1749)
);


endmodule