module fake_jpeg_16575_n_92 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_2),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_2),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_36),
.Y(n_44)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_1),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_38),
.B(n_32),
.C(n_31),
.Y(n_48)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_54),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_35),
.B1(n_33),
.B2(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_53),
.B1(n_56),
.B2(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_46),
.B1(n_18),
.B2(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_17),
.B1(n_21),
.B2(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_28),
.Y(n_78)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_78),
.C(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_79),
.B(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_63),
.C(n_62),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_83),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_61),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_84),
.B1(n_77),
.B2(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_63),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_88),
.B(n_74),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_80),
.C(n_73),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_25),
.Y(n_91)
);

XNOR2x2_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_26),
.Y(n_92)
);


endmodule