module real_jpeg_32745_n_27 (n_17, n_199, n_8, n_0, n_21, n_2, n_196, n_191, n_10, n_9, n_12, n_24, n_6, n_190, n_194, n_192, n_198, n_23, n_11, n_14, n_25, n_195, n_7, n_22, n_18, n_3, n_193, n_197, n_5, n_4, n_1, n_26, n_200, n_20, n_19, n_16, n_15, n_13, n_27);

input n_17;
input n_199;
input n_8;
input n_0;
input n_21;
input n_2;
input n_196;
input n_191;
input n_10;
input n_9;
input n_12;
input n_24;
input n_6;
input n_190;
input n_194;
input n_192;
input n_198;
input n_23;
input n_11;
input n_14;
input n_25;
input n_195;
input n_7;
input n_22;
input n_18;
input n_3;
input n_193;
input n_197;
input n_5;
input n_4;
input n_1;
input n_26;
input n_200;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI221xp5_ASAP7_75t_SL g125 ( 
.A1(n_0),
.A2(n_2),
.B1(n_126),
.B2(n_130),
.C(n_131),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_0),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_1),
.B(n_109),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_126),
.C(n_130),
.Y(n_134)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_4),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_79),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_6),
.B(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_9),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_9),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_10),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_68),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_12),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_13),
.B(n_86),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_14),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_15),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_16),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_17),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_17),
.B(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_18),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_20),
.A2(n_41),
.B1(n_43),
.B2(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_21),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_21),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_24),
.B(n_72),
.Y(n_186)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_25),
.A2(n_99),
.A3(n_101),
.B1(n_107),
.B2(n_160),
.C1(n_162),
.C2(n_200),
.Y(n_159)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_92),
.B(n_165),
.Y(n_39)
);

NAND4xp25_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_54),
.C(n_77),
.D(n_84),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_50),
.Y(n_153)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_66),
.C(n_70),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_56),
.B(n_177),
.C(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_65),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_57),
.B(n_65),
.Y(n_181)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp67_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_73),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_74),
.Y(n_185)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_196),
.Y(n_130)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_77),
.B(n_168),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_77),
.A2(n_183),
.B(n_187),
.Y(n_182)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI221xp5_ASAP7_75t_L g166 ( 
.A1(n_78),
.A2(n_167),
.B1(n_179),
.B2(n_180),
.C(n_182),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

AOI31xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_118),
.A3(n_148),
.B(n_155),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_106),
.C(n_113),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_156),
.B(n_159),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_113),
.C(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_191),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

OA21x2_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_143),
.C(n_144),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_135),
.B(n_142),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_125),
.B1(n_133),
.B2(n_134),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_141),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B(n_172),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_190),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_192),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_193),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_194),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_195),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_197),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_198),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_199),
.Y(n_151)
);


endmodule