module real_aes_10335_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_0), .Y(n_789) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_1), .A2(n_145), .B1(n_1415), .B2(n_1482), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_2), .A2(n_9), .B1(n_665), .B2(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1500 ( .A(n_2), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_3), .A2(n_219), .B1(n_927), .B2(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g940 ( .A(n_3), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_4), .A2(n_207), .B1(n_957), .B2(n_959), .Y(n_956) );
INVx1_ASAP7_75t_L g1004 ( .A(n_4), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_5), .A2(n_66), .B1(n_1196), .B2(n_1212), .Y(n_1219) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_6), .Y(n_809) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_7), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_7), .B(n_186), .Y(n_384) );
AND2x2_ASAP7_75t_L g394 ( .A(n_7), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g422 ( .A(n_7), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_8), .A2(n_154), .B1(n_346), .B2(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g448 ( .A(n_8), .Y(n_448) );
INVx1_ASAP7_75t_L g1501 ( .A(n_9), .Y(n_1501) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_10), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_10), .A2(n_239), .B1(n_747), .B2(n_749), .C(n_750), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_11), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g968 ( .A(n_12), .Y(n_968) );
INVx1_ASAP7_75t_L g901 ( .A(n_13), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_13), .A2(n_74), .B1(n_937), .B2(n_938), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g1404 ( .A1(n_14), .A2(n_1405), .B1(n_1444), .B2(n_1445), .Y(n_1404) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_14), .Y(n_1444) );
INVxp33_ASAP7_75t_SL g697 ( .A(n_15), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_15), .A2(n_77), .B1(n_672), .B2(n_734), .C(n_736), .Y(n_733) );
CKINVDCx5p33_ASAP7_75t_R g1463 ( .A(n_16), .Y(n_1463) );
XNOR2x2_ASAP7_75t_L g1026 ( .A(n_17), .B(n_1027), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_17), .A2(n_75), .B1(n_1192), .B2(n_1196), .Y(n_1203) );
AOI21xp33_ASAP7_75t_L g1043 ( .A1(n_18), .A2(n_508), .B(n_509), .Y(n_1043) );
INVx1_ASAP7_75t_L g1066 ( .A(n_18), .Y(n_1066) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_19), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_20), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g825 ( .A(n_21), .B(n_826), .Y(n_825) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_22), .A2(n_88), .B1(n_597), .B2(n_604), .C(n_607), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_22), .A2(n_88), .B1(n_657), .B2(n_660), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_23), .A2(n_47), .B1(n_973), .B2(n_975), .Y(n_972) );
INVx1_ASAP7_75t_L g1021 ( .A(n_23), .Y(n_1021) );
INVx1_ASAP7_75t_L g1092 ( .A(n_24), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_24), .A2(n_183), .B1(n_555), .B2(n_931), .Y(n_1114) );
OR2x2_ASAP7_75t_L g290 ( .A(n_25), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g329 ( .A(n_25), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_26), .A2(n_161), .B1(n_1051), .B2(n_1052), .Y(n_1050) );
INVx1_ASAP7_75t_L g1062 ( .A(n_26), .Y(n_1062) );
CKINVDCx5p33_ASAP7_75t_R g1045 ( .A(n_27), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_28), .A2(n_136), .B1(n_1180), .B2(n_1188), .Y(n_1202) );
INVx1_ASAP7_75t_L g491 ( .A(n_29), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_29), .A2(n_168), .B1(n_558), .B2(n_561), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_30), .Y(n_318) );
INVx1_ASAP7_75t_L g755 ( .A(n_31), .Y(n_755) );
INVx1_ASAP7_75t_L g292 ( .A(n_32), .Y(n_292) );
BUFx2_ASAP7_75t_L g344 ( .A(n_32), .Y(n_344) );
BUFx2_ASAP7_75t_L g366 ( .A(n_32), .Y(n_366) );
OR2x2_ASAP7_75t_L g603 ( .A(n_32), .B(n_384), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_33), .A2(n_95), .B1(n_868), .B2(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_33), .A2(n_95), .B1(n_923), .B2(n_924), .Y(n_922) );
INVx1_ASAP7_75t_L g839 ( .A(n_34), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_34), .A2(n_182), .B1(n_849), .B2(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g475 ( .A(n_35), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_35), .A2(n_144), .B1(n_363), .B2(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g1229 ( .A(n_36), .Y(n_1229) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_37), .A2(n_61), .B1(n_597), .B2(n_607), .C(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_37), .A2(n_61), .B1(n_657), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_38), .A2(n_100), .B1(n_776), .B2(n_778), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_38), .A2(n_100), .B1(n_485), .B2(n_486), .C(n_588), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g1053 ( .A1(n_39), .A2(n_44), .B1(n_390), .B2(n_431), .Y(n_1053) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_39), .A2(n_44), .B1(n_358), .B2(n_783), .C(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1295 ( .A(n_40), .Y(n_1295) );
CKINVDCx5p33_ASAP7_75t_R g1152 ( .A(n_41), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_42), .A2(n_208), .B1(n_776), .B2(n_783), .Y(n_842) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_42), .A2(n_208), .B1(n_853), .B2(n_859), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_43), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g1124 ( .A(n_45), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_46), .A2(n_50), .B1(n_313), .B2(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g797 ( .A(n_46), .Y(n_797) );
INVx1_ASAP7_75t_L g964 ( .A(n_47), .Y(n_964) );
INVx1_ASAP7_75t_L g905 ( .A(n_48), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_48), .A2(n_228), .B1(n_915), .B2(n_917), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_49), .Y(n_1031) );
INVx1_ASAP7_75t_L g796 ( .A(n_50), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g988 ( .A(n_51), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_52), .A2(n_245), .B1(n_912), .B2(n_913), .Y(n_1101) );
AOI22xp33_ASAP7_75t_SL g1108 ( .A1(n_52), .A2(n_245), .B1(n_664), .B2(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1076 ( .A(n_53), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_53), .A2(n_148), .B1(n_915), .B2(n_917), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_54), .A2(n_210), .B1(n_832), .B2(n_833), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_54), .A2(n_210), .B1(n_874), .B2(n_876), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g1425 ( .A1(n_55), .A2(n_73), .B1(n_485), .B2(n_486), .C(n_854), .Y(n_1425) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_55), .A2(n_73), .B1(n_352), .B2(n_1432), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_56), .A2(n_97), .B1(n_1180), .B2(n_1188), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_57), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_58), .Y(n_1033) );
INVx1_ASAP7_75t_L g720 ( .A(n_59), .Y(n_720) );
INVx1_ASAP7_75t_L g302 ( .A(n_60), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_60), .A2(n_62), .B1(n_413), .B2(n_415), .C(n_418), .Y(n_412) );
INVx1_ASAP7_75t_L g293 ( .A(n_62), .Y(n_293) );
INVx1_ASAP7_75t_L g1081 ( .A(n_63), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_63), .A2(n_115), .B1(n_1104), .B2(n_1106), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g1039 ( .A(n_64), .Y(n_1039) );
AO22x2_ASAP7_75t_L g892 ( .A1(n_65), .A2(n_893), .B1(n_945), .B2(n_946), .Y(n_892) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_65), .Y(n_945) );
AO221x1_ASAP7_75t_L g804 ( .A1(n_67), .A2(n_81), .B1(n_508), .B2(n_509), .C(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g820 ( .A(n_67), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_68), .A2(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g518 ( .A(n_68), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_69), .A2(n_234), .B1(n_649), .B2(n_1486), .Y(n_1489) );
INVx1_ASAP7_75t_L g1495 ( .A(n_69), .Y(n_1495) );
INVx1_ASAP7_75t_L g1117 ( .A(n_70), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1244 ( .A1(n_71), .A2(n_147), .B1(n_1180), .B2(n_1188), .Y(n_1244) );
INVx1_ASAP7_75t_L g1468 ( .A(n_72), .Y(n_1468) );
AOI22xp33_ASAP7_75t_L g1480 ( .A1(n_72), .A2(n_247), .B1(n_1018), .B2(n_1412), .Y(n_1480) );
INVx1_ASAP7_75t_L g902 ( .A(n_74), .Y(n_902) );
INVx1_ASAP7_75t_L g1137 ( .A(n_76), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_76), .A2(n_92), .B1(n_672), .B2(n_927), .Y(n_1170) );
INVxp33_ASAP7_75t_L g699 ( .A(n_77), .Y(n_699) );
XNOR2x2_ASAP7_75t_L g1071 ( .A(n_78), .B(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_79), .A2(n_162), .B1(n_362), .B2(n_364), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_79), .A2(n_162), .B1(n_456), .B2(n_461), .Y(n_455) );
INVxp33_ASAP7_75t_L g705 ( .A(n_80), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_80), .A2(n_126), .B1(n_555), .B2(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g822 ( .A(n_81), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g1414 ( .A1(n_82), .A2(n_99), .B1(n_418), .B2(n_935), .C(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1437 ( .A(n_82), .Y(n_1437) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_83), .Y(n_998) );
INVx1_ASAP7_75t_L g291 ( .A(n_84), .Y(n_291) );
INVx1_ASAP7_75t_L g342 ( .A(n_84), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_85), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_86), .A2(n_157), .B1(n_783), .B2(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g886 ( .A(n_86), .Y(n_886) );
AOI22xp33_ASAP7_75t_SL g843 ( .A1(n_87), .A2(n_137), .B1(n_347), .B2(n_362), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_87), .A2(n_137), .B1(n_500), .B2(n_857), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_89), .A2(n_121), .B1(n_1180), .B2(n_1188), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_90), .A2(n_191), .B1(n_1180), .B2(n_1188), .Y(n_1179) );
INVx1_ASAP7_75t_L g1473 ( .A(n_91), .Y(n_1473) );
OAI22xp33_ASAP7_75t_L g1497 ( .A1(n_91), .A2(n_181), .B1(n_938), .B2(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1144 ( .A(n_92), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_93), .A2(n_223), .B1(n_500), .B2(n_501), .C(n_504), .Y(n_499) );
INVx1_ASAP7_75t_L g523 ( .A(n_93), .Y(n_523) );
AOI22x1_ASAP7_75t_L g766 ( .A1(n_94), .A2(n_767), .B1(n_768), .B2(n_823), .Y(n_766) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_94), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_94), .A2(n_141), .B1(n_1192), .B2(n_1196), .Y(n_1199) );
CKINVDCx5p33_ASAP7_75t_R g995 ( .A(n_96), .Y(n_995) );
INVx1_ASAP7_75t_L g1213 ( .A(n_98), .Y(n_1213) );
INVx1_ASAP7_75t_L g1439 ( .A(n_99), .Y(n_1439) );
INVx1_ASAP7_75t_L g1140 ( .A(n_101), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_101), .A2(n_213), .B1(n_644), .B2(n_734), .C(n_1168), .Y(n_1167) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_102), .Y(n_628) );
INVx1_ASAP7_75t_L g1421 ( .A(n_103), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_103), .A2(n_221), .B1(n_644), .B2(n_928), .Y(n_1434) );
INVx1_ASAP7_75t_L g586 ( .A(n_104), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_104), .A2(n_205), .B1(n_647), .B2(n_648), .C(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g726 ( .A(n_105), .Y(n_726) );
INVx1_ASAP7_75t_L g829 ( .A(n_106), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_106), .A2(n_180), .B1(n_853), .B2(n_854), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g970 ( .A(n_107), .B(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g1019 ( .A(n_107), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_108), .A2(n_203), .B1(n_1412), .B2(n_1427), .Y(n_1426) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_108), .A2(n_203), .B1(n_644), .B2(n_655), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1476 ( .A1(n_109), .A2(n_218), .B1(n_503), .B2(n_800), .Y(n_1476) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_109), .A2(n_218), .B1(n_313), .B2(n_673), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_110), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_111), .A2(n_175), .B1(n_780), .B2(n_783), .Y(n_779) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_111), .A2(n_390), .B1(n_804), .B2(n_806), .C(n_810), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_112), .A2(n_197), .B1(n_364), .B2(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_112), .A2(n_197), .B1(n_503), .B2(n_800), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_113), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_114), .A2(n_225), .B1(n_912), .B2(n_913), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_114), .A2(n_225), .B1(n_653), .B2(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1075 ( .A(n_115), .Y(n_1075) );
INVx1_ASAP7_75t_L g255 ( .A(n_116), .Y(n_255) );
OA22x2_ASAP7_75t_L g952 ( .A1(n_117), .A2(n_953), .B1(n_1024), .B2(n_1025), .Y(n_952) );
INVxp67_ASAP7_75t_SL g1025 ( .A(n_117), .Y(n_1025) );
AO22x1_ASAP7_75t_SL g1209 ( .A1(n_118), .A2(n_198), .B1(n_1180), .B2(n_1188), .Y(n_1209) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_119), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_120), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_122), .Y(n_896) );
AOI21xp33_ASAP7_75t_L g484 ( .A1(n_123), .A2(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g553 ( .A(n_123), .Y(n_553) );
XOR2xp5_ASAP7_75t_L g577 ( .A(n_124), .B(n_578), .Y(n_577) );
AO221x2_ASAP7_75t_L g1223 ( .A1(n_124), .A2(n_237), .B1(n_1212), .B2(n_1224), .C(n_1225), .Y(n_1223) );
INVx1_ASAP7_75t_L g1293 ( .A(n_125), .Y(n_1293) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_126), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_127), .Y(n_1151) );
XNOR2xp5_ASAP7_75t_L g276 ( .A(n_128), .B(n_277), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_129), .A2(n_204), .B1(n_1412), .B2(n_1413), .Y(n_1411) );
INVx1_ASAP7_75t_L g1440 ( .A(n_129), .Y(n_1440) );
INVx1_ASAP7_75t_L g1424 ( .A(n_130), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_130), .A2(n_238), .B1(n_304), .B2(n_371), .Y(n_1433) );
INVx1_ASAP7_75t_L g615 ( .A(n_131), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_131), .A2(n_167), .B1(n_664), .B2(n_666), .C(n_668), .Y(n_663) );
INVx1_ASAP7_75t_L g624 ( .A(n_132), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_132), .A2(n_158), .B1(n_672), .B2(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g1089 ( .A(n_133), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_133), .A2(n_187), .B1(n_672), .B2(n_1112), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_134), .A2(n_229), .B1(n_672), .B2(n_924), .Y(n_929) );
INVx1_ASAP7_75t_L g943 ( .A(n_134), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_135), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_138), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_138), .A2(n_320), .B1(n_333), .B2(n_370), .C(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g593 ( .A(n_139), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_139), .A2(n_244), .B1(n_653), .B2(n_654), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g1146 ( .A(n_140), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_142), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_143), .A2(n_201), .B1(n_428), .B2(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1443 ( .A(n_143), .Y(n_1443) );
INVx1_ASAP7_75t_L g476 ( .A(n_144), .Y(n_476) );
INVx1_ASAP7_75t_L g1467 ( .A(n_145), .Y(n_1467) );
INVx1_ASAP7_75t_L g1122 ( .A(n_146), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_146), .A2(n_233), .B1(n_665), .B2(n_928), .Y(n_1163) );
INVx1_ASAP7_75t_L g1079 ( .A(n_148), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g1191 ( .A1(n_149), .A2(n_232), .B1(n_1192), .B2(n_1196), .Y(n_1191) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_150), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_151), .A2(n_215), .B1(n_364), .B2(n_774), .Y(n_864) );
INVx1_ASAP7_75t_L g880 ( .A(n_151), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_152), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_153), .A2(n_173), .B1(n_868), .B2(n_910), .Y(n_1100) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_153), .A2(n_173), .B1(n_923), .B2(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g450 ( .A(n_154), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_155), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_156), .A2(n_196), .B1(n_352), .B2(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g439 ( .A(n_156), .Y(n_439) );
INVx1_ASAP7_75t_L g867 ( .A(n_157), .Y(n_867) );
INVx1_ASAP7_75t_L g612 ( .A(n_158), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g1148 ( .A(n_159), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_160), .A2(n_227), .B1(n_854), .B2(n_1478), .Y(n_1477) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_160), .A2(n_227), .B1(n_649), .B2(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1061 ( .A(n_161), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_163), .Y(n_311) );
INVx1_ASAP7_75t_L g724 ( .A(n_164), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_165), .A2(n_220), .B1(n_1196), .B2(n_1212), .Y(n_1245) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_166), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_166), .B(n_255), .Y(n_1187) );
AND3x2_ASAP7_75t_L g1193 ( .A(n_166), .B(n_255), .C(n_1184), .Y(n_1193) );
INVx1_ASAP7_75t_L g618 ( .A(n_167), .Y(n_618) );
INVx1_ASAP7_75t_L g480 ( .A(n_168), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_169), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_170), .Y(n_505) );
INVx2_ASAP7_75t_L g268 ( .A(n_171), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_172), .Y(n_495) );
XOR2xp5_ASAP7_75t_L g690 ( .A(n_174), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g802 ( .A(n_175), .Y(n_802) );
INVx1_ASAP7_75t_L g1215 ( .A(n_176), .Y(n_1215) );
INVx1_ASAP7_75t_L g1184 ( .A(n_177), .Y(n_1184) );
INVx1_ASAP7_75t_L g1082 ( .A(n_178), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_178), .A2(n_200), .B1(n_876), .B2(n_937), .Y(n_1090) );
INVx1_ASAP7_75t_L g374 ( .A(n_179), .Y(n_374) );
INVx1_ASAP7_75t_L g835 ( .A(n_180), .Y(n_835) );
INVx1_ASAP7_75t_L g1472 ( .A(n_181), .Y(n_1472) );
INVx1_ASAP7_75t_L g838 ( .A(n_182), .Y(n_838) );
INVx1_ASAP7_75t_L g1094 ( .A(n_183), .Y(n_1094) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_184), .A2(n_188), .B1(n_597), .B2(n_604), .C(n_1130), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g1157 ( .A1(n_184), .A2(n_188), .B1(n_660), .B2(n_1158), .C(n_1160), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g1226 ( .A(n_185), .Y(n_1226) );
INVx1_ASAP7_75t_L g270 ( .A(n_186), .Y(n_270) );
INVx2_ASAP7_75t_L g395 ( .A(n_186), .Y(n_395) );
INVx1_ASAP7_75t_L g1096 ( .A(n_187), .Y(n_1096) );
AO22x2_ASAP7_75t_L g466 ( .A1(n_189), .A2(n_467), .B1(n_571), .B2(n_572), .Y(n_466) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_189), .Y(n_571) );
INVx1_ASAP7_75t_L g1035 ( .A(n_190), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_190), .A2(n_216), .B1(n_783), .B2(n_1056), .C(n_1058), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1449 ( .A1(n_191), .A2(n_1450), .B1(n_1455), .B2(n_1504), .Y(n_1449) );
XNOR2xp5_ASAP7_75t_L g1459 ( .A(n_191), .B(n_1460), .Y(n_1459) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_192), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g1289 ( .A1(n_193), .A2(n_194), .B1(n_1290), .B2(n_1291), .C(n_1292), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1407 ( .A(n_195), .B(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g443 ( .A(n_196), .Y(n_443) );
INVx1_ASAP7_75t_L g729 ( .A(n_199), .Y(n_729) );
INVx1_ASAP7_75t_L g1084 ( .A(n_200), .Y(n_1084) );
INVx1_ASAP7_75t_L g1442 ( .A(n_201), .Y(n_1442) );
INVx1_ASAP7_75t_L g904 ( .A(n_202), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_202), .A2(n_209), .B1(n_868), .B2(n_910), .Y(n_918) );
INVx1_ASAP7_75t_L g1436 ( .A(n_204), .Y(n_1436) );
INVx1_ASAP7_75t_L g590 ( .A(n_205), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_206), .Y(n_1042) );
INVx1_ASAP7_75t_L g1005 ( .A(n_207), .Y(n_1005) );
INVx1_ASAP7_75t_L g899 ( .A(n_209), .Y(n_899) );
OAI211xp5_ASAP7_75t_L g976 ( .A1(n_211), .A2(n_977), .B(n_979), .C(n_983), .Y(n_976) );
INVx1_ASAP7_75t_L g1022 ( .A(n_211), .Y(n_1022) );
INVx1_ASAP7_75t_L g1048 ( .A(n_212), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_212), .Y(n_1064) );
INVx1_ASAP7_75t_L g1138 ( .A(n_213), .Y(n_1138) );
INVxp33_ASAP7_75t_SL g700 ( .A(n_214), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_214), .A2(n_222), .B1(n_740), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g883 ( .A(n_215), .Y(n_883) );
AOI21xp33_ASAP7_75t_L g1037 ( .A1(n_216), .A2(n_385), .B(n_486), .Y(n_1037) );
INVx1_ASAP7_75t_L g1185 ( .A(n_217), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_217), .B(n_1183), .Y(n_1190) );
INVx1_ASAP7_75t_L g941 ( .A(n_219), .Y(n_941) );
INVx1_ASAP7_75t_L g1422 ( .A(n_221), .Y(n_1422) );
INVxp33_ASAP7_75t_SL g695 ( .A(n_222), .Y(n_695) );
INVx1_ASAP7_75t_L g531 ( .A(n_223), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_224), .Y(n_282) );
OAI211xp5_ASAP7_75t_L g960 ( .A1(n_226), .A2(n_434), .B(n_961), .C(n_962), .Y(n_960) );
INVx1_ASAP7_75t_L g1002 ( .A(n_226), .Y(n_1002) );
INVx1_ASAP7_75t_L g897 ( .A(n_228), .Y(n_897) );
INVx1_ASAP7_75t_L g934 ( .A(n_229), .Y(n_934) );
INVx1_ASAP7_75t_L g1126 ( .A(n_230), .Y(n_1126) );
AOI21xp33_ASAP7_75t_L g1164 ( .A1(n_230), .A2(n_782), .B(n_1165), .Y(n_1164) );
INVx2_ASAP7_75t_L g267 ( .A(n_231), .Y(n_267) );
INVx1_ASAP7_75t_L g1127 ( .A(n_233), .Y(n_1127) );
INVx1_ASAP7_75t_L g1503 ( .A(n_234), .Y(n_1503) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_235), .A2(n_236), .B1(n_353), .B2(n_358), .Y(n_357) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_235), .A2(n_390), .B(n_400), .C(n_423), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_236), .A2(n_431), .B1(n_433), .B2(n_447), .C(n_453), .Y(n_430) );
INVx1_ASAP7_75t_L g1416 ( .A(n_238), .Y(n_1416) );
INVxp33_ASAP7_75t_SL g709 ( .A(n_239), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_240), .Y(n_1154) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_241), .Y(n_991) );
INVx1_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
BUFx3_ASAP7_75t_L g308 ( .A(n_242), .Y(n_308) );
BUFx3_ASAP7_75t_L g287 ( .A(n_243), .Y(n_287) );
INVx1_ASAP7_75t_L g300 ( .A(n_243), .Y(n_300) );
INVx1_ASAP7_75t_L g582 ( .A(n_244), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_246), .Y(n_473) );
INVx1_ASAP7_75t_L g1464 ( .A(n_247), .Y(n_1464) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_248), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_271), .B(n_1172), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_258), .Y(n_252) );
AND2x4_ASAP7_75t_L g1454 ( .A(n_253), .B(n_259), .Y(n_1454) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_SL g1448 ( .A(n_254), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_254), .B(n_256), .Y(n_1506) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_256), .B(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g889 ( .A(n_261), .B(n_366), .Y(n_889) );
OR2x2_ASAP7_75t_L g944 ( .A(n_261), .B(n_366), .Y(n_944) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g446 ( .A(n_262), .B(n_270), .Y(n_446) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g486 ( .A(n_263), .B(n_487), .Y(n_486) );
INVx8_ASAP7_75t_L g885 ( .A(n_264), .Y(n_885) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_265), .Y(n_442) );
INVx1_ASAP7_75t_L g614 ( .A(n_265), .Y(n_614) );
OR2x2_ASAP7_75t_L g688 ( .A(n_265), .B(n_603), .Y(n_688) );
INVx2_ASAP7_75t_SL g708 ( .A(n_265), .Y(n_708) );
OR2x6_ASAP7_75t_L g888 ( .A(n_265), .B(n_879), .Y(n_888) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_265), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g387 ( .A(n_267), .B(n_268), .Y(n_387) );
INVx1_ASAP7_75t_L g398 ( .A(n_267), .Y(n_398) );
INVx2_ASAP7_75t_L g405 ( .A(n_267), .Y(n_405) );
AND2x4_ASAP7_75t_L g411 ( .A(n_267), .B(n_399), .Y(n_411) );
INVx1_ASAP7_75t_L g438 ( .A(n_267), .Y(n_438) );
INVx2_ASAP7_75t_L g399 ( .A(n_268), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_268), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g426 ( .A(n_268), .Y(n_426) );
INVx1_ASAP7_75t_L g437 ( .A(n_268), .Y(n_437) );
INVx1_ASAP7_75t_L g460 ( .A(n_268), .Y(n_460) );
AND2x4_ASAP7_75t_L g875 ( .A(n_269), .B(n_426), .Y(n_875) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g876 ( .A(n_270), .B(n_815), .Y(n_876) );
OR2x2_ASAP7_75t_L g938 ( .A(n_270), .B(n_815), .Y(n_938) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_948), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_759), .B1(n_760), .B2(n_947), .Y(n_272) );
INVx2_ASAP7_75t_L g947 ( .A(n_273), .Y(n_947) );
AOI22x1_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_575), .B1(n_757), .B2(n_758), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g757 ( .A(n_275), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_466), .B1(n_573), .B2(n_574), .Y(n_275) );
INVx1_ASAP7_75t_L g573 ( .A(n_276), .Y(n_573) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_373), .C(n_388), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_316), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_301), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_293), .B2(n_294), .Y(n_281) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_282), .A2(n_311), .B1(n_401), .B2(n_406), .C(n_412), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g819 ( .A1(n_283), .A2(n_303), .B1(n_376), .B2(n_807), .C1(n_811), .C2(n_820), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_283), .A2(n_294), .B1(n_1040), .B2(n_1042), .Y(n_1067) );
AOI22xp5_ASAP7_75t_L g1435 ( .A1(n_283), .A2(n_294), .B1(n_1436), .B2(n_1437), .Y(n_1435) );
CKINVDCx6p67_ASAP7_75t_R g283 ( .A(n_284), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_285), .B(n_289), .Y(n_284) );
INVx2_ASAP7_75t_L g655 ( .A(n_285), .Y(n_655) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g350 ( .A(n_286), .Y(n_350) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_286), .Y(n_533) );
INVx1_ASAP7_75t_L g556 ( .A(n_286), .Y(n_556) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_286), .Y(n_928) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
AND2x2_ASAP7_75t_L g356 ( .A(n_287), .B(n_308), .Y(n_356) );
INVx1_ASAP7_75t_L g298 ( .A(n_288), .Y(n_298) );
OR2x6_ASAP7_75t_L g295 ( .A(n_289), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g310 ( .A(n_289), .Y(n_310) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx2_ASAP7_75t_L g645 ( .A(n_290), .Y(n_645) );
OR2x2_ASAP7_75t_L g682 ( .A(n_290), .B(n_552), .Y(n_682) );
OR2x2_ASAP7_75t_L g684 ( .A(n_290), .B(n_350), .Y(n_684) );
INVx1_ASAP7_75t_L g327 ( .A(n_291), .Y(n_327) );
INVx1_ASAP7_75t_L g330 ( .A(n_292), .Y(n_330) );
AND2x4_ASAP7_75t_L g585 ( .A(n_292), .B(n_394), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_294), .A2(n_312), .B1(n_809), .B2(n_822), .Y(n_821) );
CKINVDCx6p67_ASAP7_75t_R g294 ( .A(n_295), .Y(n_294) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_296), .Y(n_1001) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g565 ( .A(n_297), .Y(n_565) );
BUFx4f_ASAP7_75t_L g1162 ( .A(n_297), .Y(n_1162) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g552 ( .A(n_298), .B(n_299), .Y(n_552) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g315 ( .A(n_300), .B(n_308), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_311), .B2(n_312), .Y(n_301) );
AOI222xp33_ASAP7_75t_L g1065 ( .A1(n_303), .A2(n_312), .B1(n_376), .B2(n_1039), .C1(n_1045), .C2(n_1066), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_303), .A2(n_312), .B1(n_1439), .B2(n_1440), .Y(n_1438) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_310), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g672 ( .A(n_305), .Y(n_672) );
INVx1_ASAP7_75t_L g1486 ( .A(n_305), .Y(n_1486) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
INVx6_ASAP7_75t_L g360 ( .A(n_306), .Y(n_360) );
AND2x2_ASAP7_75t_L g377 ( .A(n_306), .B(n_326), .Y(n_377) );
AND2x4_ASAP7_75t_L g528 ( .A(n_306), .B(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
AND2x2_ASAP7_75t_L g312 ( .A(n_310), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g774 ( .A(n_314), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_314), .A2(n_1004), .B1(n_1005), .B2(n_1006), .Y(n_1003) );
INVx2_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_315), .Y(n_363) );
AND2x6_ASAP7_75t_L g524 ( .A(n_315), .B(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_315), .Y(n_560) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_315), .Y(n_644) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_315), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_337), .C(n_368), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_331), .B2(n_332), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_318), .A2(n_331), .B1(n_424), .B2(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g788 ( .A(n_320), .Y(n_788) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g659 ( .A(n_322), .Y(n_659) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g540 ( .A(n_323), .Y(n_540) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
OR2x6_ASAP7_75t_L g333 ( .A(n_325), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_326), .B(n_330), .Y(n_325) );
AND2x4_ASAP7_75t_L g658 ( .A(n_326), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_326), .B(n_335), .Y(n_661) );
INVx1_ASAP7_75t_L g678 ( .A(n_326), .Y(n_678) );
AND2x4_ASAP7_75t_L g1159 ( .A(n_326), .B(n_659), .Y(n_1159) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x4_ASAP7_75t_L g367 ( .A(n_328), .B(n_342), .Y(n_367) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g341 ( .A(n_329), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g521 ( .A(n_329), .Y(n_521) );
INVx1_ASAP7_75t_L g526 ( .A(n_329), .Y(n_526) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_329), .Y(n_530) );
OR2x6_ASAP7_75t_L g637 ( .A(n_330), .B(n_420), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_332), .A2(n_788), .B1(n_789), .B2(n_790), .C(n_791), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g1441 ( .A1(n_332), .A2(n_788), .B1(n_791), .B2(n_1442), .C(n_1443), .Y(n_1441) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g744 ( .A(n_334), .B(n_678), .Y(n_744) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x6_ASAP7_75t_L g541 ( .A(n_336), .B(n_526), .Y(n_541) );
AOI33xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_345), .A3(n_351), .B1(n_357), .B2(n_361), .B3(n_365), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g1054 ( .A1(n_338), .A2(n_570), .B1(n_1055), .B2(n_1059), .C(n_1063), .Y(n_1054) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_339), .A2(n_548), .B1(n_562), .B2(n_568), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_339), .Y(n_921) );
OR2x6_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
OR2x2_ASAP7_75t_L g772 ( .A(n_340), .B(n_343), .Y(n_772) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g670 ( .A(n_341), .Y(n_670) );
INVx1_ASAP7_75t_L g750 ( .A(n_341), .Y(n_750) );
INVx1_ASAP7_75t_L g846 ( .A(n_341), .Y(n_846) );
BUFx3_ASAP7_75t_L g1169 ( .A(n_341), .Y(n_1169) );
INVx1_ASAP7_75t_L g514 ( .A(n_342), .Y(n_514) );
INVx2_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
BUFx2_ASAP7_75t_L g465 ( .A(n_343), .Y(n_465) );
OR2x2_ASAP7_75t_L g845 ( .A(n_343), .B(n_846), .Y(n_845) );
AND2x4_ASAP7_75t_L g860 ( .A(n_343), .B(n_446), .Y(n_860) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_343), .B(n_419), .Y(n_1483) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g515 ( .A(n_344), .Y(n_515) );
OR2x6_ASAP7_75t_L g610 ( .A(n_344), .B(n_486), .Y(n_610) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g364 ( .A(n_348), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_348), .A2(n_559), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g742 ( .A(n_349), .Y(n_742) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g993 ( .A(n_350), .Y(n_993) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g1112 ( .A(n_354), .Y(n_1112) );
INVx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_355), .Y(n_371) );
INVx1_ASAP7_75t_L g536 ( .A(n_355), .Y(n_536) );
AND2x4_ASAP7_75t_L g675 ( .A(n_355), .B(n_645), .Y(n_675) );
BUFx4f_ASAP7_75t_L g778 ( .A(n_355), .Y(n_778) );
BUFx3_ASAP7_75t_L g1471 ( .A(n_355), .Y(n_1471) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_356), .Y(n_546) );
INVx4_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g647 ( .A(n_359), .Y(n_647) );
INVx2_ASAP7_75t_L g863 ( .A(n_359), .Y(n_863) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g522 ( .A(n_360), .Y(n_522) );
INVx2_ASAP7_75t_L g753 ( .A(n_360), .Y(n_753) );
INVx2_ASAP7_75t_L g777 ( .A(n_360), .Y(n_777) );
INVx2_ASAP7_75t_SL g782 ( .A(n_360), .Y(n_782) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_360), .Y(n_1057) );
BUFx4f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g931 ( .A(n_363), .Y(n_931) );
AOI33xp33_ASAP7_75t_L g770 ( .A1(n_365), .A2(n_771), .A3(n_773), .B1(n_775), .B2(n_779), .B3(n_785), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g861 ( .A(n_365), .B(n_862), .C(n_864), .Y(n_861) );
AOI33xp33_ASAP7_75t_L g1429 ( .A1(n_365), .A2(n_844), .A3(n_1430), .B1(n_1431), .B2(n_1433), .B3(n_1434), .Y(n_1429) );
NAND3xp33_ASAP7_75t_L g1488 ( .A(n_365), .B(n_1489), .C(n_1490), .Y(n_1488) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x4_ASAP7_75t_L g376 ( .A(n_366), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g570 ( .A(n_366), .B(n_367), .Y(n_570) );
INVx2_ASAP7_75t_L g651 ( .A(n_367), .Y(n_651) );
INVx2_ASAP7_75t_SL g738 ( .A(n_367), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g1165 ( .A(n_367), .Y(n_1165) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_371), .Y(n_561) );
BUFx2_ASAP7_75t_SL g749 ( .A(n_371), .Y(n_749) );
AND2x2_ASAP7_75t_L g791 ( .A(n_372), .B(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g1408 ( .A(n_375), .Y(n_1408) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx2_ASAP7_75t_L g689 ( .A(n_376), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_L g640 ( .A(n_379), .Y(n_640) );
INVx1_ASAP7_75t_L g471 ( .A(n_380), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_385), .Y(n_380) );
AND2x2_ASAP7_75t_L g424 ( .A(n_381), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x6_ASAP7_75t_L g428 ( .A(n_382), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g453 ( .A(n_382), .B(n_454), .Y(n_453) );
OR2x6_ASAP7_75t_L g511 ( .A(n_382), .B(n_454), .Y(n_511) );
INVx1_ASAP7_75t_L g816 ( .A(n_382), .Y(n_816) );
INVx1_ASAP7_75t_L g1419 ( .A(n_382), .Y(n_1419) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g853 ( .A(n_385), .Y(n_853) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g508 ( .A(n_386), .Y(n_508) );
INVx2_ASAP7_75t_SL g592 ( .A(n_386), .Y(n_592) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
OAI31xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_430), .A3(n_455), .B(n_463), .Y(n_388) );
INVx8_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_391), .A2(n_432), .B1(n_470), .B2(n_471), .C1(n_472), .C2(n_473), .Y(n_469) );
AOI221xp5_ASAP7_75t_SL g1410 ( .A1(n_391), .A2(n_1411), .B1(n_1414), .B2(n_1416), .C(n_1417), .Y(n_1410) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
AND2x4_ASAP7_75t_L g462 ( .A(n_392), .B(n_409), .Y(n_462) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g432 ( .A(n_394), .B(n_417), .Y(n_432) );
AND2x2_ASAP7_75t_L g457 ( .A(n_394), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
INVx1_ASAP7_75t_L g487 ( .A(n_395), .Y(n_487) );
INVx1_ASAP7_75t_L g414 ( .A(n_396), .Y(n_414) );
BUFx6f_ASAP7_75t_L g1482 ( .A(n_396), .Y(n_1482) );
BUFx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g588 ( .A(n_397), .Y(n_588) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_397), .Y(n_805) );
BUFx6f_ASAP7_75t_L g854 ( .A(n_397), .Y(n_854) );
AND2x4_ASAP7_75t_L g870 ( .A(n_397), .B(n_871), .Y(n_870) );
AND2x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g490 ( .A(n_404), .Y(n_490) );
INVx1_ASAP7_75t_L g623 ( .A(n_404), .Y(n_623) );
INVx1_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
AND2x4_ASAP7_75t_L g458 ( .A(n_405), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g857 ( .A(n_408), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_408), .A2(n_988), .B1(n_991), .B2(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g1427 ( .A(n_410), .Y(n_1427) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g452 ( .A(n_411), .Y(n_452) );
INVx3_ASAP7_75t_L g494 ( .A(n_411), .Y(n_494) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_411), .Y(n_503) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g935 ( .A(n_414), .Y(n_935) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_415), .A2(n_811), .B(n_812), .C(n_816), .Y(n_810) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g963 ( .A(n_416), .Y(n_963) );
INVx2_ASAP7_75t_SL g1478 ( .A(n_416), .Y(n_1478) );
INVx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_417), .Y(n_485) );
BUFx2_ASAP7_75t_L g1415 ( .A(n_417), .Y(n_1415) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g509 ( .A(n_420), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g872 ( .A(n_421), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_424), .A2(n_427), .B1(n_497), .B2(n_498), .Y(n_496) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g601 ( .A(n_426), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g1047 ( .A1(n_426), .A2(n_606), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
CKINVDCx11_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g606 ( .A(n_429), .Y(n_606) );
CKINVDCx6p67_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_432), .A2(n_799), .B1(n_801), .B2(n_802), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g1423 ( .A1(n_432), .A2(n_510), .B1(n_1424), .B2(n_1425), .C(n_1426), .Y(n_1423) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_439), .B1(n_440), .B2(n_443), .C(n_444), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g1134 ( .A1(n_434), .A2(n_1135), .B1(n_1137), .B2(n_1138), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g1149 ( .A1(n_434), .A2(n_1150), .B1(n_1151), .B2(n_1152), .Y(n_1149) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g454 ( .A(n_436), .Y(n_454) );
INVx2_ASAP7_75t_L g506 ( .A(n_436), .Y(n_506) );
INVx3_ASAP7_75t_L g1036 ( .A(n_436), .Y(n_1036) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_437), .B(n_438), .Y(n_483) );
INVx1_ASAP7_75t_L g815 ( .A(n_438), .Y(n_815) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g1009 ( .A1(n_442), .A2(n_995), .B1(n_998), .B2(n_1010), .Y(n_1009) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_442), .A2(n_727), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_442), .Y(n_1150) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_449), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_449), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_449), .A2(n_808), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g626 ( .A(n_451), .Y(n_626) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g882 ( .A(n_452), .Y(n_882) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_454), .Y(n_710) );
INVx1_ASAP7_75t_L g1011 ( .A(n_454), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_454), .B(n_1047), .Y(n_1046) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_457), .A2(n_462), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_457), .A2(n_462), .B1(n_796), .B2(n_797), .Y(n_795) );
INVx3_ASAP7_75t_L g1051 ( .A(n_457), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_457), .A2(n_462), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
BUFx2_ASAP7_75t_L g500 ( .A(n_458), .Y(n_500) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_458), .Y(n_595) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_458), .Y(n_800) );
INVx1_ASAP7_75t_L g850 ( .A(n_458), .Y(n_850) );
AND2x4_ASAP7_75t_L g878 ( .A(n_458), .B(n_879), .Y(n_878) );
BUFx2_ASAP7_75t_L g912 ( .A(n_458), .Y(n_912) );
BUFx6f_ASAP7_75t_L g1412 ( .A(n_458), .Y(n_1412) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g1052 ( .A(n_462), .Y(n_1052) );
AOI31xp33_ASAP7_75t_L g1155 ( .A1(n_463), .A2(n_1156), .A3(n_1166), .B(n_1171), .Y(n_1155) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
CKINVDCx8_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
AOI221x1_ASAP7_75t_SL g467 ( .A1(n_465), .A2(n_468), .B1(n_512), .B2(n_516), .C(n_547), .Y(n_467) );
INVx2_ASAP7_75t_SL g574 ( .A(n_466), .Y(n_574) );
INVx1_ASAP7_75t_L g572 ( .A(n_467), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_474), .C(n_477), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_470), .A2(n_528), .B1(n_531), .B2(n_532), .Y(n_527) );
OAI221xp5_ASAP7_75t_L g562 ( .A1(n_472), .A2(n_473), .B1(n_550), .B2(n_563), .C(n_566), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_499), .C(n_510), .Y(n_477) );
OAI21xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_488), .B(n_496), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_484), .Y(n_479) );
BUFx3_ASAP7_75t_L g616 ( .A(n_481), .Y(n_616) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g728 ( .A(n_482), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_482), .B(n_813), .Y(n_812) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g1044 ( .A1(n_485), .A2(n_816), .B(n_1045), .C(n_1046), .Y(n_1044) );
INVx1_ASAP7_75t_L g1105 ( .A(n_485), .Y(n_1105) );
INVx1_ASAP7_75t_L g879 ( .A(n_487), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_491), .B1(n_492), .B2(n_495), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_489), .A2(n_720), .B1(n_721), .B2(n_724), .Y(n_719) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g957 ( .A(n_490), .B(n_958), .Y(n_957) );
INVx2_ASAP7_75t_L g1014 ( .A(n_490), .Y(n_1014) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g584 ( .A(n_493), .B(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g718 ( .A(n_494), .Y(n_718) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_494), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_495), .A2(n_549), .B1(n_553), .B2(n_554), .C(n_557), .Y(n_548) );
AOI222xp33_ASAP7_75t_L g534 ( .A1(n_497), .A2(n_498), .B1(n_505), .B2(n_535), .C1(n_537), .C2(n_541), .Y(n_534) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_SL g913 ( .A(n_502), .Y(n_913) );
INVx4_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_SL g629 ( .A(n_503), .Y(n_629) );
BUFx3_ASAP7_75t_L g917 ( .A(n_503), .Y(n_917) );
OAI21xp5_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_506), .B(n_507), .Y(n_504) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_506), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g1041 ( .A1(n_506), .A2(n_1042), .B(n_1043), .Y(n_1041) );
BUFx3_ASAP7_75t_L g910 ( .A(n_508), .Y(n_910) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AOI211x1_ASAP7_75t_L g1072 ( .A1(n_512), .A2(n_1073), .B(n_1085), .C(n_1098), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AO211x2_ASAP7_75t_L g826 ( .A1(n_513), .A2(n_827), .B(n_840), .C(n_865), .Y(n_826) );
AOI211x1_ASAP7_75t_SL g893 ( .A1(n_513), .A2(n_894), .B(n_906), .C(n_932), .Y(n_893) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
AND2x4_ASAP7_75t_L g984 ( .A(n_514), .B(n_515), .Y(n_984) );
INVx2_ASAP7_75t_L g818 ( .A(n_515), .Y(n_818) );
NAND4xp25_ASAP7_75t_SL g516 ( .A(n_517), .B(n_527), .C(n_534), .D(n_542), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_523), .B2(n_524), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_519), .A2(n_528), .B1(n_835), .B2(n_836), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_519), .A2(n_524), .B1(n_904), .B2(n_905), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_519), .A2(n_524), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
AND2x6_ASAP7_75t_L g532 ( .A(n_520), .B(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g1466 ( .A(n_520), .B(n_522), .Y(n_1466) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_524), .A2(n_532), .B1(n_838), .B2(n_839), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1465 ( .A1(n_524), .A2(n_1466), .B1(n_1467), .B2(n_1468), .Y(n_1465) );
INVx1_ASAP7_75t_L g545 ( .A(n_525), .Y(n_545) );
INVx1_ASAP7_75t_L g974 ( .A(n_525), .Y(n_974) );
AND2x2_ASAP7_75t_L g978 ( .A(n_525), .B(n_649), .Y(n_978) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_528), .A2(n_532), .B1(n_896), .B2(n_897), .Y(n_895) );
INVx4_ASAP7_75t_L g975 ( .A(n_528), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_528), .A2(n_532), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1462 ( .A1(n_528), .A2(n_532), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
AND2x4_ASAP7_75t_L g538 ( .A(n_529), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_SL g982 ( .A(n_529), .B(n_539), .Y(n_982) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g971 ( .A(n_532), .Y(n_971) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_533), .Y(n_673) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_533), .Y(n_786) );
INVx1_ASAP7_75t_L g1006 ( .A(n_533), .Y(n_1006) );
INVx2_ASAP7_75t_L g1110 ( .A(n_533), .Y(n_1110) );
INVx1_ASAP7_75t_L g1492 ( .A(n_533), .Y(n_1492) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI222xp33_ASAP7_75t_L g898 ( .A1(n_537), .A2(n_541), .B1(n_899), .B2(n_900), .C1(n_901), .C2(n_902), .Y(n_898) );
BUFx4f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g832 ( .A(n_538), .Y(n_832) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g833 ( .A(n_541), .Y(n_833) );
AOI322xp5_ASAP7_75t_L g979 ( .A1(n_541), .A2(n_560), .A3(n_965), .B1(n_968), .B2(n_980), .C1(n_981), .C2(n_982), .Y(n_979) );
AOI222xp33_ASAP7_75t_L g1080 ( .A1(n_541), .A2(n_778), .B1(n_1081), .B2(n_1082), .C1(n_1083), .C2(n_1084), .Y(n_1080) );
AOI222xp33_ASAP7_75t_L g1469 ( .A1(n_541), .A2(n_982), .B1(n_1470), .B2(n_1471), .C1(n_1472), .C2(n_1473), .Y(n_1469) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND4xp25_ASAP7_75t_L g894 ( .A(n_543), .B(n_895), .C(n_898), .D(n_903), .Y(n_894) );
NAND4xp25_ASAP7_75t_SL g1073 ( .A(n_543), .B(n_1074), .C(n_1077), .D(n_1080), .Y(n_1073) );
NAND4xp25_ASAP7_75t_L g1461 ( .A(n_543), .B(n_1462), .C(n_1465), .D(n_1469), .Y(n_1461) );
INVx5_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI211xp5_ASAP7_75t_L g828 ( .A1(n_544), .A2(n_829), .B(n_830), .C(n_831), .Y(n_828) );
CKINVDCx8_ASAP7_75t_R g983 ( .A(n_544), .Y(n_983) );
AND2x4_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_546), .Y(n_649) );
INVx1_ASAP7_75t_L g667 ( .A(n_546), .Y(n_667) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_546), .Y(n_679) );
INVx2_ASAP7_75t_L g784 ( .A(n_546), .Y(n_784) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g973 ( .A(n_552), .B(n_974), .Y(n_973) );
INVx2_ASAP7_75t_L g997 ( .A(n_552), .Y(n_997) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g567 ( .A(n_556), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_556), .A2(n_748), .B1(n_1031), .B2(n_1033), .Y(n_1058) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g990 ( .A(n_559), .Y(n_990) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g999 ( .A(n_565), .Y(n_999) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
BUFx4f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI33xp33_ASAP7_75t_L g920 ( .A1(n_570), .A2(n_921), .A3(n_922), .B1(n_926), .B2(n_929), .B3(n_930), .Y(n_920) );
INVx4_ASAP7_75t_L g1007 ( .A(n_570), .Y(n_1007) );
BUFx4f_ASAP7_75t_L g1115 ( .A(n_570), .Y(n_1115) );
INVx1_ASAP7_75t_L g758 ( .A(n_575), .Y(n_758) );
AO22x2_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_690), .B2(n_756), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_638), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_596), .C(n_609), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_589), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_586), .B2(n_587), .Y(n_581) );
BUFx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g696 ( .A(n_584), .Y(n_696) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_584), .Y(n_1123) );
AND2x6_ASAP7_75t_L g587 ( .A(n_585), .B(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g591 ( .A(n_585), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g594 ( .A(n_585), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_585), .B(n_595), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_587), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_587), .A2(n_1122), .B1(n_1123), .B2(n_1124), .Y(n_1121) );
NAND2x1p5_ASAP7_75t_L g608 ( .A(n_588), .B(n_602), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_593), .B2(n_594), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_591), .A2(n_594), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_591), .A2(n_1126), .B1(n_1127), .B2(n_1128), .Y(n_1125) );
INVx2_ASAP7_75t_SL g916 ( .A(n_595), .Y(n_916) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2x1_ASAP7_75t_SL g599 ( .A(n_600), .B(n_602), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_600), .A2(n_789), .B1(n_790), .B2(n_814), .Y(n_813) );
NAND2x1p5_ASAP7_75t_L g1418 ( .A(n_600), .B(n_1419), .Y(n_1418) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g605 ( .A(n_602), .B(n_606), .Y(n_605) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx4f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx4f_ASAP7_75t_L g702 ( .A(n_605), .Y(n_702) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g1130 ( .A(n_608), .Y(n_1130) );
OAI33xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .A3(n_617), .B1(n_627), .B2(n_631), .B3(n_635), .Y(n_609) );
OAI33xp33_ASAP7_75t_L g703 ( .A1(n_610), .A2(n_635), .A3(n_704), .B1(n_711), .B2(n_719), .B3(n_725), .Y(n_703) );
OAI33xp33_ASAP7_75t_L g1008 ( .A1(n_610), .A2(n_1009), .A3(n_1012), .B1(n_1015), .B2(n_1020), .B3(n_1023), .Y(n_1008) );
INVx1_ASAP7_75t_L g1133 ( .A(n_610), .Y(n_1133) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_615), .B2(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g632 ( .A(n_614), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_624), .B2(n_625), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_619), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g713 ( .A(n_622), .Y(n_713) );
INVx2_ASAP7_75t_SL g1016 ( .A(n_622), .Y(n_1016) );
BUFx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g1143 ( .A(n_623), .Y(n_1143) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_628), .A2(n_643), .B1(n_646), .B2(n_652), .C(n_656), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_630), .A2(n_633), .B1(n_681), .B2(n_683), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_634), .A2(n_663), .B1(n_671), .B2(n_674), .C(n_676), .Y(n_662) );
OAI33xp33_ASAP7_75t_L g1131 ( .A1(n_635), .A2(n_1132), .A3(n_1134), .B1(n_1139), .B2(n_1145), .B3(n_1149), .Y(n_1131) );
CKINVDCx8_ASAP7_75t_R g635 ( .A(n_636), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g847 ( .A(n_636), .B(n_848), .C(n_852), .Y(n_847) );
INVx5_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx6_ASAP7_75t_L g919 ( .A(n_637), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B1(n_685), .B2(n_686), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_639), .A2(n_686), .B1(n_731), .B2(n_755), .Y(n_730) );
AOI31xp33_ASAP7_75t_L g1409 ( .A1(n_639), .A2(n_1410), .A3(n_1420), .B(n_1423), .Y(n_1409) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI31xp33_ASAP7_75t_L g1028 ( .A1(n_640), .A2(n_1029), .A3(n_1050), .B(n_1053), .Y(n_1028) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_662), .C(n_680), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_643), .A2(n_720), .B1(n_733), .B2(n_739), .C(n_743), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g1156 ( .A1(n_643), .A2(n_1146), .B(n_1157), .Y(n_1156) );
AND2x4_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
BUFx3_ASAP7_75t_L g653 ( .A(n_644), .Y(n_653) );
INVx1_ASAP7_75t_L g741 ( .A(n_644), .Y(n_741) );
INVx2_ASAP7_75t_SL g748 ( .A(n_644), .Y(n_748) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_649), .Y(n_830) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_649), .Y(n_900) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
BUFx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g792 ( .A(n_667), .Y(n_792) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_674), .A2(n_676), .B1(n_729), .B2(n_746), .C(n_751), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g1166 ( .A1(n_674), .A2(n_676), .B1(n_1152), .B2(n_1167), .C(n_1170), .Y(n_1166) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x4_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g735 ( .A(n_679), .Y(n_735) );
INVx1_ASAP7_75t_L g925 ( .A(n_679), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_681), .A2(n_683), .B1(n_724), .B2(n_726), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_681), .A2(n_683), .B1(n_1148), .B2(n_1151), .Y(n_1171) );
INVx6_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx4_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g1153 ( .A1(n_686), .A2(n_1154), .B(n_1155), .Y(n_1153) );
INVx5_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g756 ( .A(n_690), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_730), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_701), .C(n_703), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_698), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_709), .B2(n_710), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_706), .A2(n_726), .B1(n_727), .B2(n_729), .Y(n_725) );
BUFx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g808 ( .A(n_718), .Y(n_808) );
INVx2_ASAP7_75t_L g1032 ( .A(n_718), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1413 ( .A(n_718), .Y(n_1413) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g1018 ( .A(n_723), .Y(n_1018) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_745), .C(n_754), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
BUFx3_ASAP7_75t_L g923 ( .A(n_753), .Y(n_923) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
XNOR2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_891), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_824), .B2(n_890), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND4xp75_ASAP7_75t_L g768 ( .A(n_769), .B(n_793), .C(n_819), .D(n_821), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_787), .Y(n_769) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
OAI33xp33_ASAP7_75t_L g986 ( .A1(n_772), .A2(n_987), .A3(n_994), .B1(n_1000), .B2(n_1003), .B3(n_1007), .Y(n_986) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g1432 ( .A(n_784), .Y(n_1432) );
OAI21xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_803), .B(n_817), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_798), .Y(n_794) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_805), .Y(n_859) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_805), .Y(n_1088) );
INVx2_ASAP7_75t_L g851 ( .A(n_808), .Y(n_851) );
AND2x4_ASAP7_75t_L g966 ( .A(n_814), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx8_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g890 ( .A(n_824), .Y(n_890) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_834), .C(n_837), .Y(n_827) );
INVx1_ASAP7_75t_L g1083 ( .A(n_832), .Y(n_1083) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_836), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_884) );
NAND4xp25_ASAP7_75t_L g840 ( .A(n_841), .B(n_847), .C(n_855), .D(n_861), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .C(n_844), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g1484 ( .A(n_844), .B(n_1485), .C(n_1487), .Y(n_1484) );
INVx3_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_SL g869 ( .A(n_854), .Y(n_869) );
BUFx6f_ASAP7_75t_L g1496 ( .A(n_854), .Y(n_1496) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_858), .C(n_860), .Y(n_855) );
BUFx3_ASAP7_75t_L g908 ( .A(n_860), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g1475 ( .A(n_860), .B(n_1476), .C(n_1477), .Y(n_1475) );
AOI31xp33_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_877), .A3(n_884), .B(n_889), .Y(n_865) );
AOI211xp5_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B(n_870), .C(n_873), .Y(n_866) );
INVx2_ASAP7_75t_SL g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g1106 ( .A(n_869), .Y(n_1106) );
AOI211xp5_ASAP7_75t_L g933 ( .A1(n_870), .A2(n_934), .B(n_935), .C(n_936), .Y(n_933) );
CKINVDCx11_ASAP7_75t_R g961 ( .A(n_870), .Y(n_961) );
AOI211xp5_ASAP7_75t_L g1086 ( .A1(n_870), .A2(n_1087), .B(n_1089), .C(n_1090), .Y(n_1086) );
AOI211xp5_ASAP7_75t_L g1494 ( .A1(n_870), .A2(n_1495), .B(n_1496), .C(n_1497), .Y(n_1494) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVxp67_ASAP7_75t_L g967 ( .A(n_872), .Y(n_967) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g937 ( .A(n_875), .Y(n_937) );
AOI322xp5_ASAP7_75t_L g962 ( .A1(n_875), .A2(n_958), .A3(n_963), .B1(n_964), .B2(n_965), .C1(n_966), .C2(n_968), .Y(n_962) );
INVx2_ASAP7_75t_L g1498 ( .A(n_875), .Y(n_1498) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_878), .A2(n_880), .B1(n_881), .B2(n_883), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_878), .A2(n_881), .B1(n_940), .B2(n_941), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_878), .A2(n_1092), .B1(n_1093), .B2(n_1094), .Y(n_1091) );
AOI22xp33_ASAP7_75t_SL g1499 ( .A1(n_878), .A2(n_1093), .B1(n_1500), .B2(n_1501), .Y(n_1499) );
AND2x4_ASAP7_75t_L g881 ( .A(n_879), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g958 ( .A(n_879), .Y(n_958) );
AND2x4_ASAP7_75t_L g1093 ( .A(n_879), .B(n_882), .Y(n_1093) );
INVx5_ASAP7_75t_SL g959 ( .A(n_881), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_885), .A2(n_887), .B1(n_896), .B2(n_943), .Y(n_942) );
AOI211xp5_ASAP7_75t_L g954 ( .A1(n_885), .A2(n_955), .B(n_956), .C(n_960), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_885), .A2(n_1078), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
AOI22xp33_ASAP7_75t_SL g1502 ( .A1(n_885), .A2(n_1097), .B1(n_1463), .B2(n_1503), .Y(n_1502) );
INVx5_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx4_ASAP7_75t_L g1097 ( .A(n_888), .Y(n_1097) );
AOI31xp33_ASAP7_75t_L g1085 ( .A1(n_889), .A2(n_1086), .A3(n_1091), .B(n_1095), .Y(n_1085) );
AOI31xp33_ASAP7_75t_L g1493 ( .A1(n_889), .A2(n_1494), .A3(n_1499), .B(n_1502), .Y(n_1493) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g946 ( .A(n_893), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_920), .Y(n_906) );
AOI33xp33_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_909), .A3(n_911), .B1(n_914), .B2(n_918), .B3(n_919), .Y(n_907) );
AOI33xp33_ASAP7_75t_L g1099 ( .A1(n_908), .A2(n_919), .A3(n_1100), .B1(n_1101), .B2(n_1102), .B3(n_1103), .Y(n_1099) );
INVx3_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g1147 ( .A(n_917), .Y(n_1147) );
INVx2_ASAP7_75t_L g1023 ( .A(n_919), .Y(n_1023) );
AOI33xp33_ASAP7_75t_L g1107 ( .A1(n_921), .A2(n_1108), .A3(n_1111), .B1(n_1113), .B2(n_1114), .B3(n_1115), .Y(n_1107) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
AOI31xp33_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_939), .A3(n_942), .B(n_944), .Y(n_932) );
OAI211xp5_ASAP7_75t_L g953 ( .A1(n_944), .A2(n_954), .B(n_969), .C(n_985), .Y(n_953) );
XOR2xp5_ASAP7_75t_L g948 ( .A(n_949), .B(n_1068), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
XNOR2x1_ASAP7_75t_L g951 ( .A(n_952), .B(n_1026), .Y(n_951) );
INVx1_ASAP7_75t_L g1024 ( .A(n_953), .Y(n_1024) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_955), .A2(n_996), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
OAI31xp33_ASAP7_75t_SL g969 ( .A1(n_970), .A2(n_972), .A3(n_976), .B(n_984), .Y(n_969) );
INVx1_ASAP7_75t_L g980 ( .A(n_974), .Y(n_980) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_981), .A2(n_1016), .B1(n_1017), .B2(n_1019), .Y(n_1015) );
AOI211xp5_ASAP7_75t_L g1460 ( .A1(n_984), .A2(n_1461), .B(n_1474), .C(n_1493), .Y(n_1460) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_1008), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B1(n_991), .B2(n_992), .Y(n_987) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
OAI22xp33_ASAP7_75t_SL g994 ( .A1(n_995), .A2(n_996), .B1(n_998), .B2(n_999), .Y(n_994) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_1017), .A2(n_1140), .B1(n_1141), .B2(n_1144), .Y(n_1139) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
NAND4xp25_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1054), .C(n_1065), .D(n_1067), .Y(n_1027) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1034), .B1(n_1038), .B2(n_1041), .C(n_1044), .Y(n_1029) );
OAI21xp5_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1036), .B(n_1037), .Y(n_1034) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
XNOR2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1116), .Y(n_1070) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1107), .Y(n_1098) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
XNOR2x1_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1118), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1153), .Y(n_1118) );
NOR3xp33_ASAP7_75t_SL g1119 ( .A(n_1120), .B(n_1129), .C(n_1131), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1125), .Y(n_1120) );
OAI211xp5_ASAP7_75t_L g1160 ( .A1(n_1124), .A2(n_1161), .B(n_1163), .C(n_1164), .Y(n_1160) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx3_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_1141), .A2(n_1146), .B1(n_1147), .B2(n_1148), .Y(n_1145) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_SL g1158 ( .A(n_1159), .Y(n_1158) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
OAI221xp5_ASAP7_75t_L g1172 ( .A1(n_1173), .A2(n_1400), .B1(n_1404), .B2(n_1446), .C(n_1449), .Y(n_1172) );
AOI211xp5_ASAP7_75t_SL g1173 ( .A1(n_1174), .A2(n_1284), .B(n_1298), .C(n_1359), .Y(n_1173) );
A2O1A1Ixp33_ASAP7_75t_L g1174 ( .A1(n_1175), .A2(n_1246), .B(n_1253), .C(n_1256), .Y(n_1174) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1204), .B1(n_1206), .B2(n_1236), .Y(n_1175) );
NOR4xp25_ASAP7_75t_L g1253 ( .A(n_1176), .B(n_1220), .C(n_1236), .D(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1176), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1200), .Y(n_1176) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1177), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1177), .B(n_1260), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1177), .B(n_1201), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1197), .Y(n_1177) );
INVxp67_ASAP7_75t_SL g1249 ( .A(n_1178), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1178), .B(n_1235), .Y(n_1251) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1178), .Y(n_1266) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1178), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1178), .B(n_1201), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1191), .Y(n_1178) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1186), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1182), .B(n_1187), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1185), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1185), .Y(n_1195) );
AND2x4_ASAP7_75t_L g1188 ( .A(n_1186), .B(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1187), .B(n_1190), .Y(n_1231) );
HB1xp67_ASAP7_75t_L g1505 ( .A(n_1189), .Y(n_1505) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1194), .Y(n_1192) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_1193), .B(n_1195), .Y(n_1196) );
AND2x4_ASAP7_75t_L g1212 ( .A(n_1193), .B(n_1194), .Y(n_1212) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1196), .Y(n_1214) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1197), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1197), .B(n_1249), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1200), .B(n_1223), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1200), .B(n_1265), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1200), .B(n_1320), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1200), .B(n_1251), .Y(n_1338) );
OAI22xp33_ASAP7_75t_L g1341 ( .A1(n_1200), .A2(n_1342), .B1(n_1344), .B2(n_1347), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1378 ( .A(n_1200), .B(n_1335), .Y(n_1378) );
CKINVDCx5p33_ASAP7_75t_R g1200 ( .A(n_1201), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1201), .B(n_1233), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1201), .B(n_1248), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1201), .B(n_1222), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1201), .B(n_1265), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1201), .B(n_1271), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g1346 ( .A(n_1201), .B(n_1234), .Y(n_1346) );
AND2x4_ASAP7_75t_SL g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
INVxp67_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1220), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1216), .Y(n_1206) );
NAND2xp5_ASAP7_75t_SL g1276 ( .A(n_1207), .B(n_1277), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1207), .B(n_1243), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1207), .B(n_1254), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1207), .B(n_1255), .Y(n_1385) );
CKINVDCx6p67_ASAP7_75t_R g1207 ( .A(n_1208), .Y(n_1207) );
CKINVDCx5p33_ASAP7_75t_R g1272 ( .A(n_1208), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1208), .B(n_1216), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1208), .B(n_1275), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1208), .B(n_1277), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1208), .B(n_1217), .Y(n_1358) );
OR2x2_ASAP7_75t_L g1362 ( .A(n_1208), .B(n_1241), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1208), .B(n_1370), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1208), .B(n_1216), .Y(n_1379) );
OR2x6_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1209), .B(n_1210), .Y(n_1300) );
OAI22xp5_ASAP7_75t_SL g1210 ( .A1(n_1211), .A2(n_1213), .B1(n_1214), .B2(n_1215), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_1212), .Y(n_1290) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1214), .Y(n_1224) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1214), .Y(n_1291) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1216), .Y(n_1261) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1217), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1217), .B(n_1255), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1217), .B(n_1243), .Y(n_1269) );
BUFx6f_ASAP7_75t_L g1312 ( .A(n_1217), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1219), .Y(n_1217) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1220), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1232), .Y(n_1220) );
NOR2x1p5_ASAP7_75t_L g1320 ( .A(n_1221), .B(n_1321), .Y(n_1320) );
INVxp67_ASAP7_75t_L g1370 ( .A(n_1221), .Y(n_1370) );
INVx2_ASAP7_75t_SL g1221 ( .A(n_1222), .Y(n_1221) );
BUFx3_ASAP7_75t_L g1239 ( .A(n_1222), .Y(n_1239) );
BUFx2_ASAP7_75t_L g1260 ( .A(n_1222), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1222), .B(n_1281), .Y(n_1326) );
INVx2_ASAP7_75t_SL g1222 ( .A(n_1223), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1223), .B(n_1255), .Y(n_1275) );
OAI22xp33_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1227), .B1(n_1229), .B2(n_1230), .Y(n_1225) );
BUFx3_ASAP7_75t_L g1294 ( .A(n_1227), .Y(n_1294) );
BUFx6f_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1231), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1232), .B(n_1239), .Y(n_1304) );
INVxp67_ASAP7_75t_L g1371 ( .A(n_1232), .Y(n_1371) );
AOI311xp33_ASAP7_75t_L g1331 ( .A1(n_1233), .A2(n_1272), .A3(n_1332), .B(n_1334), .C(n_1341), .Y(n_1331) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
O2A1O1Ixp33_ASAP7_75t_L g1328 ( .A1(n_1234), .A2(n_1241), .B(n_1329), .C(n_1330), .Y(n_1328) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1235), .B(n_1266), .Y(n_1265) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1240), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_1238), .B(n_1362), .Y(n_1389) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1239), .B(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1241), .Y(n_1303) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1241), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1243), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1242), .B(n_1255), .Y(n_1277) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1243), .Y(n_1255) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1243), .Y(n_1281) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1243), .Y(n_1305) );
AOI211xp5_ASAP7_75t_SL g1318 ( .A1(n_1243), .A2(n_1319), .B(n_1322), .C(n_1328), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1245), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1250), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1248), .B(n_1283), .Y(n_1282) );
NAND3xp33_ASAP7_75t_L g1325 ( .A(n_1248), .B(n_1326), .C(n_1327), .Y(n_1325) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1248), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1248), .B(n_1252), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1252), .Y(n_1250) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1251), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1251), .B(n_1283), .Y(n_1350) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1254), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1254), .B(n_1260), .Y(n_1333) );
AOI21xp5_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1272), .B(n_1273), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1262), .B1(n_1267), .B2(n_1270), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1261), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1260), .B(n_1269), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1260), .B(n_1311), .Y(n_1310) );
INVx2_ASAP7_75t_L g1329 ( .A(n_1260), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_1260), .B(n_1336), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1264), .Y(n_1262) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1269), .Y(n_1383) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1270), .Y(n_1372) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_1272), .A2(n_1389), .B1(n_1390), .B2(n_1391), .C(n_1395), .Y(n_1388) );
A2O1A1Ixp33_ASAP7_75t_L g1273 ( .A1(n_1274), .A2(n_1276), .B(n_1278), .C(n_1280), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1277), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_1278), .A2(n_1329), .B1(n_1355), .B2(n_1356), .Y(n_1354) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
NAND2xp67_ASAP7_75t_L g1392 ( .A(n_1281), .B(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1282), .Y(n_1397) );
AOI32xp33_ASAP7_75t_L g1298 ( .A1(n_1284), .A2(n_1299), .A3(n_1318), .B1(n_1331), .B2(n_1349), .Y(n_1298) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
OAI211xp5_ASAP7_75t_L g1322 ( .A1(n_1285), .A2(n_1323), .B(n_1324), .C(n_1325), .Y(n_1322) );
INVx3_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
AOI211xp5_ASAP7_75t_L g1382 ( .A1(n_1287), .A2(n_1383), .B(n_1384), .C(n_1386), .Y(n_1382) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_1293), .A2(n_1294), .B1(n_1295), .B2(n_1296), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1403 ( .A(n_1296), .Y(n_1403) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
AOI211xp5_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1301), .B(n_1306), .C(n_1309), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g1301 ( .A1(n_1302), .A2(n_1303), .B1(n_1304), .B2(n_1305), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1305), .B(n_1307), .Y(n_1306) );
INVx3_ASAP7_75t_L g1353 ( .A(n_1305), .Y(n_1353) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1308), .Y(n_1330) );
OAI222xp33_ASAP7_75t_L g1309 ( .A1(n_1310), .A2(n_1311), .B1(n_1312), .B2(n_1313), .C1(n_1314), .C2(n_1316), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1364 ( .A1(n_1310), .A2(n_1316), .B1(n_1365), .B2(n_1367), .Y(n_1364) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1311), .Y(n_1399) );
CKINVDCx14_ASAP7_75t_R g1327 ( .A(n_1312), .Y(n_1327) );
A2O1A1Ixp33_ASAP7_75t_L g1395 ( .A1(n_1313), .A2(n_1396), .B(n_1397), .C(n_1398), .Y(n_1395) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1319), .Y(n_1394) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1323), .Y(n_1390) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1329), .Y(n_1355) );
AOI221xp5_ASAP7_75t_L g1377 ( .A1(n_1329), .A2(n_1335), .B1(n_1344), .B2(n_1378), .C(n_1379), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1329), .B(n_1357), .Y(n_1387) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
AOI21xp33_ASAP7_75t_SL g1334 ( .A1(n_1335), .A2(n_1337), .B(n_1339), .Y(n_1334) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1335), .Y(n_1363) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1338), .B(n_1343), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g1339 ( .A(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
HB1xp67_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1348), .B(n_1399), .Y(n_1398) );
A2O1A1Ixp33_ASAP7_75t_SL g1349 ( .A1(n_1350), .A2(n_1351), .B(n_1354), .C(n_1358), .Y(n_1349) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
AOI21xp33_ASAP7_75t_L g1373 ( .A1(n_1356), .A2(n_1374), .B(n_1375), .Y(n_1373) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND3xp33_ASAP7_75t_SL g1359 ( .A(n_1360), .B(n_1376), .C(n_1388), .Y(n_1359) );
AOI211xp5_ASAP7_75t_L g1360 ( .A1(n_1361), .A2(n_1363), .B(n_1364), .C(n_1373), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
NAND3xp33_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1371), .C(n_1372), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
NOR3xp33_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1380), .C(n_1382), .Y(n_1376) );
INVxp67_ASAP7_75t_SL g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
NAND2xp5_ASAP7_75t_SL g1391 ( .A(n_1392), .B(n_1394), .Y(n_1391) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1393), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_SL g1401 ( .A(n_1402), .Y(n_1401) );
BUFx2_ASAP7_75t_SL g1402 ( .A(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1405), .Y(n_1445) );
HB1xp67_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
NOR3xp33_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1409), .C(n_1428), .Y(n_1406) );
NAND4xp25_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1435), .C(n_1438), .D(n_1441), .Y(n_1428) );
CKINVDCx5p33_ASAP7_75t_R g1446 ( .A(n_1447), .Y(n_1446) );
OAI21xp5_ASAP7_75t_L g1504 ( .A1(n_1448), .A2(n_1505), .B(n_1506), .Y(n_1504) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
HB1xp67_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
NAND4xp25_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1479), .C(n_1484), .D(n_1488), .Y(n_1474) );
NAND3xp33_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1481), .C(n_1483), .Y(n_1479) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
endmodule