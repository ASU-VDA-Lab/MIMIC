module fake_jpeg_2104_n_219 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_219);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_51),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_81),
.C(n_65),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_0),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_69),
.B1(n_76),
.B2(n_75),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_60),
.B(n_67),
.Y(n_112)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_72),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_57),
.C(n_55),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_74),
.C(n_71),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_69),
.B1(n_76),
.B2(n_63),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_82),
.B1(n_60),
.B2(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_118),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_109),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_104),
.B1(n_52),
.B2(n_4),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_66),
.B1(n_58),
.B2(n_62),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_71),
.B1(n_85),
.B2(n_75),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_89),
.B(n_88),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_68),
.B(n_73),
.C(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_74),
.B1(n_64),
.B2(n_63),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_89),
.B1(n_78),
.B2(n_98),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_117),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_78),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_95),
.Y(n_120)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_25),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_131),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_122),
.A2(n_134),
.B1(n_114),
.B2(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_127),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_119),
.B(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_23),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_52),
.B1(n_4),
.B2(n_6),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_3),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_13),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_7),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_145),
.B1(n_156),
.B2(n_166),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_147),
.B(n_27),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_29),
.C(n_48),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_163),
.C(n_166),
.Y(n_171)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_15),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_14),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_165),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_30),
.C(n_46),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_33),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_172),
.B1(n_41),
.B2(n_44),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_128),
.B1(n_141),
.B2(n_122),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g173 ( 
.A(n_148),
.B(n_37),
.C(n_45),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_176),
.C(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_28),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_24),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_185),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_39),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_161),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_17),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_163),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_161),
.C(n_40),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_198),
.C(n_184),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_193),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_181),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_49),
.C(n_19),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_200),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_195),
.B(n_177),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_203),
.A2(n_205),
.B(n_168),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_194),
.C(n_202),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_176),
.B(n_179),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_190),
.C(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_170),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_211),
.C(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_187),
.B1(n_168),
.B2(n_204),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_210),
.A3(n_192),
.B1(n_173),
.B2(n_20),
.C1(n_19),
.C2(n_18),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_215),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_217),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_218),
.Y(n_219)
);


endmodule