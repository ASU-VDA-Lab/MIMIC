module fake_jpeg_14473_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

AOI21xp33_ASAP7_75t_L g10 ( 
.A1(n_6),
.A2(n_3),
.B(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_19),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_21),
.B(n_24),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_2),
.B1(n_8),
.B2(n_7),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_15),
.B1(n_9),
.B2(n_13),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_25),
.B1(n_20),
.B2(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_14),
.A2(n_2),
.B1(n_12),
.B2(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_13),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_14),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_15),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_21),
.B1(n_17),
.B2(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_31),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_36),
.B(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp67_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_36),
.Y(n_42)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_41),
.A3(n_43),
.B1(n_29),
.B2(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_44),
.Y(n_46)
);


endmodule