module real_jpeg_20718_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_0),
.B(n_40),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_0),
.A2(n_21),
.B(n_25),
.C(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_0),
.A2(n_75),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_0),
.B(n_75),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_0),
.A2(n_10),
.B(n_49),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_0),
.B(n_91),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_0),
.A2(n_21),
.B1(n_22),
.B2(n_50),
.Y(n_168)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_3),
.B(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_3),
.B(n_121),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_23),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_4),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_36),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_6),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_27),
.B(n_63),
.C(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_10),
.B(n_27),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_114),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_112),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_70),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_15),
.B(n_70),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_56),
.C(n_61),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_16),
.A2(n_17),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_18),
.B(n_39),
.C(n_43),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_31),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_24),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_20),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_24),
.B(n_25),
.C(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_42),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_22),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g59 ( 
.A1(n_26),
.A2(n_27),
.B(n_50),
.Y(n_59)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_28),
.A2(n_50),
.B(n_64),
.C(n_125),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_35),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_74),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_75),
.B(n_79),
.C(n_80),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_45),
.B(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_46),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_52),
.B(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_48),
.B(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_50),
.B(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_50),
.B(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_51),
.B(n_121),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_54),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_58),
.A2(n_60),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_61),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_63),
.B(n_69),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_63),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_67),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_66),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_67),
.B(n_150),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_96),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_83),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_79),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_95),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_90),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_93),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_110),
.B2(n_111),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_109),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_104)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_172),
.B(n_178),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_155),
.B(n_171),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_141),
.B(n_154),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_130),
.B(n_140),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_122),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_126),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_135),
.B(n_139),
.Y(n_130)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_148),
.C(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_157),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B1(n_162),
.B2(n_170),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_169),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_173),
.B(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);


endmodule