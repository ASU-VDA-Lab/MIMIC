module fake_jpeg_3227_n_77 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_25),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_23),
.B(n_26),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_23),
.B(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_45),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_22),
.B(n_11),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_39),
.B1(n_27),
.B2(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_51),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_21),
.B(n_36),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_21),
.B1(n_22),
.B2(n_3),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_49),
.C(n_47),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_1),
.C(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVxp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_45),
.B(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_65),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_12),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_56),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_69),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_66),
.C(n_67),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_72),
.B(n_66),
.Y(n_74)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_20),
.A3(n_18),
.B1(n_17),
.B2(n_13),
.C1(n_8),
.C2(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_5),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_71),
.Y(n_77)
);


endmodule