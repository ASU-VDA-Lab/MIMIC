module fake_jpeg_29291_n_265 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_27),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_18),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_18),
.Y(n_86)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_24),
.B1(n_34),
.B2(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_63),
.B1(n_58),
.B2(n_43),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_93),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_34),
.B1(n_35),
.B2(n_32),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_63),
.B1(n_51),
.B2(n_58),
.Y(n_100)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_88),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_28),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_35),
.B1(n_23),
.B2(n_30),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_19),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_96),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_38),
.C(n_28),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_41),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_19),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_105),
.Y(n_151)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_59),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_103),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_122),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_54),
.CON(n_103),
.SN(n_103)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_69),
.B1(n_74),
.B2(n_80),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_51),
.C(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_106),
.B(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_33),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_31),
.B(n_29),
.C(n_26),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_116),
.B(n_128),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_60),
.B1(n_47),
.B2(n_31),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_121),
.B1(n_79),
.B2(n_74),
.Y(n_141)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_29),
.B1(n_23),
.B2(n_2),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_23),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_14),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_0),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_90),
.B1(n_79),
.B2(n_81),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_103),
.B1(n_110),
.B2(n_108),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_140),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_94),
.B(n_90),
.C(n_81),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_83),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_144),
.B1(n_151),
.B2(n_95),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_83),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_107),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_160),
.B(n_161),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_174),
.B1(n_123),
.B2(n_80),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_137),
.C(n_133),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_127),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_169),
.A3(n_19),
.B1(n_67),
.B2(n_120),
.C1(n_131),
.C2(n_152),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_78),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_172),
.B(n_175),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_101),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_177),
.C(n_139),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_117),
.B(n_112),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_121),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_100),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_129),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_149),
.A2(n_117),
.B(n_124),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_182),
.Y(n_200)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_138),
.B(n_140),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_185),
.B(n_198),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_151),
.B(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_151),
.B1(n_141),
.B2(n_95),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_177),
.B1(n_173),
.B2(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_192),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_153),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_114),
.B1(n_69),
.B2(n_98),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_196),
.A2(n_134),
.B1(n_166),
.B2(n_167),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_135),
.B(n_146),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_154),
.C(n_148),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_164),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_180),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_216),
.B1(n_191),
.B2(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_206),
.B1(n_218),
.B2(n_183),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_169),
.B1(n_165),
.B2(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_159),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_217),
.C(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_201),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_214),
.A2(n_199),
.B(n_186),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_182),
.B1(n_147),
.B2(n_142),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_164),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_147),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_192),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_192),
.CI(n_184),
.CON(n_221),
.SN(n_221)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_222),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_206),
.B1(n_203),
.B2(n_202),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_185),
.B(n_198),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_230),
.A2(n_219),
.B(n_217),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_202),
.C(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_209),
.C(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_233),
.B1(n_237),
.B2(n_226),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_215),
.B1(n_202),
.B2(n_187),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_239),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_191),
.B1(n_209),
.B2(n_216),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_227),
.C(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_146),
.C(n_1),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_222),
.C(n_225),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_221),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_247),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_224),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_238),
.A3(n_230),
.B1(n_240),
.B2(n_5),
.C1(n_7),
.C2(n_8),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_238),
.C(n_2),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_4),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_0),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_253),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_11),
.B(n_8),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_258),
.A2(n_252),
.B1(n_8),
.B2(n_9),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_259),
.A2(n_260),
.B1(n_256),
.B2(n_255),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_5),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_169),
.C2(n_165),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_259),
.Y(n_265)
);


endmodule