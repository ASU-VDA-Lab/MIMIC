module real_aes_638_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_0), .B(n_120), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_1), .A2(n_133), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_2), .B(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_3), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g127 ( .A(n_4), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_5), .B(n_142), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_6), .B(n_129), .Y(n_502) );
INVx1_ASAP7_75t_L g478 ( .A(n_7), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g812 ( .A(n_8), .Y(n_812) );
XNOR2xp5_ASAP7_75t_L g104 ( .A(n_9), .B(n_105), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_10), .Y(n_493) );
NAND2xp33_ASAP7_75t_L g205 ( .A(n_11), .B(n_140), .Y(n_205) );
INVx2_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
AOI221x1_ASAP7_75t_L g149 ( .A1(n_13), .A2(n_25), .B1(n_120), .B2(n_133), .C(n_150), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_14), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_15), .B(n_120), .Y(n_201) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_16), .A2(n_199), .B(n_200), .Y(n_198) );
INVx1_ASAP7_75t_L g510 ( .A(n_17), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_18), .B(n_147), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_19), .B(n_142), .Y(n_193) );
AO21x1_ASAP7_75t_L g119 ( .A1(n_20), .A2(n_120), .B(n_128), .Y(n_119) );
INVx1_ASAP7_75t_L g443 ( .A(n_21), .Y(n_443) );
INVx1_ASAP7_75t_L g508 ( .A(n_22), .Y(n_508) );
INVx1_ASAP7_75t_SL g559 ( .A(n_23), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_24), .B(n_121), .Y(n_522) );
NAND2x1_ASAP7_75t_L g160 ( .A(n_26), .B(n_142), .Y(n_160) );
AOI33xp33_ASAP7_75t_L g546 ( .A1(n_27), .A2(n_54), .A3(n_459), .B1(n_466), .B2(n_547), .B3(n_548), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_28), .A2(n_103), .B1(n_805), .B2(n_816), .C1(n_830), .C2(n_832), .Y(n_102) );
AOI22xp5_ASAP7_75t_SL g819 ( .A1(n_28), .A2(n_820), .B1(n_823), .B2(n_824), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_28), .Y(n_824) );
NAND2x1_ASAP7_75t_L g219 ( .A(n_29), .B(n_140), .Y(n_219) );
INVx1_ASAP7_75t_L g486 ( .A(n_30), .Y(n_486) );
OR2x2_ASAP7_75t_L g130 ( .A(n_31), .B(n_88), .Y(n_130) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_31), .A2(n_88), .B(n_131), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_32), .B(n_457), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_33), .B(n_140), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_34), .B(n_142), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_35), .A2(n_65), .B1(n_821), .B2(n_822), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_35), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_36), .B(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_37), .A2(n_133), .B(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g126 ( .A(n_38), .B(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g134 ( .A(n_38), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g465 ( .A(n_38), .Y(n_465) );
OR2x6_ASAP7_75t_L g441 ( .A(n_39), .B(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_40), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_41), .B(n_120), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_42), .B(n_457), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_43), .A2(n_129), .B1(n_165), .B2(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_44), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_45), .B(n_121), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_46), .A2(n_96), .B1(n_106), .B2(n_107), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_46), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_47), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_48), .B(n_140), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_49), .B(n_199), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_50), .B(n_121), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_51), .A2(n_133), .B(n_218), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_52), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_53), .B(n_140), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_55), .B(n_121), .Y(n_471) );
INVx1_ASAP7_75t_L g123 ( .A(n_56), .Y(n_123) );
INVx1_ASAP7_75t_L g137 ( .A(n_56), .Y(n_137) );
AND2x2_ASAP7_75t_L g472 ( .A(n_57), .B(n_147), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_58), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_59), .A2(n_77), .B1(n_457), .B2(n_463), .C(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_60), .B(n_457), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_61), .B(n_142), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_62), .B(n_165), .Y(n_495) );
AOI21xp5_ASAP7_75t_SL g530 ( .A1(n_63), .A2(n_463), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_64), .A2(n_133), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_65), .Y(n_821) );
INVx1_ASAP7_75t_L g505 ( .A(n_66), .Y(n_505) );
AO21x1_ASAP7_75t_L g132 ( .A1(n_67), .A2(n_133), .B(n_138), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_68), .B(n_120), .Y(n_210) );
INVx1_ASAP7_75t_L g469 ( .A(n_69), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_70), .A2(n_104), .B1(n_796), .B2(n_801), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_71), .B(n_120), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_72), .A2(n_463), .B(n_468), .Y(n_462) );
AND2x2_ASAP7_75t_L g177 ( .A(n_73), .B(n_148), .Y(n_177) );
INVx1_ASAP7_75t_L g125 ( .A(n_74), .Y(n_125) );
INVx1_ASAP7_75t_L g135 ( .A(n_74), .Y(n_135) );
AND2x2_ASAP7_75t_L g223 ( .A(n_75), .B(n_164), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_76), .B(n_457), .Y(n_549) );
AND2x2_ASAP7_75t_L g561 ( .A(n_78), .B(n_164), .Y(n_561) );
INVx1_ASAP7_75t_L g506 ( .A(n_79), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_80), .A2(n_463), .B(n_558), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_81), .A2(n_463), .B(n_521), .C(n_525), .Y(n_520) );
INVx1_ASAP7_75t_L g444 ( .A(n_82), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_83), .B(n_120), .Y(n_195) );
AND2x2_ASAP7_75t_L g208 ( .A(n_84), .B(n_164), .Y(n_208) );
AND2x2_ASAP7_75t_SL g528 ( .A(n_85), .B(n_164), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_86), .A2(n_463), .B1(n_544), .B2(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g128 ( .A(n_87), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g167 ( .A(n_89), .B(n_164), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_90), .B(n_140), .Y(n_194) );
INVx1_ASAP7_75t_L g532 ( .A(n_91), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_92), .B(n_142), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_93), .B(n_140), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_94), .A2(n_133), .B(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g550 ( .A(n_95), .B(n_164), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_96), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_97), .B(n_142), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_98), .A2(n_484), .B(n_485), .C(n_488), .Y(n_483) );
BUFx2_ASAP7_75t_L g813 ( .A(n_99), .Y(n_813) );
BUFx2_ASAP7_75t_SL g838 ( .A(n_99), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_100), .A2(n_133), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_101), .B(n_121), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_108), .B(n_795), .Y(n_103) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_436), .B1(n_445), .B2(n_791), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_111), .A2(n_797), .B1(n_799), .B2(n_800), .Y(n_796) );
XOR2x1_ASAP7_75t_SL g818 ( .A(n_111), .B(n_819), .Y(n_818) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_335), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_272), .C(n_295), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_224), .C(n_241), .Y(n_113) );
OAI31xp33_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_154), .A3(n_178), .B(n_185), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_115), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_146), .Y(n_116) );
AND2x4_ASAP7_75t_L g227 ( .A(n_117), .B(n_146), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_117), .B(n_169), .Y(n_256) );
AND2x4_ASAP7_75t_L g258 ( .A(n_117), .B(n_252), .Y(n_258) );
AND2x2_ASAP7_75t_L g389 ( .A(n_117), .B(n_182), .Y(n_389) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g234 ( .A(n_118), .Y(n_234) );
OAI21x1_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_132), .B(n_144), .Y(n_118) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_126), .Y(n_120) );
INVx1_ASAP7_75t_L g487 ( .A(n_121), .Y(n_487) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
AND2x6_ASAP7_75t_L g140 ( .A(n_122), .B(n_135), .Y(n_140) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g142 ( .A(n_124), .B(n_137), .Y(n_142) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx5_ASAP7_75t_L g143 ( .A(n_126), .Y(n_143) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_126), .Y(n_488) );
AND2x2_ASAP7_75t_L g136 ( .A(n_127), .B(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_127), .Y(n_460) );
INVx1_ASAP7_75t_L g145 ( .A(n_128), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_129), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_SL g189 ( .A(n_129), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_129), .A2(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_129), .B(n_143), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_129), .A2(n_530), .B(n_534), .Y(n_529) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_130), .B(n_131), .Y(n_148) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
BUFx3_ASAP7_75t_L g461 ( .A(n_134), .Y(n_461) );
INVx2_ASAP7_75t_L g467 ( .A(n_135), .Y(n_467) );
AND2x4_ASAP7_75t_L g463 ( .A(n_136), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g459 ( .A(n_137), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_141), .B(n_143), .Y(n_138) );
INVxp67_ASAP7_75t_L g509 ( .A(n_140), .Y(n_509) );
INVxp67_ASAP7_75t_L g511 ( .A(n_142), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_143), .A2(n_151), .B(n_152), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_143), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_143), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_143), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_143), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_143), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_143), .A2(n_219), .B(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_143), .A2(n_469), .B(n_470), .C(n_471), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_143), .A2(n_470), .B(n_478), .C(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_143), .A2(n_522), .B(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_143), .A2(n_470), .B(n_532), .C(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g544 ( .A(n_143), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_SL g558 ( .A1(n_143), .A2(n_470), .B(n_559), .C(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g168 ( .A(n_146), .B(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_146), .B(n_233), .Y(n_325) );
AND2x2_ASAP7_75t_L g331 ( .A(n_146), .B(n_170), .Y(n_331) );
AND2x2_ASAP7_75t_L g420 ( .A(n_146), .B(n_421), .Y(n_420) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_153), .Y(n_146) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_147), .A2(n_149), .B(n_153), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_147), .A2(n_210), .B(n_211), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_147), .Y(n_222) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_SL g402 ( .A(n_154), .Y(n_402) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_168), .Y(n_154) );
BUFx2_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
AND2x2_ASAP7_75t_L g265 ( .A(n_155), .B(n_169), .Y(n_265) );
AND2x2_ASAP7_75t_L g314 ( .A(n_155), .B(n_170), .Y(n_314) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g271 ( .A(n_156), .B(n_170), .Y(n_271) );
INVxp67_ASAP7_75t_L g283 ( .A(n_156), .Y(n_283) );
BUFx3_ASAP7_75t_L g328 ( .A(n_156), .Y(n_328) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_163), .B(n_167), .Y(n_156) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_157), .A2(n_163), .B(n_167), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_163), .A2(n_171), .B(n_177), .Y(n_170) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_163), .A2(n_171), .B(n_177), .Y(n_184) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_163), .A2(n_455), .B(n_472), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_163), .A2(n_164), .B1(n_483), .B2(n_489), .Y(n_482) );
AO21x2_ASAP7_75t_L g611 ( .A1(n_163), .A2(n_455), .B(n_472), .Y(n_611) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_165), .B(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx4f_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
OAI31xp33_ASAP7_75t_L g224 ( .A1(n_168), .A2(n_225), .A3(n_230), .B(n_235), .Y(n_224) );
AND2x2_ASAP7_75t_L g232 ( .A(n_169), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g251 ( .A(n_170), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_172), .B(n_176), .Y(n_171) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_178), .A2(n_300), .A3(n_329), .B1(n_334), .B2(n_426), .C1(n_429), .C2(n_430), .Y(n_425) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_179), .B(n_271), .Y(n_276) );
NAND2x1_ASAP7_75t_L g313 ( .A(n_179), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g357 ( .A(n_179), .B(n_261), .Y(n_357) );
INVx1_ASAP7_75t_SL g371 ( .A(n_179), .Y(n_371) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g252 ( .A(n_180), .Y(n_252) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_180), .Y(n_395) );
AND2x2_ASAP7_75t_L g324 ( .A(n_181), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_181), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_SL g181 ( .A(n_182), .B(n_183), .Y(n_181) );
BUFx2_ASAP7_75t_L g229 ( .A(n_182), .Y(n_229) );
INVx1_ASAP7_75t_L g421 ( .A(n_182), .Y(n_421) );
OR2x2_ASAP7_75t_L g288 ( .A(n_183), .B(n_233), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_183), .B(n_258), .Y(n_322) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x4_ASAP7_75t_L g261 ( .A(n_184), .B(n_233), .Y(n_261) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_206), .Y(n_185) );
INVxp67_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g317 ( .A(n_187), .Y(n_317) );
OR2x2_ASAP7_75t_L g344 ( .A(n_187), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_198), .Y(n_187) );
NOR2x1_ASAP7_75t_SL g238 ( .A(n_188), .B(n_207), .Y(n_238) );
AND2x2_ASAP7_75t_L g245 ( .A(n_188), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g417 ( .A(n_188), .B(n_279), .Y(n_417) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_196), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_189), .B(n_197), .Y(n_196) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_189), .A2(n_190), .B(n_196), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_195), .Y(n_190) );
OR2x2_ASAP7_75t_L g239 ( .A(n_198), .B(n_240), .Y(n_239) );
BUFx3_ASAP7_75t_L g248 ( .A(n_198), .Y(n_248) );
INVx2_ASAP7_75t_L g279 ( .A(n_198), .Y(n_279) );
INVx1_ASAP7_75t_L g320 ( .A(n_198), .Y(n_320) );
AND2x2_ASAP7_75t_L g351 ( .A(n_198), .B(n_207), .Y(n_351) );
AND2x2_ASAP7_75t_L g382 ( .A(n_198), .B(n_309), .Y(n_382) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_199), .A2(n_476), .B(n_480), .Y(n_475) );
INVx2_ASAP7_75t_SL g525 ( .A(n_199), .Y(n_525) );
AND2x2_ASAP7_75t_L g278 ( .A(n_206), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_206), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_SL g381 ( .A(n_206), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g386 ( .A(n_206), .B(n_248), .Y(n_386) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_215), .Y(n_206) );
INVx5_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_207), .B(n_240), .Y(n_318) );
BUFx2_ASAP7_75t_L g378 ( .A(n_207), .Y(n_378) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
INVx4_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
AND2x2_ASAP7_75t_L g363 ( .A(n_215), .B(n_246), .Y(n_363) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_222), .B(n_223), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_222), .A2(n_555), .B(n_561), .Y(n_554) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_226), .A2(n_353), .B1(n_356), .B2(n_358), .C(n_359), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AND2x2_ASAP7_75t_L g374 ( .A(n_227), .B(n_265), .Y(n_374) );
INVx1_ASAP7_75t_SL g400 ( .A(n_227), .Y(n_400) );
AND2x2_ASAP7_75t_L g385 ( .A(n_228), .B(n_357), .Y(n_385) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_229), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
AND2x2_ASAP7_75t_L g254 ( .A(n_231), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g260 ( .A(n_231), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g284 ( .A(n_232), .Y(n_284) );
AND2x2_ASAP7_75t_L g342 ( .A(n_232), .B(n_270), .Y(n_342) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
BUFx2_ASAP7_75t_L g267 ( .A(n_234), .Y(n_267) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
OR2x2_ASAP7_75t_L g431 ( .A(n_239), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g247 ( .A(n_240), .Y(n_247) );
AND2x4_ASAP7_75t_L g303 ( .A(n_240), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_240), .B(n_308), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_240), .B(n_246), .Y(n_345) );
AND2x2_ASAP7_75t_L g405 ( .A(n_240), .B(n_308), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_249), .B1(n_262), .B2(n_264), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_242), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND3x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .C(n_248), .Y(n_244) );
AND2x4_ASAP7_75t_L g262 ( .A(n_245), .B(n_263), .Y(n_262) );
INVx4_ASAP7_75t_L g302 ( .A(n_246), .Y(n_302) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_246), .B(n_303), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_247), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g347 ( .A(n_248), .Y(n_347) );
AOI322xp5_ASAP7_75t_L g412 ( .A1(n_248), .A2(n_377), .A3(n_413), .B1(n_415), .B2(n_418), .C1(n_422), .C2(n_423), .Y(n_412) );
NAND4xp25_ASAP7_75t_SL g249 ( .A(n_250), .B(n_253), .C(n_257), .D(n_259), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_SL g379 ( .A(n_251), .B(n_267), .Y(n_379) );
BUFx2_ASAP7_75t_L g270 ( .A(n_252), .Y(n_270) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g394 ( .A(n_255), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g408 ( .A(n_256), .B(n_283), .Y(n_408) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g274 ( .A(n_258), .B(n_275), .Y(n_274) );
OAI211xp5_ASAP7_75t_L g326 ( .A1(n_258), .A2(n_327), .B(n_329), .C(n_332), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_258), .B(n_265), .Y(n_384) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_260), .A2(n_342), .B1(n_343), .B2(n_346), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_261), .A2(n_297), .B1(n_301), .B2(n_305), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_261), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_261), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_261), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g428 ( .A(n_261), .Y(n_428) );
INVx1_ASAP7_75t_L g367 ( .A(n_262), .Y(n_367) );
OAI21xp33_ASAP7_75t_SL g264 ( .A1(n_265), .A2(n_266), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_265), .B(n_270), .Y(n_424) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g360 ( .A(n_267), .B(n_271), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_269), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g427 ( .A(n_270), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g401 ( .A(n_271), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_277), .C(n_280), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI22xp33_ASAP7_75t_SL g387 ( .A1(n_275), .A2(n_306), .B1(n_353), .B2(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_279), .B(n_302), .Y(n_310) );
OR2x2_ASAP7_75t_L g339 ( .A(n_279), .B(n_340), .Y(n_339) );
OAI21xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_285), .B(n_289), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g300 ( .A(n_283), .Y(n_300) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI211xp5_ASAP7_75t_SL g338 ( .A1(n_286), .A2(n_339), .B(n_341), .C(n_349), .Y(n_338) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp67_ASAP7_75t_SL g372 ( .A(n_291), .B(n_318), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_291), .Y(n_375) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_293), .B(n_302), .Y(n_432) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g304 ( .A(n_294), .Y(n_304) );
INVx2_ASAP7_75t_L g309 ( .A(n_294), .Y(n_309) );
NAND4xp25_ASAP7_75t_L g295 ( .A(n_296), .B(n_311), .C(n_323), .D(n_326), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_299), .A2(n_431), .B1(n_433), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x4_ASAP7_75t_L g398 ( .A(n_302), .B(n_328), .Y(n_398) );
AND2x2_ASAP7_75t_L g319 ( .A(n_303), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g340 ( .A(n_303), .Y(n_340) );
AND2x2_ASAP7_75t_L g350 ( .A(n_303), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_310), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_309), .Y(n_364) );
INVx1_ASAP7_75t_L g354 ( .A(n_310), .Y(n_354) );
AOI32xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .A3(n_318), .B1(n_319), .B2(n_321), .Y(n_311) );
OAI21xp33_ASAP7_75t_L g359 ( .A1(n_312), .A2(n_360), .B(n_361), .Y(n_359) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_315), .A2(n_392), .B1(n_394), .B2(n_396), .C(n_399), .Y(n_391) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g376 ( .A(n_317), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g334 ( .A(n_318), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_319), .A2(n_357), .B1(n_407), .B2(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g333 ( .A(n_320), .Y(n_333) );
AND2x2_ASAP7_75t_L g411 ( .A(n_320), .B(n_364), .Y(n_411) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_327), .B(n_379), .Y(n_414) );
INVx1_ASAP7_75t_L g433 ( .A(n_327), .Y(n_433) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g335 ( .A(n_336), .B(n_390), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_380), .Y(n_336) );
NOR3xp33_ASAP7_75t_SL g337 ( .A(n_338), .B(n_352), .C(n_365), .Y(n_337) );
INVx1_ASAP7_75t_L g355 ( .A(n_340), .Y(n_355) );
INVx1_ASAP7_75t_SL g366 ( .A(n_342), .Y(n_366) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g348 ( .A(n_345), .Y(n_348) );
INVx2_ASAP7_75t_L g358 ( .A(n_346), .Y(n_358) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x4_ASAP7_75t_L g404 ( .A(n_347), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g422 ( .A(n_351), .B(n_405), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
AOI32xp33_ASAP7_75t_L g373 ( .A1(n_362), .A2(n_374), .A3(n_375), .B1(n_376), .B2(n_379), .Y(n_373) );
NOR2xp33_ASAP7_75t_SL g392 ( .A(n_362), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g393 ( .A(n_364), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_368), .C(n_373), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g429 ( .A(n_377), .B(n_417), .Y(n_429) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_378), .B(n_417), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B1(n_385), .B2(n_386), .C(n_387), .Y(n_380) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g388 ( .A(n_389), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_391), .B(n_406), .C(n_412), .D(n_425), .Y(n_390) );
INVxp33_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_402), .C(n_403), .Y(n_399) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
CKINVDCx11_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
INVx4_ASAP7_75t_SL g800 ( .A(n_437), .Y(n_800) );
INVx3_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
AND2x6_ASAP7_75t_SL g439 ( .A(n_440), .B(n_441), .Y(n_439) );
OR2x6_ASAP7_75t_SL g793 ( .A(n_440), .B(n_794), .Y(n_793) );
OR2x2_ASAP7_75t_L g804 ( .A(n_440), .B(n_441), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_440), .B(n_794), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_441), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx2_ASAP7_75t_L g799 ( .A(n_445), .Y(n_799) );
NAND4xp75_ASAP7_75t_L g445 ( .A(n_446), .B(n_663), .C(n_708), .D(n_777), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_623), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_579), .C(n_604), .Y(n_448) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_497), .B1(n_535), .B2(n_551), .C1(n_566), .C2(n_573), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_473), .Y(n_451) );
AND2x2_ASAP7_75t_L g788 ( .A(n_452), .B(n_602), .Y(n_788) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_454), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_454), .B(n_481), .Y(n_578) );
INVx3_ASAP7_75t_L g593 ( .A(n_454), .Y(n_593) );
AND2x2_ASAP7_75t_L g726 ( .A(n_454), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_462), .Y(n_455) );
INVx1_ASAP7_75t_L g496 ( .A(n_457), .Y(n_496) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g517 ( .A(n_458), .Y(n_517) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
OR2x6_ASAP7_75t_L g470 ( .A(n_459), .B(n_467), .Y(n_470) );
INVxp33_ASAP7_75t_L g547 ( .A(n_459), .Y(n_547) );
INVx1_ASAP7_75t_L g518 ( .A(n_461), .Y(n_518) );
INVxp67_ASAP7_75t_L g494 ( .A(n_463), .Y(n_494) );
NOR2x1p5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g548 ( .A(n_466), .Y(n_548) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g484 ( .A(n_470), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_470), .A2(n_487), .B1(n_505), .B2(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g524 ( .A(n_470), .Y(n_524) );
AND2x2_ASAP7_75t_L g656 ( .A(n_473), .B(n_609), .Y(n_656) );
AND2x2_ASAP7_75t_L g658 ( .A(n_473), .B(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g693 ( .A(n_473), .Y(n_693) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_481), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g576 ( .A(n_475), .Y(n_576) );
INVx1_ASAP7_75t_L g595 ( .A(n_475), .Y(n_595) );
AND2x4_ASAP7_75t_L g602 ( .A(n_475), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_475), .B(n_541), .Y(n_618) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_475), .Y(n_727) );
INVx1_ASAP7_75t_L g737 ( .A(n_475), .Y(n_737) );
INVx1_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
INVx2_ASAP7_75t_L g590 ( .A(n_481), .Y(n_590) );
INVx1_ASAP7_75t_L g671 ( .A(n_481), .Y(n_671) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_SL g498 ( .A(n_499), .B(n_526), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_499), .B(n_553), .Y(n_646) );
INVx2_ASAP7_75t_L g667 ( .A(n_499), .Y(n_667) );
AND2x2_ASAP7_75t_L g675 ( .A(n_499), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_513), .Y(n_499) );
AND2x4_ASAP7_75t_L g565 ( .A(n_500), .B(n_514), .Y(n_565) );
INVx1_ASAP7_75t_L g572 ( .A(n_500), .Y(n_572) );
AND2x2_ASAP7_75t_L g748 ( .A(n_500), .B(n_554), .Y(n_748) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g586 ( .A(n_501), .B(n_514), .Y(n_586) );
INVx2_ASAP7_75t_L g622 ( .A(n_501), .Y(n_622) );
AND2x2_ASAP7_75t_L g701 ( .A(n_501), .B(n_554), .Y(n_701) );
NOR2x1_ASAP7_75t_SL g744 ( .A(n_501), .B(n_527), .Y(n_744) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_507), .B(n_512), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g598 ( .A(n_514), .B(n_527), .Y(n_598) );
INVx1_ASAP7_75t_L g614 ( .A(n_514), .Y(n_614) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_514), .Y(n_722) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .C(n_519), .Y(n_516) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_525), .A2(n_542), .B(n_550), .Y(n_541) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_525), .A2(n_542), .B(n_550), .Y(n_591) );
AND2x2_ASAP7_75t_L g585 ( .A(n_526), .B(n_586), .Y(n_585) );
OR2x6_ASAP7_75t_L g666 ( .A(n_526), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g704 ( .A(n_526), .B(n_701), .Y(n_704) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx4_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_527), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g633 ( .A(n_527), .Y(n_633) );
OR2x2_ASAP7_75t_L g639 ( .A(n_527), .B(n_554), .Y(n_639) );
AND2x4_ASAP7_75t_L g653 ( .A(n_527), .B(n_614), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_527), .B(n_622), .Y(n_654) );
OR2x6_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g698 ( .A(n_538), .B(n_617), .Y(n_698) );
BUFx2_ASAP7_75t_L g750 ( .A(n_538), .Y(n_750) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g781 ( .A(n_540), .B(n_693), .Y(n_781) );
INVx2_ASAP7_75t_L g575 ( .A(n_541), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_543), .B(n_549), .Y(n_542) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_562), .Y(n_551) );
AND2x2_ASAP7_75t_L g597 ( .A(n_552), .B(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_SL g582 ( .A(n_553), .B(n_572), .Y(n_582) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g570 ( .A(n_554), .Y(n_570) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_554), .Y(n_676) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_554), .Y(n_743) );
INVx1_ASAP7_75t_L g783 ( .A(n_554), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
BUFx2_ASAP7_75t_L g697 ( .A(n_562), .Y(n_697) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x4_ASAP7_75t_L g613 ( .A(n_563), .B(n_614), .Y(n_613) );
NOR2xp67_ASAP7_75t_SL g645 ( .A(n_563), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g718 ( .A(n_563), .B(n_701), .Y(n_718) );
AND2x4_ASAP7_75t_SL g721 ( .A(n_563), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g770 ( .A(n_563), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g637 ( .A(n_564), .Y(n_637) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g632 ( .A(n_565), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_565), .B(n_630), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_565), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_565), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g715 ( .A(n_569), .B(n_716), .Y(n_715) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g631 ( .A(n_570), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
AND2x2_ASAP7_75t_L g749 ( .A(n_574), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g757 ( .A(n_574), .B(n_686), .Y(n_757) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g626 ( .A(n_575), .B(n_611), .Y(n_626) );
AND2x4_ASAP7_75t_L g659 ( .A(n_575), .B(n_593), .Y(n_659) );
INVx1_ASAP7_75t_L g776 ( .A(n_575), .Y(n_776) );
AND2x2_ASAP7_75t_L g662 ( .A(n_577), .B(n_602), .Y(n_662) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g683 ( .A(n_578), .B(n_618), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_587), .B1(n_596), .B2(n_599), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .B(n_585), .Y(n_580) );
OAI22xp5_ASAP7_75t_SL g762 ( .A1(n_581), .A2(n_650), .B1(n_758), .B2(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_582), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g651 ( .A(n_582), .B(n_583), .Y(n_651) );
AND2x2_ASAP7_75t_SL g681 ( .A(n_582), .B(n_653), .Y(n_681) );
AOI211xp5_ASAP7_75t_SL g769 ( .A1(n_582), .A2(n_770), .B(n_772), .C(n_773), .Y(n_769) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_583), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_583), .B(n_629), .Y(n_755) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g660 ( .A(n_585), .Y(n_660) );
INVx2_ASAP7_75t_L g716 ( .A(n_586), .Y(n_716) );
AND2x2_ASAP7_75t_L g790 ( .A(n_586), .B(n_783), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_587), .A2(n_739), .B(n_745), .Y(n_738) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_592), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g725 ( .A(n_589), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g735 ( .A(n_589), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g642 ( .A(n_590), .B(n_595), .Y(n_642) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_590), .B(n_611), .Y(n_644) );
AND2x2_ASAP7_75t_L g686 ( .A(n_590), .B(n_611), .Y(n_686) );
INVx2_ASAP7_75t_L g603 ( .A(n_591), .Y(n_603) );
AND2x4_ASAP7_75t_L g609 ( .A(n_591), .B(n_610), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx3_ASAP7_75t_L g601 ( .A(n_593), .Y(n_601) );
INVx3_ASAP7_75t_L g607 ( .A(n_594), .Y(n_607) );
BUFx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g784 ( .A1(n_598), .A2(n_704), .B(n_780), .Y(n_784) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g616 ( .A(n_601), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_601), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_601), .B(n_676), .Y(n_691) );
OR2x2_ASAP7_75t_L g706 ( .A(n_601), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g713 ( .A(n_601), .B(n_617), .Y(n_713) );
AND2x2_ASAP7_75t_L g669 ( .A(n_602), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g685 ( .A(n_602), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g702 ( .A(n_602), .B(n_671), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_612), .B1(n_615), .B2(n_619), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp67_ASAP7_75t_L g679 ( .A(n_607), .B(n_608), .Y(n_679) );
NOR2xp67_ASAP7_75t_SL g717 ( .A(n_607), .B(n_625), .Y(n_717) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2x1_ASAP7_75t_L g736 ( .A(n_611), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g620 ( .A(n_613), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g684 ( .A(n_613), .B(n_630), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_613), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g787 ( .A(n_621), .B(n_653), .Y(n_787) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2x1_ASAP7_75t_L g732 ( .A(n_622), .B(n_733), .Y(n_732) );
NOR2xp67_ASAP7_75t_SL g623 ( .A(n_624), .B(n_647), .Y(n_623) );
OAI211xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_634), .C(n_643), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_625), .A2(n_678), .B(n_688), .C(n_692), .Y(n_687) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g767 ( .A(n_626), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g678 ( .A(n_630), .B(n_654), .Y(n_678) );
AND2x2_ASAP7_75t_L g765 ( .A(n_630), .B(n_744), .Y(n_765) );
INVx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g733 ( .A(n_633), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_640), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_637), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g707 ( .A(n_642), .Y(n_707) );
NAND2xp33_ASAP7_75t_SL g643 ( .A(n_644), .B(n_645), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_655), .B1(n_657), .B2(n_660), .C(n_661), .Y(n_647) );
NOR4xp25_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .C(n_652), .D(n_654), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g766 ( .A(n_653), .B(n_729), .Y(n_766) );
INVx2_ASAP7_75t_L g772 ( .A(n_653), .Y(n_772) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_656), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g759 ( .A(n_659), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND4xp75_ASAP7_75t_L g664 ( .A(n_665), .B(n_687), .C(n_694), .D(n_703), .Y(n_664) );
OA211x2_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_672), .C(n_680), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_666), .B(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g760 ( .A(n_670), .Y(n_760) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g768 ( .A(n_671), .Y(n_768) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_673), .B(n_679), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g729 ( .A(n_676), .Y(n_729) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_684), .B2(n_685), .Y(n_680) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g789 ( .A1(n_684), .A2(n_735), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_SL g763 ( .A(n_685), .Y(n_763) );
NAND2x1p5_ASAP7_75t_L g775 ( .A(n_686), .B(n_776), .Y(n_775) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_699), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVxp67_ASAP7_75t_L g761 ( .A(n_697), .Y(n_761) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_701), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_702), .A2(n_765), .B1(n_787), .B2(n_788), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND3x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_751), .C(n_764), .Y(n_709) );
NOR3x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_723), .C(n_738), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_719), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_717), .B2(n_718), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_728), .B1(n_730), .B2(n_734), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g782 ( .A(n_732), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
INVxp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g771 ( .A(n_748), .Y(n_771) );
OAI21xp5_ASAP7_75t_SL g779 ( .A1(n_749), .A2(n_780), .B(n_782), .Y(n_779) );
NOR2x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_762), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .B1(n_758), .B2(n_761), .Y(n_752) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
O2A1O1Ixp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B(n_767), .C(n_769), .Y(n_764) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NOR2x1_ASAP7_75t_SL g777 ( .A(n_778), .B(n_785), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_784), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g785 ( .A(n_786), .B(n_789), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_792), .Y(n_798) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
BUFx4f_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
INVx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_814), .Y(n_807) );
INVxp67_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g809 ( .A(n_810), .B(n_813), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OR2x2_ASAP7_75t_SL g831 ( .A(n_811), .B(n_813), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_811), .A2(n_836), .B(n_839), .Y(n_835) );
INVx1_ASAP7_75t_SL g826 ( .A(n_814), .Y(n_826) );
BUFx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx2_ASAP7_75t_R g828 ( .A(n_815), .Y(n_828) );
BUFx2_ASAP7_75t_L g840 ( .A(n_815), .Y(n_840) );
INVxp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AOI21xp33_ASAP7_75t_SL g817 ( .A1(n_818), .A2(n_825), .B(n_827), .Y(n_817) );
INVx1_ASAP7_75t_L g823 ( .A(n_820), .Y(n_823) );
INVx1_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_SL g827 ( .A(n_828), .B(n_829), .Y(n_827) );
CKINVDCx9p33_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_SL g834 ( .A(n_835), .Y(n_834) );
CKINVDCx11_ASAP7_75t_R g836 ( .A(n_837), .Y(n_836) );
CKINVDCx8_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
endmodule