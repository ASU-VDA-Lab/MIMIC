module fake_ariane_2622_n_1765 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1765);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1765;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx10_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_52),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_37),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_36),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_16),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_60),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_62),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_111),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_8),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_59),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_47),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_55),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_105),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_98),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_51),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_90),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_32),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_33),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_39),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_31),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_40),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_77),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_14),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_125),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_71),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_28),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_11),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_91),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_15),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_69),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_154),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_78),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_136),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_38),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_89),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_137),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_19),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_19),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_124),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_129),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_99),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_114),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_43),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_1),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_155),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_102),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_108),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_5),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_104),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_33),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_97),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_61),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_74),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_31),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_65),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_51),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_46),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_66),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_83),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_53),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_12),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_86),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_35),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_18),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_147),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_48),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_2),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_95),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_45),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_75),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_140),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_151),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_27),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_110),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_122),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_88),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_54),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_42),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_0),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_117),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_50),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_58),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_134),
.Y(n_269)
);

BUFx8_ASAP7_75t_SL g270 ( 
.A(n_17),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_24),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_34),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_120),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_73),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_25),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_79),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_93),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_72),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_3),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_121),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_27),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_29),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_100),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_25),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_48),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_26),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_142),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_135),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_109),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_30),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_46),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_21),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_112),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_26),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_64),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_40),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_4),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_92),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_38),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_44),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_20),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_44),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_162),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_204),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_185),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_270),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_226),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_185),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_185),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_156),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_185),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_185),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_185),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_162),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_185),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_164),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_156),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_231),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_204),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_231),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_231),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_231),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_231),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_231),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_164),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_159),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_160),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_263),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_263),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_249),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_263),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_263),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_186),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_165),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_192),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_211),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_198),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_200),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_209),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_213),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_165),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_177),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_177),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_170),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_190),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_190),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_238),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_238),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_179),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_179),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_211),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_181),
.B(n_1),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_197),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_220),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_197),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_156),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_300),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_217),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_183),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_170),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_184),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_249),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_245),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_196),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_218),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_203),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_227),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_171),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_349),
.A2(n_181),
.B1(n_274),
.B2(n_225),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_348),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_268),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_317),
.A2(n_176),
.B(n_168),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_313),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_220),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_189),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_310),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_335),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_322),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_362),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_319),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_320),
.A2(n_324),
.B(n_321),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_315),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_311),
.B(n_288),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_321),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_353),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_328),
.B(n_219),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_329),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_330),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_331),
.B(n_194),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_366),
.A2(n_206),
.B1(n_225),
.B2(n_195),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_318),
.B(n_245),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_333),
.B(n_215),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_342),
.B(n_288),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_366),
.A2(n_274),
.B1(n_206),
.B2(n_195),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_334),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_378),
.B(n_166),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_336),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_375),
.B(n_219),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_362),
.B(n_294),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_339),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_363),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_375),
.B(n_219),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_340),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_364),
.B(n_294),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_379),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_318),
.A2(n_259),
.B1(n_267),
.B2(n_171),
.Y(n_447)
);

BUFx8_ASAP7_75t_L g448 ( 
.A(n_326),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_337),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_340),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_341),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_364),
.B(n_166),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_341),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_414),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_408),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_387),
.B(n_326),
.Y(n_458)
);

OAI22x1_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_368),
.B1(n_265),
.B2(n_182),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

AND2x6_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_223),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_409),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_413),
.A2(n_376),
.B1(n_259),
.B2(n_267),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_387),
.B(n_370),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_391),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_438),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_409),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_417),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_SL g472 ( 
.A(n_449),
.B(n_338),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_387),
.B(n_438),
.Y(n_474)
);

BUFx6f_ASAP7_75t_SL g475 ( 
.A(n_413),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_370),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_405),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_443),
.B(n_345),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_417),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_425),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_382),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_435),
.B(n_347),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_419),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_421),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_400),
.B(n_350),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_394),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_433),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_435),
.B(n_351),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_400),
.B(n_352),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_434),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_434),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_418),
.B(n_371),
.Y(n_504)
);

AND3x2_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_239),
.C(n_234),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_413),
.B(n_430),
.Y(n_506)
);

NOR2x1p5_ASAP7_75t_L g507 ( 
.A(n_395),
.B(n_374),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_412),
.B(n_381),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_418),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_434),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_440),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_440),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_413),
.A2(n_307),
.B1(n_247),
.B2(n_261),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_442),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_418),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_L g518 ( 
.A1(n_386),
.A2(n_282),
.B1(n_306),
.B2(n_308),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_453),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_397),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_425),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_385),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_412),
.B(n_377),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_413),
.B(n_343),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_385),
.B(n_344),
.C(n_343),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_430),
.A2(n_284),
.B1(n_279),
.B2(n_272),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_397),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_420),
.B(n_367),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_425),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_401),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_447),
.A2(n_306),
.B1(n_308),
.B2(n_243),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_430),
.B(n_169),
.Y(n_540)
);

BUFx6f_ASAP7_75t_SL g541 ( 
.A(n_430),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_420),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_430),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_420),
.B(n_367),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_389),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_452),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_397),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_398),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_411),
.Y(n_549)
);

OA22x2_ASAP7_75t_L g550 ( 
.A1(n_407),
.A2(n_360),
.B1(n_346),
.B2(n_354),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_401),
.Y(n_551)
);

INVx8_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_392),
.B(n_169),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_403),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_398),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_452),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_452),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_404),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_398),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_404),
.B(n_344),
.C(n_369),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_410),
.B(n_372),
.C(n_369),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_396),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_420),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_452),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_398),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_392),
.B(n_172),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_398),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_451),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_451),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_407),
.B(n_372),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_406),
.Y(n_572)
);

CKINVDCx6p67_ASAP7_75t_R g573 ( 
.A(n_389),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_406),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_410),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_415),
.B(n_373),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_388),
.B(n_373),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_411),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_415),
.B(n_377),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_406),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_392),
.B(n_172),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_406),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_406),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_426),
.Y(n_584)
);

OAI22xp33_ASAP7_75t_L g585 ( 
.A1(n_432),
.A2(n_277),
.B1(n_236),
.B2(n_246),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_392),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_396),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_392),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_451),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_451),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_426),
.B(n_380),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_388),
.B(n_173),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_451),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_427),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_450),
.B(n_380),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_446),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_396),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_448),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_427),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_396),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_439),
.B(n_383),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_431),
.B(n_383),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_448),
.B(n_173),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_552),
.B(n_431),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_546),
.A2(n_428),
.B1(n_450),
.B2(n_436),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_543),
.A2(n_428),
.B1(n_447),
.B2(n_448),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_460),
.Y(n_607)
);

INVx4_ASAP7_75t_SL g608 ( 
.A(n_461),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_543),
.B(n_436),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_506),
.B(n_437),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_552),
.B(n_437),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_484),
.A2(n_445),
.B1(n_439),
.B2(n_448),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_530),
.B(n_598),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_526),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_521),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_506),
.B(n_444),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_469),
.B(n_444),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_469),
.B(n_422),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_509),
.B(n_422),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_509),
.B(n_429),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_516),
.B(n_429),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_526),
.B(n_423),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_516),
.B(n_448),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_393),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_524),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_571),
.B(n_393),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_474),
.B(n_439),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_466),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_488),
.B(n_489),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_482),
.B(n_396),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_524),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_460),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_525),
.A2(n_390),
.B(n_439),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_482),
.B(n_390),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_504),
.B(n_439),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_477),
.A2(n_390),
.B(n_445),
.C(n_271),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_550),
.A2(n_445),
.B1(n_423),
.B2(n_216),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_454),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_488),
.B(n_445),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_482),
.B(n_486),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_499),
.B(n_445),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_527),
.A2(n_564),
.B(n_542),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_546),
.B(n_174),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_557),
.B(n_558),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_482),
.B(n_174),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_529),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_529),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_478),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_537),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_458),
.B(n_250),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_552),
.Y(n_651)
);

AO221x1_ASAP7_75t_L g652 ( 
.A1(n_518),
.A2(n_187),
.B1(n_207),
.B2(n_237),
.C(n_241),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_461),
.A2(n_475),
.B1(n_541),
.B2(n_557),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_478),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_558),
.B(n_175),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_486),
.B(n_175),
.Y(n_656)
);

AND2x6_ASAP7_75t_SL g657 ( 
.A(n_495),
.B(n_394),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_565),
.B(n_252),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_483),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_537),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_486),
.B(n_216),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_565),
.B(n_256),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_464),
.B(n_266),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_461),
.B(n_586),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_466),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_486),
.B(n_242),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_530),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_483),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_461),
.B(n_273),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_501),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_502),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_461),
.B(n_285),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_502),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_550),
.A2(n_461),
.B1(n_541),
.B2(n_475),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_454),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_502),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_536),
.B(n_244),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_461),
.B(n_287),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_586),
.B(n_290),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_552),
.B(n_178),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_510),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_SL g682 ( 
.A1(n_463),
.A2(n_441),
.B1(n_416),
.B2(n_402),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_588),
.B(n_595),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_588),
.B(n_291),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_530),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_510),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_536),
.B(n_248),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_531),
.B(n_292),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_550),
.A2(n_475),
.B1(n_541),
.B2(n_585),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_530),
.A2(n_301),
.B1(n_297),
.B2(n_298),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_480),
.B(n_299),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_601),
.B(n_303),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_536),
.B(n_251),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_552),
.A2(n_255),
.B1(n_258),
.B2(n_264),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_538),
.A2(n_346),
.B(n_361),
.C(n_360),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_536),
.B(n_269),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_601),
.B(n_304),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_545),
.B(n_399),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_598),
.B(n_354),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_535),
.B(n_309),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_539),
.B(n_283),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_544),
.B(n_157),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_573),
.B(n_399),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_573),
.B(n_402),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_569),
.B(n_161),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_569),
.B(n_163),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_569),
.B(n_570),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_569),
.B(n_167),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_527),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_570),
.B(n_527),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_459),
.A2(n_228),
.B1(n_260),
.B2(n_223),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_551),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_553),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_553),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_540),
.B(n_289),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_570),
.B(n_180),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_596),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_539),
.B(n_293),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_527),
.B(n_188),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_473),
.B(n_355),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_555),
.A2(n_355),
.B(n_356),
.C(n_358),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_539),
.B(n_178),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_562),
.B(n_356),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_454),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_510),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_512),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_538),
.A2(n_579),
.B1(n_602),
.B2(n_591),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_592),
.B(n_2),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_539),
.B(n_6),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_542),
.B(n_191),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_505),
.B(n_358),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_520),
.B(n_178),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_512),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_512),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_542),
.B(n_193),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_508),
.B(n_416),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_507),
.B(n_359),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_542),
.B(n_199),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_555),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_564),
.B(n_201),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_559),
.A2(n_295),
.B1(n_221),
.B2(n_214),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_603),
.A2(n_240),
.B1(n_205),
.B2(n_208),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_564),
.B(n_202),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_559),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_472),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_520),
.B(n_178),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_513),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_575),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_564),
.B(n_212),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_575),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_507),
.B(n_441),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_584),
.B(n_222),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_584),
.B(n_467),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_520),
.Y(n_756)
);

AND2x6_ASAP7_75t_SL g757 ( 
.A(n_468),
.B(n_496),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_549),
.A2(n_257),
.B1(n_224),
.B2(n_305),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_467),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_594),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_513),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_459),
.A2(n_228),
.B1(n_260),
.B2(n_361),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_594),
.A2(n_359),
.B(n_7),
.C(n_9),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_554),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_599),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_467),
.B(n_302),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_599),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_467),
.B(n_296),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_514),
.A2(n_187),
.B1(n_207),
.B2(n_178),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_476),
.B(n_281),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_549),
.B(n_178),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_476),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_576),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_476),
.B(n_280),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_700),
.Y(n_775)
);

BUFx8_ASAP7_75t_L g776 ( 
.A(n_705),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_628),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_757),
.B(n_476),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_670),
.B(n_567),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_615),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_651),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_628),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_671),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_614),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_637),
.A2(n_533),
.B1(n_562),
.B2(n_455),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_625),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_719),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_622),
.B(n_581),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_631),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_738),
.B(n_522),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_629),
.B(n_455),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_651),
.B(n_549),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_613),
.B(n_589),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_706),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_731),
.B(n_578),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_671),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_739),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_731),
.B(n_578),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_624),
.B(n_456),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_626),
.B(n_456),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_756),
.A2(n_578),
.B(n_600),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_729),
.B(n_589),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_635),
.B(n_619),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_682),
.B(n_522),
.Y(n_804)
);

NOR2x1p5_ASAP7_75t_L g805 ( 
.A(n_753),
.B(n_561),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_646),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_657),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_683),
.B(n_590),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_647),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_635),
.B(n_457),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_R g811 ( 
.A(n_680),
.B(n_457),
.Y(n_811)
);

AO22x1_ASAP7_75t_L g812 ( 
.A1(n_667),
.A2(n_462),
.B1(n_465),
.B2(n_470),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_620),
.B(n_462),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_621),
.B(n_465),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_686),
.A2(n_532),
.B1(n_470),
.B2(n_491),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_613),
.B(n_590),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_649),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_660),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_747),
.B(n_561),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_618),
.B(n_471),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_739),
.Y(n_821)
);

NAND2x1p5_ASAP7_75t_L g822 ( 
.A(n_726),
.B(n_597),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_773),
.B(n_471),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_664),
.B(n_593),
.Y(n_824)
);

OR2x2_ASAP7_75t_SL g825 ( 
.A(n_606),
.B(n_523),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_613),
.B(n_593),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_673),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_726),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_688),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_628),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_759),
.B(n_466),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_714),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_759),
.B(n_466),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_639),
.B(n_641),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_650),
.B(n_479),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_701),
.Y(n_836)
);

NOR2x2_ASAP7_75t_L g837 ( 
.A(n_692),
.B(n_572),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_650),
.A2(n_532),
.B1(n_479),
.B2(n_481),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_739),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_674),
.A2(n_652),
.B1(n_691),
.B2(n_717),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_772),
.B(n_466),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_701),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_772),
.B(n_492),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_608),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_684),
.A2(n_500),
.B1(n_494),
.B2(n_481),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_717),
.A2(n_485),
.B1(n_515),
.B2(n_511),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_701),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_673),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_715),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_733),
.Y(n_850)
);

INVx5_ASAP7_75t_L g851 ( 
.A(n_628),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_663),
.A2(n_500),
.B1(n_511),
.B2(n_485),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_733),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_663),
.B(n_491),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_722),
.B(n_494),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_730),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_716),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_694),
.B(n_515),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_610),
.B(n_519),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_638),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_676),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_676),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_608),
.B(n_523),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_665),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_608),
.B(n_764),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_681),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_681),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_733),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_693),
.Y(n_869)
);

CKINVDCx6p67_ASAP7_75t_R g870 ( 
.A(n_623),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_693),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_687),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_665),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_653),
.B(n_597),
.Y(n_874)
);

BUFx6f_ASAP7_75t_SL g875 ( 
.A(n_741),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_746),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_616),
.B(n_519),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_699),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_730),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_605),
.B(n_528),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_750),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_687),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_644),
.B(n_492),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_752),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_638),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_696),
.A2(n_572),
.B1(n_574),
.B2(n_580),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_675),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_760),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_675),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_665),
.B(n_492),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_609),
.A2(n_572),
.B1(n_574),
.B2(n_580),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_SL g892 ( 
.A1(n_680),
.A2(n_498),
.B1(n_487),
.B2(n_490),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_627),
.B(n_528),
.Y(n_893)
);

CKINVDCx14_ASAP7_75t_R g894 ( 
.A(n_758),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_702),
.B(n_534),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_697),
.A2(n_513),
.B(n_487),
.C(n_498),
.Y(n_896)
);

AND3x1_ASAP7_75t_SL g897 ( 
.A(n_765),
.B(n_6),
.C(n_9),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_727),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_727),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_744),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_697),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_665),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_612),
.A2(n_574),
.B1(n_580),
.B2(n_582),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_640),
.B(n_492),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_767),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_679),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_728),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_658),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_R g909 ( 
.A(n_604),
.B(n_600),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_728),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_617),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_735),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_642),
.A2(n_493),
.B(n_490),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_690),
.B(n_597),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_735),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_736),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_662),
.B(n_534),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_736),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_SL g919 ( 
.A1(n_669),
.A2(n_493),
.B1(n_497),
.B2(n_503),
.Y(n_919)
);

INVx5_ASAP7_75t_L g920 ( 
.A(n_749),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_749),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_761),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_640),
.B(n_492),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_761),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_725),
.B(n_685),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_709),
.B(n_547),
.Y(n_926)
);

INVxp67_ASAP7_75t_SL g927 ( 
.A(n_611),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_607),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_643),
.B(n_547),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_630),
.B(n_636),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_754),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_762),
.B(n_497),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_704),
.B(n_548),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_607),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_632),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_655),
.B(n_548),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_711),
.B(n_563),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_712),
.A2(n_600),
.B(n_597),
.Y(n_938)
);

BUFx4f_ASAP7_75t_L g939 ( 
.A(n_632),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_755),
.B(n_556),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_666),
.A2(n_582),
.B1(n_556),
.B2(n_583),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_648),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_648),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_654),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_666),
.B(n_600),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_677),
.B(n_560),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_L g947 ( 
.A(n_743),
.B(n_560),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_672),
.B(n_563),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_636),
.B(n_566),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_654),
.B(n_659),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_677),
.B(n_566),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_633),
.B(n_563),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_659),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_668),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_668),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_713),
.B(n_568),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_689),
.A2(n_582),
.B1(n_583),
.B2(n_568),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_689),
.B(n_517),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_695),
.B(n_698),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_695),
.B(n_517),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_769),
.A2(n_503),
.B1(n_563),
.B2(n_587),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_698),
.B(n_587),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_SL g963 ( 
.A1(n_678),
.A2(n_235),
.B1(n_276),
.B2(n_229),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_634),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_795),
.A2(n_634),
.B(n_771),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_795),
.A2(n_734),
.B(n_771),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_803),
.A2(n_645),
.B1(n_656),
.B2(n_703),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_SL g968 ( 
.A(n_869),
.B(n_645),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_856),
.A2(n_720),
.B(n_703),
.C(n_763),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_911),
.B(n_720),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_879),
.A2(n_656),
.B1(n_661),
.B2(n_708),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_871),
.B(n_707),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_788),
.B(n_821),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_784),
.B(n_710),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_781),
.B(n_721),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_779),
.A2(n_723),
.B(n_661),
.C(n_718),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_834),
.B(n_630),
.Y(n_977)
);

OAI22x1_ASAP7_75t_L g978 ( 
.A1(n_900),
.A2(n_734),
.B1(n_748),
.B2(n_724),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_777),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_781),
.B(n_732),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_779),
.B(n_766),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_878),
.A2(n_835),
.B(n_854),
.C(n_802),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_836),
.B(n_737),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_787),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_775),
.B(n_11),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_781),
.B(n_740),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_836),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_842),
.B(n_745),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_780),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_801),
.A2(n_748),
.B(n_724),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_781),
.B(n_751),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_802),
.A2(n_742),
.B(n_770),
.C(n_768),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_847),
.B(n_774),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_794),
.B(n_12),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_797),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_799),
.B(n_587),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_839),
.B(n_587),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_798),
.A2(n_587),
.B(n_563),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_894),
.A2(n_278),
.B1(n_275),
.B2(n_262),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_793),
.B(n_254),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_798),
.A2(n_253),
.B(n_233),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_800),
.B(n_13),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_810),
.A2(n_232),
.B(n_230),
.Y(n_1003)
);

NAND2x1p5_ASAP7_75t_L g1004 ( 
.A(n_844),
.B(n_207),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_944),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_894),
.B(n_13),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_SL g1007 ( 
.A1(n_807),
.A2(n_207),
.B1(n_187),
.B2(n_178),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_931),
.B(n_16),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_927),
.A2(n_207),
.B(n_187),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_850),
.B(n_17),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_927),
.A2(n_952),
.B(n_877),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_791),
.B(n_18),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_790),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_844),
.B(n_853),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_804),
.B(n_20),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_858),
.B(n_21),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_906),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1017)
);

O2A1O1Ixp5_ASAP7_75t_L g1018 ( 
.A1(n_952),
.A2(n_792),
.B(n_914),
.C(n_904),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_944),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_859),
.A2(n_187),
.B1(n_29),
.B2(n_30),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_786),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_819),
.A2(n_22),
.B(n_32),
.C(n_35),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_793),
.B(n_37),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_908),
.B(n_41),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_823),
.A2(n_41),
.B(n_42),
.C(n_49),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_901),
.B(n_789),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_955),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_806),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_809),
.B(n_49),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_813),
.A2(n_814),
.B(n_820),
.C(n_959),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_777),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_868),
.B(n_50),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_955),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_964),
.A2(n_56),
.B(n_57),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_805),
.A2(n_63),
.B1(n_68),
.B2(n_70),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_817),
.B(n_76),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_SL g1037 ( 
.A1(n_937),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_SL g1038 ( 
.A1(n_792),
.A2(n_85),
.B(n_87),
.C(n_94),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_964),
.A2(n_96),
.B(n_106),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_818),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_829),
.B(n_113),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_832),
.A2(n_857),
.B1(n_849),
.B2(n_884),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_796),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_937),
.A2(n_115),
.B(n_116),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_870),
.B(n_118),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_876),
.A2(n_119),
.B(n_123),
.C(n_143),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_881),
.B(n_149),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_776),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_816),
.B(n_153),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_888),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_875),
.B(n_825),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_872),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_816),
.B(n_826),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_785),
.B(n_840),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_933),
.A2(n_914),
.B(n_895),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_826),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_SL g1057 ( 
.A(n_939),
.B(n_875),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_845),
.A2(n_938),
.B(n_883),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_840),
.B(n_846),
.C(n_852),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_872),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_828),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_777),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_785),
.B(n_808),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_905),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_917),
.A2(n_936),
.B(n_893),
.C(n_889),
.Y(n_1065)
);

AND3x1_ASAP7_75t_L g1066 ( 
.A(n_778),
.B(n_808),
.C(n_776),
.Y(n_1066)
);

AOI22x1_ASAP7_75t_L g1067 ( 
.A1(n_885),
.A2(n_889),
.B1(n_887),
.B2(n_860),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_865),
.B(n_932),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_882),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_882),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_865),
.B(n_828),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_939),
.Y(n_1072)
);

BUFx2_ASAP7_75t_R g1073 ( 
.A(n_830),
.Y(n_1073)
);

BUFx8_ASAP7_75t_L g1074 ( 
.A(n_778),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_SL g1075 ( 
.A1(n_945),
.A2(n_860),
.B(n_887),
.C(n_951),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_940),
.A2(n_890),
.B(n_913),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_777),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_R g1078 ( 
.A(n_851),
.B(n_925),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_L g1079 ( 
.A(n_925),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_880),
.A2(n_846),
.B1(n_930),
.B2(n_838),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_890),
.A2(n_923),
.B(n_904),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_930),
.B(n_910),
.Y(n_1082)
);

OAI22x1_ASAP7_75t_L g1083 ( 
.A1(n_837),
.A2(n_815),
.B1(n_897),
.B2(n_903),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_934),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_910),
.B(n_916),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_960),
.A2(n_945),
.B(n_946),
.C(n_951),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_916),
.B(n_924),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_960),
.A2(n_946),
.B(n_947),
.C(n_929),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_783),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_830),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_885),
.A2(n_923),
.B(n_891),
.C(n_843),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_864),
.Y(n_1092)
);

AO32x1_ASAP7_75t_L g1093 ( 
.A1(n_941),
.A2(n_957),
.A3(n_897),
.B1(n_954),
.B2(n_953),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_855),
.A2(n_896),
.B(n_949),
.C(n_962),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_831),
.A2(n_843),
.B(n_841),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_942),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_831),
.A2(n_833),
.B(n_841),
.C(n_896),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_812),
.B(n_924),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_851),
.B(n_902),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_833),
.A2(n_824),
.B(n_958),
.C(n_926),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_864),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_918),
.B(n_921),
.Y(n_1102)
);

BUFx4f_ASAP7_75t_L g1103 ( 
.A(n_782),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_886),
.A2(n_892),
.B1(n_961),
.B2(n_956),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_961),
.A2(n_851),
.B1(n_920),
.B2(n_874),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_873),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_824),
.A2(n_926),
.B(n_822),
.C(n_922),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_782),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_928),
.A2(n_935),
.B(n_863),
.C(n_873),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_950),
.A2(n_822),
.B(n_920),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_963),
.A2(n_863),
.B1(n_902),
.B2(n_907),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_851),
.B(n_920),
.Y(n_1112)
);

AO32x1_ASAP7_75t_L g1113 ( 
.A1(n_943),
.A2(n_899),
.A3(n_912),
.B1(n_827),
.B2(n_848),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_811),
.B(n_920),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_1080),
.B(n_874),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_990),
.A2(n_867),
.B(n_898),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_978),
.A2(n_861),
.A3(n_862),
.B(n_866),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1013),
.B(n_935),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1014),
.B(n_782),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_972),
.B(n_782),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1076),
.A2(n_915),
.B(n_928),
.Y(n_1121)
);

OA21x2_ASAP7_75t_L g1122 ( 
.A1(n_1018),
.A2(n_919),
.B(n_811),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_981),
.A2(n_907),
.B(n_909),
.C(n_948),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1086),
.A2(n_909),
.B(n_948),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_1080),
.A2(n_907),
.B(n_967),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_984),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1055),
.A2(n_907),
.B(n_1058),
.Y(n_1127)
);

AOI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_1054),
.A2(n_1059),
.B(n_1083),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1011),
.A2(n_965),
.B(n_998),
.Y(n_1129)
);

O2A1O1Ixp5_ASAP7_75t_L g1130 ( 
.A1(n_968),
.A2(n_971),
.B(n_967),
.C(n_991),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_1099),
.B(n_1103),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1026),
.B(n_987),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1014),
.B(n_1053),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1108),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_L g1135 ( 
.A(n_977),
.B(n_1067),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_989),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_1014),
.B(n_1071),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_982),
.A2(n_1030),
.B(n_1065),
.C(n_1008),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1072),
.B(n_1056),
.Y(n_1139)
);

NAND2x1p5_ASAP7_75t_L g1140 ( 
.A(n_1099),
.B(n_1103),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_1082),
.Y(n_1141)
);

BUFx4_ASAP7_75t_SL g1142 ( 
.A(n_1048),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1020),
.A2(n_1015),
.B(n_1006),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_1068),
.B(n_1114),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_971),
.A2(n_1063),
.B(n_1002),
.C(n_1016),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1073),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_966),
.A2(n_1081),
.B(n_1095),
.Y(n_1147)
);

AO21x1_ASAP7_75t_L g1148 ( 
.A1(n_1020),
.A2(n_1104),
.B(n_1098),
.Y(n_1148)
);

OAI22x1_ASAP7_75t_L g1149 ( 
.A1(n_1051),
.A2(n_999),
.B1(n_1035),
.B2(n_1010),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1061),
.B(n_1021),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1012),
.A2(n_969),
.B(n_976),
.C(n_1088),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_1074),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1010),
.A2(n_1023),
.B1(n_1000),
.B2(n_1032),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1077),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_1072),
.B(n_1077),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1090),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1061),
.B(n_1028),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_L g1158 ( 
.A1(n_1104),
.A2(n_1025),
.B(n_1075),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1024),
.B(n_1040),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1057),
.B(n_985),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1097),
.A2(n_1037),
.B(n_1110),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_977),
.B(n_1082),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1094),
.A2(n_1009),
.B(n_996),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1105),
.A2(n_1085),
.A3(n_1109),
.B(n_1027),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_992),
.A2(n_1105),
.B(n_1091),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1107),
.A2(n_1100),
.B(n_1044),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_975),
.A2(n_980),
.B(n_986),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1034),
.A2(n_1039),
.B(n_1004),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1042),
.B(n_995),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1012),
.A2(n_970),
.B(n_1047),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1085),
.A2(n_1033),
.A3(n_1019),
.B(n_1005),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_1077),
.B(n_1101),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1043),
.A2(n_1052),
.A3(n_1070),
.B(n_1069),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_983),
.A2(n_1029),
.B(n_1036),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1092),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_997),
.A2(n_1087),
.B(n_1102),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1004),
.A2(n_1087),
.B(n_1112),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_1077),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1112),
.A2(n_1041),
.B(n_1046),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1042),
.A2(n_1093),
.B(n_1038),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1057),
.B(n_1079),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1022),
.A2(n_1017),
.B(n_988),
.C(n_993),
.Y(n_1182)
);

AO32x2_ASAP7_75t_L g1183 ( 
.A1(n_1093),
.A2(n_1113),
.A3(n_1084),
.B1(n_1096),
.B2(n_1066),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1093),
.A2(n_1049),
.B(n_1003),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1060),
.A2(n_1111),
.B(n_1064),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_1078),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1106),
.B(n_1050),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_L g1188 ( 
.A(n_994),
.B(n_1007),
.C(n_1045),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_L g1189 ( 
.A(n_979),
.B(n_1031),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1106),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1001),
.A2(n_1079),
.B(n_1031),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_979),
.B(n_1031),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1074),
.B(n_979),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1062),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1062),
.B(n_1113),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1062),
.A2(n_981),
.B(n_856),
.C(n_1059),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_1113),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_989),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1013),
.B(n_670),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1103),
.Y(n_1200)
);

INVx6_ASAP7_75t_L g1201 ( 
.A(n_1074),
.Y(n_1201)
);

NAND2x1_ASAP7_75t_SL g1202 ( 
.A(n_1045),
.B(n_753),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1013),
.B(n_670),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1013),
.B(n_670),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_972),
.B(n_869),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1089),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_981),
.B(n_879),
.C(n_871),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1086),
.A2(n_967),
.B(n_965),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1080),
.A2(n_879),
.B1(n_871),
.B2(n_869),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1013),
.B(n_670),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_973),
.B(n_622),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1055),
.A2(n_756),
.B(n_795),
.Y(n_1215)
);

AO21x2_ASAP7_75t_L g1216 ( 
.A1(n_1055),
.A2(n_965),
.B(n_966),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_SL g1217 ( 
.A1(n_981),
.A2(n_538),
.B(n_670),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1013),
.B(n_670),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1055),
.A2(n_756),
.B(n_795),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_1055),
.A2(n_965),
.B(n_966),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1086),
.A2(n_967),
.B(n_965),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1013),
.B(n_670),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_978),
.A2(n_1055),
.A3(n_1104),
.B(n_1094),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1074),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1014),
.B(n_1053),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1014),
.B(n_1053),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1080),
.A2(n_879),
.B1(n_871),
.B2(n_869),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_972),
.A2(n_981),
.B(n_779),
.C(n_974),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_973),
.B(n_622),
.Y(n_1234)
);

O2A1O1Ixp5_ASAP7_75t_L g1235 ( 
.A1(n_968),
.A2(n_795),
.B(n_798),
.C(n_1058),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_978),
.A2(n_1055),
.A3(n_1104),
.B(n_1094),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_989),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1055),
.A2(n_756),
.B(n_795),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1073),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_989),
.Y(n_1242)
);

O2A1O1Ixp5_ASAP7_75t_SL g1243 ( 
.A1(n_1020),
.A2(n_952),
.B(n_364),
.C(n_367),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_981),
.B(n_879),
.C(n_871),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1086),
.A2(n_967),
.B(n_965),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1013),
.B(n_670),
.Y(n_1246)
);

NOR4xp25_ASAP7_75t_L g1247 ( 
.A(n_1020),
.B(n_1025),
.C(n_1022),
.D(n_1017),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1013),
.B(n_670),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1013),
.B(n_670),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_989),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1013),
.B(n_670),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_990),
.A2(n_1076),
.B(n_1058),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_973),
.B(n_622),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1086),
.A2(n_967),
.B(n_965),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1055),
.A2(n_756),
.B(n_795),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1063),
.B(n_1054),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_973),
.B(n_622),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1055),
.A2(n_756),
.B(n_795),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_973),
.B(n_622),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_973),
.B(n_622),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1080),
.A2(n_879),
.B1(n_803),
.B2(n_856),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1180),
.A2(n_1165),
.B(n_1158),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1171),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1210),
.B(n_1222),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1217),
.B(n_1261),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1261),
.A2(n_1188),
.B1(n_1148),
.B2(n_1128),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1221),
.A2(n_1227),
.B(n_1223),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1212),
.A2(n_1231),
.B1(n_1217),
.B2(n_1209),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1128),
.A2(n_1115),
.B1(n_1260),
.B2(n_1259),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1119),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_1257),
.B1(n_1214),
.B2(n_1253),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1229),
.A2(n_1239),
.B(n_1252),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1198),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1231),
.A2(n_1244),
.B1(n_1209),
.B2(n_1143),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1142),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1119),
.B(n_1133),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1244),
.B(n_1143),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1171),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1184),
.A2(n_1158),
.B(n_1170),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1126),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1145),
.A2(n_1151),
.B(n_1138),
.C(n_1130),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1238),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1206),
.B(n_1196),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1134),
.Y(n_1285)
);

BUFx4f_ASAP7_75t_L g1286 ( 
.A(n_1131),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1242),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1233),
.A2(n_1237),
.B(n_1129),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1175),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1127),
.A2(n_1258),
.B(n_1215),
.Y(n_1290)
);

AOI31xp67_ASAP7_75t_L g1291 ( 
.A1(n_1195),
.A2(n_1162),
.A3(n_1256),
.B(n_1192),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1234),
.A2(n_1125),
.B1(n_1149),
.B2(n_1153),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1147),
.A2(n_1161),
.B(n_1168),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1160),
.A2(n_1256),
.B1(n_1174),
.B2(n_1207),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1250),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1199),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1219),
.A2(n_1255),
.B(n_1240),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1116),
.A2(n_1121),
.B(n_1254),
.Y(n_1298)
);

AND2x6_ASAP7_75t_L g1299 ( 
.A(n_1133),
.B(n_1228),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1245),
.A2(n_1254),
.B(n_1166),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1245),
.A2(n_1124),
.B(n_1182),
.C(n_1235),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1179),
.A2(n_1177),
.B(n_1243),
.Y(n_1302)
);

AO21x2_ASAP7_75t_L g1303 ( 
.A1(n_1197),
.A2(n_1124),
.B(n_1185),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1163),
.A2(n_1176),
.B(n_1167),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1163),
.A2(n_1191),
.B(n_1122),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1247),
.A2(n_1135),
.B(n_1123),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1150),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1183),
.B(n_1236),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1157),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_SL g1310 ( 
.A1(n_1132),
.A2(n_1178),
.B(n_1118),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1122),
.A2(n_1146),
.B1(n_1241),
.B2(n_1230),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1216),
.A2(n_1220),
.B(n_1120),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1194),
.A2(n_1141),
.B(n_1190),
.Y(n_1313)
);

BUFx8_ASAP7_75t_L g1314 ( 
.A(n_1226),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1216),
.A2(n_1220),
.B(n_1189),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1194),
.A2(n_1181),
.B(n_1172),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1131),
.A2(n_1140),
.B(n_1202),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_SL g1318 ( 
.A1(n_1178),
.A2(n_1159),
.B(n_1249),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1187),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1140),
.A2(n_1155),
.B(n_1200),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1183),
.B(n_1225),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1187),
.B(n_1203),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1192),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1247),
.A2(n_1204),
.B(n_1224),
.C(n_1218),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1213),
.B(n_1251),
.C(n_1248),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1183),
.B(n_1236),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1146),
.A2(n_1241),
.B1(n_1228),
.B2(n_1230),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1173),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1154),
.Y(n_1329)
);

NAND3xp33_ASAP7_75t_L g1330 ( 
.A(n_1246),
.B(n_1144),
.C(n_1193),
.Y(n_1330)
);

AOI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1139),
.A2(n_1186),
.B1(n_1152),
.B2(n_1236),
.C(n_1225),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1225),
.B(n_1117),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1117),
.A2(n_1164),
.A3(n_1137),
.B(n_1154),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1117),
.A2(n_1164),
.B(n_1154),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1164),
.A2(n_670),
.B(n_1217),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1201),
.B(n_1169),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1201),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1171),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1217),
.B(n_1261),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1217),
.B(n_1261),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1342)
);

AO21x1_ASAP7_75t_L g1343 ( 
.A1(n_1261),
.A2(n_1143),
.B(n_1080),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1151),
.A2(n_1222),
.B(n_1210),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1171),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1142),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1154),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1261),
.A2(n_682),
.B1(n_423),
.B2(n_484),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1136),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1119),
.B(n_1133),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1171),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1156),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1136),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1181),
.B(n_1077),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1171),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1180),
.A2(n_1184),
.B(n_1158),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1154),
.Y(n_1359)
);

CKINVDCx6p67_ASAP7_75t_R g1360 ( 
.A(n_1152),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1217),
.B(n_1232),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1171),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1151),
.A2(n_1222),
.B(n_1210),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1180),
.A2(n_1184),
.B(n_1158),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1217),
.B(n_1261),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1126),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1171),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1210),
.B(n_1222),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1261),
.A2(n_322),
.B1(n_325),
.B2(n_310),
.Y(n_1372)
);

AOI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1217),
.A2(n_518),
.B1(n_386),
.B2(n_463),
.C(n_1261),
.Y(n_1373)
);

CKINVDCx8_ASAP7_75t_R g1374 ( 
.A(n_1156),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1156),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1142),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_SL g1379 ( 
.A(n_1212),
.B(n_879),
.C(n_871),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1119),
.B(n_1133),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1210),
.B(n_1222),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1119),
.B(n_1133),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1212),
.A2(n_1231),
.B1(n_1217),
.B2(n_879),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1208),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1344),
.A2(n_1364),
.B(n_1282),
.Y(n_1389)
);

AO21x1_ASAP7_75t_L g1390 ( 
.A1(n_1266),
.A2(n_1341),
.B(n_1340),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1266),
.A2(n_1367),
.B1(n_1341),
.B2(n_1340),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1276),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1313),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1278),
.B(n_1322),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1276),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1368),
.B(n_1281),
.Y(n_1396)
);

AOI211xp5_ASAP7_75t_L g1397 ( 
.A1(n_1269),
.A2(n_1367),
.B(n_1384),
.C(n_1275),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1293),
.A2(n_1300),
.B(n_1315),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1289),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1361),
.A2(n_1373),
.B(n_1278),
.C(n_1379),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1293),
.A2(n_1300),
.B(n_1305),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1343),
.A2(n_1306),
.B(n_1301),
.C(n_1336),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1264),
.A2(n_1382),
.B(n_1371),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1337),
.B(n_1354),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1264),
.A2(n_1371),
.B1(n_1382),
.B2(n_1267),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1330),
.B(n_1325),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1274),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1354),
.B(n_1375),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1294),
.B(n_1307),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1350),
.A2(n_1301),
.B1(n_1284),
.B2(n_1270),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_SL g1411 ( 
.A(n_1348),
.B(n_1377),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1319),
.B(n_1283),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1287),
.B(n_1295),
.Y(n_1413)
);

CKINVDCx14_ASAP7_75t_R g1414 ( 
.A(n_1348),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1308),
.A2(n_1326),
.B(n_1321),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1351),
.B(n_1355),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1272),
.B(n_1284),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1333),
.B(n_1323),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1331),
.A2(n_1324),
.B(n_1296),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1372),
.A2(n_1292),
.B1(n_1374),
.B2(n_1327),
.Y(n_1420)
);

NOR2xp67_ASAP7_75t_L g1421 ( 
.A(n_1338),
.B(n_1309),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1308),
.B(n_1277),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1374),
.A2(n_1311),
.B1(n_1285),
.B2(n_1286),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1305),
.A2(n_1286),
.B(n_1317),
.C(n_1312),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1285),
.A2(n_1286),
.B1(n_1377),
.B2(n_1360),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1318),
.A2(n_1310),
.B(n_1262),
.C(n_1358),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1262),
.B(n_1332),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1303),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1328),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1288),
.A2(n_1304),
.B(n_1369),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1262),
.B(n_1332),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1314),
.B(n_1329),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1280),
.B(n_1358),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1280),
.B(n_1366),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1356),
.A2(n_1383),
.B1(n_1381),
.B2(n_1352),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1381),
.A2(n_1271),
.B1(n_1329),
.B2(n_1359),
.Y(n_1436)
);

AOI221x1_ASAP7_75t_SL g1437 ( 
.A1(n_1314),
.A2(n_1366),
.B1(n_1291),
.B2(n_1339),
.C(n_1347),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1317),
.A2(n_1316),
.B(n_1320),
.C(n_1335),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1334),
.B(n_1349),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1349),
.A2(n_1359),
.B1(n_1370),
.B2(n_1363),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1334),
.B(n_1299),
.Y(n_1441)
);

AOI31xp33_ASAP7_75t_L g1442 ( 
.A1(n_1299),
.A2(n_1263),
.A3(n_1370),
.B(n_1357),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1290),
.A2(n_1388),
.B(n_1386),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1299),
.B(n_1335),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1299),
.B(n_1304),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1299),
.B(n_1298),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1290),
.A2(n_1388),
.B(n_1386),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1376),
.B(n_1388),
.Y(n_1448)
);

AND2x2_ASAP7_75t_SL g1449 ( 
.A(n_1279),
.B(n_1347),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1376),
.A2(n_1386),
.B(n_1357),
.C(n_1353),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1376),
.A2(n_1353),
.B(n_1339),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1288),
.A2(n_1265),
.B(n_1268),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1298),
.B(n_1297),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1302),
.B(n_1297),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1265),
.A2(n_1268),
.B1(n_1273),
.B2(n_1342),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1273),
.B(n_1342),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1345),
.A2(n_1346),
.B(n_1362),
.C(n_1365),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1345),
.A2(n_1346),
.B(n_1362),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_1369),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1378),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1461)
);

AOI221xp5_ASAP7_75t_L g1462 ( 
.A1(n_1385),
.A2(n_1373),
.B1(n_1217),
.B2(n_1261),
.C(n_518),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1387),
.Y(n_1463)
);

O2A1O1Ixp5_ASAP7_75t_L g1464 ( 
.A1(n_1387),
.A2(n_1148),
.B(n_1343),
.C(n_1344),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1278),
.B(n_1322),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1278),
.B(n_1322),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1266),
.A2(n_1340),
.B1(n_1367),
.B2(n_1341),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1266),
.A2(n_1340),
.B1(n_1367),
.B2(n_1341),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1266),
.A2(n_1340),
.B1(n_1367),
.B2(n_1341),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1384),
.A2(n_1232),
.B(n_1217),
.C(n_1269),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1264),
.B(n_1371),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1278),
.B(n_1322),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1384),
.A2(n_1232),
.B(n_1217),
.C(n_1269),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1471),
.B(n_1403),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1403),
.B(n_1471),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1428),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1429),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1445),
.B(n_1446),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1433),
.A2(n_1434),
.B(n_1443),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1427),
.Y(n_1480)
);

OAI21xp33_ASAP7_75t_L g1481 ( 
.A1(n_1391),
.A2(n_1469),
.B(n_1468),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1407),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1431),
.B(n_1459),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1463),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1413),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1416),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1447),
.A2(n_1451),
.B(n_1450),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_L g1488 ( 
.A(n_1426),
.B(n_1419),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1431),
.B(n_1448),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1439),
.Y(n_1490)
);

OR2x6_ASAP7_75t_L g1491 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1405),
.A2(n_1393),
.B(n_1457),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1412),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1391),
.B(n_1467),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1399),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1464),
.A2(n_1402),
.B(n_1460),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1409),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1422),
.B(n_1467),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1454),
.B(n_1468),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1456),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1410),
.A2(n_1390),
.B1(n_1420),
.B2(n_1469),
.Y(n_1502)
);

OAI21xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1389),
.A2(n_1462),
.B(n_1405),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1389),
.B(n_1472),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1394),
.B(n_1465),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1461),
.B(n_1466),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1396),
.B(n_1453),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1438),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1408),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1449),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1398),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1401),
.B(n_1404),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1440),
.A2(n_1424),
.B(n_1455),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1430),
.B(n_1452),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1437),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1476),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1477),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1502),
.A2(n_1397),
.B1(n_1410),
.B2(n_1462),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1502),
.A2(n_1420),
.B1(n_1417),
.B2(n_1406),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1501),
.B(n_1491),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1475),
.B(n_1458),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1481),
.A2(n_1503),
.B(n_1495),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1500),
.B(n_1440),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1476),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1500),
.B(n_1415),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1400),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1501),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1489),
.B(n_1473),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1484),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1474),
.B(n_1418),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1489),
.B(n_1474),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1503),
.A2(n_1423),
.B1(n_1421),
.B2(n_1435),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1489),
.B(n_1474),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1512),
.B(n_1442),
.Y(n_1535)
);

AO22x1_ASAP7_75t_L g1536 ( 
.A1(n_1488),
.A2(n_1423),
.B1(n_1435),
.B2(n_1436),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1527),
.B(n_1522),
.C(n_1518),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1516),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1522),
.A2(n_1511),
.B(n_1514),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1520),
.Y(n_1540)
);

OAI31xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1527),
.A2(n_1518),
.A3(n_1488),
.B(n_1529),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1532),
.B(n_1506),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1532),
.B(n_1506),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1519),
.A2(n_1495),
.B1(n_1515),
.B2(n_1504),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1519),
.A2(n_1470),
.B1(n_1499),
.B2(n_1504),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

OAI31xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1529),
.A2(n_1425),
.A3(n_1483),
.B(n_1508),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1536),
.A2(n_1487),
.B(n_1513),
.Y(n_1548)
);

AO21x1_ASAP7_75t_SL g1549 ( 
.A1(n_1533),
.A2(n_1499),
.B(n_1508),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_SL g1550 ( 
.A(n_1529),
.B(n_1515),
.C(n_1499),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1532),
.B(n_1480),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1517),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1535),
.A2(n_1505),
.B1(n_1491),
.B2(n_1492),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

OAI222xp33_ASAP7_75t_L g1555 ( 
.A1(n_1526),
.A2(n_1483),
.B1(n_1498),
.B2(n_1505),
.C1(n_1492),
.C2(n_1491),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1520),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1516),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1526),
.A2(n_1535),
.B1(n_1510),
.B2(n_1493),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1478),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_R g1560 ( 
.A(n_1526),
.B(n_1414),
.Y(n_1560)
);

AOI222xp33_ASAP7_75t_L g1561 ( 
.A1(n_1536),
.A2(n_1425),
.B1(n_1494),
.B2(n_1486),
.C1(n_1485),
.C2(n_1482),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1535),
.A2(n_1493),
.B1(n_1513),
.B2(n_1490),
.Y(n_1562)
);

OAI211xp5_ASAP7_75t_L g1563 ( 
.A1(n_1521),
.A2(n_1496),
.B(n_1511),
.C(n_1497),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1509),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1517),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1523),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1552),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1539),
.B(n_1521),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1539),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1538),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1552),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1539),
.Y(n_1575)
);

AND4x1_ASAP7_75t_L g1576 ( 
.A(n_1541),
.B(n_1411),
.C(n_1432),
.D(n_1524),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1540),
.B(n_1521),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1537),
.C(n_1544),
.Y(n_1578)
);

INVx4_ASAP7_75t_SL g1579 ( 
.A(n_1546),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1554),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1549),
.Y(n_1581)
);

INVx4_ASAP7_75t_SL g1582 ( 
.A(n_1546),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1554),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1565),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1551),
.B(n_1525),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1547),
.B(n_1530),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1549),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1557),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1537),
.Y(n_1589)
);

AO21x2_ASAP7_75t_L g1590 ( 
.A1(n_1548),
.A2(n_1487),
.B(n_1479),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1544),
.B(n_1524),
.C(n_1496),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1572),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1589),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1568),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1587),
.B(n_1542),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1571),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1568),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1587),
.B(n_1581),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1573),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1578),
.A2(n_1545),
.B1(n_1550),
.B2(n_1561),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1589),
.B(n_1392),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1581),
.B(n_1542),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1579),
.B(n_1556),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1573),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1581),
.B(n_1543),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1571),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1589),
.B(n_1545),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1580),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1591),
.C(n_1575),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1581),
.B(n_1569),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1591),
.B(n_1550),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1572),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1571),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1543),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1580),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1588),
.B(n_1547),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1579),
.B(n_1556),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1583),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_1559),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1574),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1583),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1581),
.B(n_1559),
.Y(n_1622)
);

NAND2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1546),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1569),
.B(n_1564),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1585),
.B(n_1588),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1569),
.B(n_1564),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1576),
.B(n_1395),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1584),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1585),
.B(n_1567),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1585),
.B(n_1567),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1584),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1586),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1531),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1623),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1607),
.B(n_1555),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1607),
.B(n_1574),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1598),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1593),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1631),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1623),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1594),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1594),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1592),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1597),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1597),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1602),
.B(n_1579),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1575),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1609),
.A2(n_1563),
.B(n_1570),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1600),
.B(n_1577),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1616),
.B(n_1577),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1612),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1577),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1632),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1601),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1599),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1599),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1609),
.A2(n_1558),
.B1(n_1562),
.B2(n_1563),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1627),
.B(n_1566),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1602),
.B(n_1579),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1604),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1604),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1611),
.B(n_1633),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1623),
.B(n_1555),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1596),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1595),
.B(n_1579),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1605),
.B(n_1582),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1655),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1655),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1667),
.B(n_1603),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1638),
.B(n_1611),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_L g1673 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1634),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1647),
.B(n_1595),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1644),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1641),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1647),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1650),
.A2(n_1664),
.B(n_1659),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1649),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1641),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1636),
.B(n_1625),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1638),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1642),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1635),
.B(n_1651),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1636),
.B(n_1629),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1648),
.B(n_1605),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1642),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1645),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1667),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_L g1691 ( 
.A(n_1634),
.B(n_1640),
.C(n_1656),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1648),
.B(n_1614),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1637),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1685),
.A2(n_1665),
.B1(n_1634),
.B2(n_1570),
.C(n_1654),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1670),
.B(n_1653),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1679),
.A2(n_1652),
.B1(n_1667),
.B2(n_1660),
.Y(n_1696)
);

AND2x2_ASAP7_75t_SL g1697 ( 
.A(n_1669),
.B(n_1661),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1686),
.B(n_1637),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1683),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1686),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1682),
.B(n_1669),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1677),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1672),
.A2(n_1570),
.B1(n_1613),
.B2(n_1606),
.C(n_1596),
.Y(n_1703)
);

AOI311xp33_ASAP7_75t_L g1704 ( 
.A1(n_1676),
.A2(n_1639),
.A3(n_1658),
.B(n_1663),
.C(n_1662),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1673),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1677),
.Y(n_1706)
);

OAI21xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1673),
.A2(n_1669),
.B(n_1687),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1681),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1691),
.A2(n_1639),
.B(n_1649),
.C(n_1668),
.Y(n_1709)
);

OAI321xp33_ASAP7_75t_L g1710 ( 
.A1(n_1682),
.A2(n_1613),
.A3(n_1596),
.B1(n_1606),
.B2(n_1620),
.C(n_1610),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1681),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1680),
.A2(n_1610),
.B(n_1613),
.C(n_1606),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1700),
.B(n_1693),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1697),
.B(n_1690),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1707),
.B(n_1671),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1701),
.Y(n_1716)
);

INVxp33_ASAP7_75t_L g1717 ( 
.A(n_1698),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1705),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1699),
.B(n_1693),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_L g1720 ( 
.A(n_1705),
.B(n_1680),
.C(n_1674),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1696),
.B(n_1675),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1709),
.B(n_1678),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1675),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1723),
.B(n_1680),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1715),
.A2(n_1674),
.B(n_1666),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_SL g1726 ( 
.A1(n_1717),
.A2(n_1671),
.B(n_1703),
.Y(n_1726)
);

OAI211xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1722),
.A2(n_1694),
.B(n_1712),
.C(n_1674),
.Y(n_1727)
);

OAI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1720),
.A2(n_1704),
.B(n_1708),
.C(n_1706),
.Y(n_1728)
);

NAND2xp33_ASAP7_75t_L g1729 ( 
.A(n_1721),
.B(n_1674),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1714),
.A2(n_1666),
.B1(n_1692),
.B2(n_1687),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

OAI322xp33_ASAP7_75t_L g1732 ( 
.A1(n_1718),
.A2(n_1711),
.A3(n_1702),
.B1(n_1684),
.B2(n_1688),
.C1(n_1689),
.C2(n_1620),
.Y(n_1732)
);

OAI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1727),
.A2(n_1720),
.B1(n_1713),
.B2(n_1719),
.C(n_1688),
.Y(n_1733)
);

AOI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1728),
.A2(n_1710),
.B(n_1689),
.C(n_1684),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1726),
.A2(n_1710),
.B1(n_1663),
.B2(n_1662),
.C(n_1645),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1724),
.Y(n_1736)
);

O2A1O1Ixp33_ASAP7_75t_SL g1737 ( 
.A1(n_1731),
.A2(n_1646),
.B(n_1657),
.C(n_1629),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1736),
.B(n_1730),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1733),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1737),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1734),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1735),
.B(n_1729),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1736),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1741),
.A2(n_1732),
.B1(n_1725),
.B2(n_1646),
.C(n_1657),
.Y(n_1744)
);

AOI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1738),
.A2(n_1671),
.B(n_1692),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1740),
.B(n_1671),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1739),
.A2(n_1668),
.B1(n_1661),
.B2(n_1590),
.C(n_1615),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_L g1748 ( 
.A(n_1743),
.B(n_1617),
.C(n_1603),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1745),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1746),
.B(n_1742),
.C(n_1617),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1748),
.B(n_1603),
.Y(n_1751)
);

CKINVDCx20_ASAP7_75t_R g1752 ( 
.A(n_1750),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1752),
.B(n_1751),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1753),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1753),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1754),
.A2(n_1749),
.B(n_1744),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1755),
.A2(n_1747),
.B(n_1615),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1756),
.A2(n_1630),
.B1(n_1614),
.B2(n_1608),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1757),
.A2(n_1617),
.B1(n_1603),
.B2(n_1622),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_R g1760 ( 
.A1(n_1758),
.A2(n_1560),
.B1(n_1628),
.B2(n_1608),
.Y(n_1760)
);

XNOR2xp5_ASAP7_75t_L g1761 ( 
.A(n_1760),
.B(n_1759),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1761),
.A2(n_1617),
.B1(n_1622),
.B2(n_1619),
.Y(n_1762)
);

AOI322xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1619),
.A3(n_1626),
.B1(n_1624),
.B2(n_1628),
.C1(n_1618),
.C2(n_1621),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1626),
.B1(n_1624),
.B2(n_1618),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1621),
.B(n_1630),
.C(n_1553),
.Y(n_1765)
);


endmodule