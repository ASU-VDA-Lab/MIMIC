module fake_jpeg_364_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_56),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_63),
.B1(n_45),
.B2(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_50),
.B1(n_49),
.B2(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_78),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_71),
.B(n_70),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_68),
.Y(n_98)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_88),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_51),
.Y(n_106)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_45),
.B1(n_44),
.B2(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_53),
.B1(n_43),
.B2(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_46),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_77),
.C(n_87),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_54),
.B(n_68),
.Y(n_90)
);

NOR4xp25_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_100),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_51),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_106),
.B1(n_10),
.B2(n_11),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_50),
.B1(n_47),
.B2(n_54),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_25),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_1),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_113),
.B1(n_98),
.B2(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_80),
.B1(n_83),
.B2(n_51),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_111),
.B1(n_119),
.B2(n_12),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_117),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_121),
.C(n_98),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_7),
.B(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_9),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_10),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_12),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

OAI322xp33_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_127),
.A3(n_131),
.B1(n_133),
.B2(n_117),
.C1(n_16),
.C2(n_15),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_28),
.C(n_39),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_126),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_109),
.B1(n_16),
.B2(n_19),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_13),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_108),
.B(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_141),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_143),
.Y(n_148)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_132),
.B1(n_128),
.B2(n_137),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_144),
.B1(n_140),
.B2(n_26),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_127),
.C(n_130),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_139),
.C(n_136),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_150),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_151),
.C(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_145),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_17),
.B(n_21),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_29),
.B(n_30),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_31),
.Y(n_157)
);

OAI311xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_32),
.A3(n_33),
.B1(n_34),
.C1(n_37),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_40),
.Y(n_159)
);


endmodule