module fake_jpeg_27759_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_23),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_58),
.Y(n_70)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_54),
.Y(n_97)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_63),
.B(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_24),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_80),
.Y(n_115)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_96),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_17),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_40),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_97),
.B1(n_79),
.B2(n_89),
.Y(n_99)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_95),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_45),
.Y(n_124)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_64),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_43),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_44),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_31),
.B1(n_43),
.B2(n_26),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_45),
.B1(n_37),
.B2(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_24),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_48),
.B(n_40),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_44),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_101),
.B(n_47),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_42),
.C(n_47),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_122),
.C(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_114),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_30),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_47),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_119),
.B(n_51),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_117),
.B(n_78),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_48),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_86),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_48),
.C(n_40),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_126),
.B1(n_97),
.B2(n_51),
.Y(n_143)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_45),
.B1(n_37),
.B2(n_83),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_77),
.C(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_134),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_151),
.C(n_153),
.Y(n_158)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_48),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_139),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_0),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_85),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_142),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_107),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_145),
.B(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_85),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_149),
.B1(n_154),
.B2(n_103),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_97),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_146),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_0),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_116),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_82),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_81),
.B1(n_71),
.B2(n_74),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_71),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_46),
.C(n_38),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_46),
.B1(n_30),
.B2(n_38),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_157),
.A2(n_165),
.B1(n_166),
.B2(n_179),
.Y(n_213)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_181),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_162),
.A2(n_168),
.B(n_170),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_119),
.B1(n_125),
.B2(n_104),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_102),
.B1(n_104),
.B2(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_168),
.B(n_170),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_147),
.C(n_141),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_119),
.C(n_126),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_38),
.C(n_109),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_175),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_132),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_109),
.B1(n_116),
.B2(n_17),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_183),
.Y(n_200)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_36),
.B1(n_34),
.B2(n_32),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_139),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_158),
.Y(n_222)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_205),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_146),
.C(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_199),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_36),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_208),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_145),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_215),
.B(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_34),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_32),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_214),
.Y(n_239)
);

INVx5_ASAP7_75t_SL g211 ( 
.A(n_176),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_25),
.B1(n_28),
.B2(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_29),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_29),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_164),
.A2(n_60),
.B(n_28),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_158),
.B(n_28),
.C(n_25),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_173),
.C(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_228),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_203),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_178),
.B1(n_159),
.B2(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_194),
.C(n_191),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_R g233 ( 
.A(n_217),
.B(n_187),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_212),
.B(n_205),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_189),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_160),
.B1(n_177),
.B2(n_20),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_223),
.B1(n_219),
.B2(n_235),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_192),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_241),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_20),
.Y(n_242)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_243),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_196),
.B(n_18),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_202),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_211),
.B1(n_195),
.B2(n_190),
.Y(n_251)
);

OAI22x1_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_206),
.B1(n_190),
.B2(n_215),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_246),
.A2(n_251),
.B1(n_226),
.B2(n_219),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_248),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_204),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_255),
.B1(n_257),
.B2(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_260),
.C(n_221),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_194),
.C(n_218),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_232),
.B(n_203),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_226),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_236),
.B(n_1),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_279),
.C(n_284),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_250),
.B(n_265),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_225),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_228),
.C(n_230),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_225),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_230),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_220),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_220),
.C(n_244),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_244),
.C(n_223),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_263),
.C(n_252),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_289),
.B(n_294),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_227),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_300),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_255),
.B(n_261),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_299),
.C(n_275),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_251),
.B(n_256),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_294),
.A2(n_292),
.B1(n_291),
.B2(n_290),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_272),
.C(n_274),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_303),
.C(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_275),
.C(n_240),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_239),
.C(n_25),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_8),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_299),
.B1(n_297),
.B2(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_16),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_6),
.B(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_5),
.C(n_6),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_315),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_322),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_8),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.C(n_312),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_9),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_313),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_9),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_320),
.B(n_314),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_328),
.C(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_330),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_308),
.C(n_309),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_310),
.B1(n_14),
.B2(n_15),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_332),
.B(n_333),
.C(n_327),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_329),
.C(n_326),
.Y(n_337)
);

NAND2x1_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_321),
.Y(n_338)
);

AND2x4_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_10),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_14),
.C(n_15),
.Y(n_340)
);


endmodule