module fake_jpeg_15550_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_2),
.B(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_6),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_14),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_20),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_15),
.B1(n_10),
.B2(n_8),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_19),
.B1(n_12),
.B2(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_1),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_7),
.A2(n_4),
.B(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_14),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_23),
.C(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_30),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_17),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_38),
.C(n_26),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_19),
.C(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_30),
.Y(n_39)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_40),
.A3(n_41),
.B1(n_13),
.B2(n_31),
.C1(n_28),
.C2(n_29),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_43),
.C(n_36),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_13),
.A3(n_24),
.B1(n_22),
.B2(n_36),
.C1(n_5),
.C2(n_33),
.Y(n_43)
);


endmodule