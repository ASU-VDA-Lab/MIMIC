module fake_netlist_1_8058_n_20 (n_1, n_2, n_4, n_3, n_0, n_20);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_20;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_7;
INVxp67_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
INVx1_ASAP7_75t_SL g6 ( .A(n_2), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_1), .B(n_3), .Y(n_8) );
OAI21x1_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_0), .B(n_1), .Y(n_9) );
AO21x2_ASAP7_75t_L g10 ( .A1(n_7), .A2(n_0), .B(n_1), .Y(n_10) );
OAI21x1_ASAP7_75t_L g11 ( .A1(n_8), .A2(n_2), .B(n_3), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
NAND3xp33_ASAP7_75t_L g15 ( .A(n_12), .B(n_10), .C(n_11), .Y(n_15) );
NOR3xp33_ASAP7_75t_L g16 ( .A(n_15), .B(n_12), .C(n_6), .Y(n_16) );
AOI321xp33_ASAP7_75t_L g17 ( .A1(n_14), .A2(n_12), .A3(n_13), .B1(n_2), .B2(n_4), .C(n_11), .Y(n_17) );
NAND4xp25_ASAP7_75t_L g18 ( .A(n_17), .B(n_6), .C(n_13), .D(n_4), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
AOI222xp33_ASAP7_75t_SL g20 ( .A1(n_18), .A2(n_4), .B1(n_9), .B2(n_10), .C1(n_19), .C2(n_6), .Y(n_20) );
endmodule