module fake_netlist_1_743_n_721 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_721);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_721;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_482;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_649;
wire n_98;
wire n_527;
wire n_276;
wire n_526;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_15), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_4), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_17), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_22), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_70), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_47), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_15), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_5), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_2), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_68), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_69), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_73), .Y(n_93) );
INVx2_ASAP7_75t_SL g94 ( .A(n_50), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_76), .Y(n_95) );
NOR2xp67_ASAP7_75t_L g96 ( .A(n_7), .B(n_18), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_45), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_4), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_66), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_11), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_41), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_23), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_24), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_39), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_33), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_72), .B(n_58), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_78), .B(n_8), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_48), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_44), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_26), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_59), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_55), .B(n_65), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_35), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_56), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_16), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_16), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_29), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_9), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_6), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_40), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_38), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_34), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_67), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_62), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_117), .B(n_0), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_94), .B(n_1), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_97), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_97), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_97), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_95), .Y(n_136) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_80), .A2(n_30), .B(n_75), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_87), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_94), .B(n_1), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_104), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_88), .B(n_3), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_84), .B(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_80), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_90), .B(n_5), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_88), .B(n_6), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_100), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_121), .B(n_7), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_85), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_104), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_86), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_86), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_121), .B(n_8), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_114), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_119), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_100), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_123), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_115), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_115), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_83), .B(n_9), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_119), .B(n_10), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_91), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_123), .B(n_10), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_92), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_126), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_81), .B(n_82), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_93), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_166), .B(n_126), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_147), .B(n_92), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_165), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_165), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_169), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_171), .B(n_109), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_149), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_160), .B(n_111), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_138), .Y(n_185) );
AND2x6_ASAP7_75t_L g186 ( .A(n_167), .B(n_93), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_138), .A2(n_98), .B1(n_111), .B2(n_124), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_167), .Y(n_188) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_167), .B(n_106), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_160), .B(n_124), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_166), .B(n_122), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_166), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
NOR2xp33_ASAP7_75t_SL g196 ( .A(n_164), .B(n_116), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_145), .B(n_122), .Y(n_199) );
OAI221xp5_ASAP7_75t_L g200 ( .A1(n_161), .A2(n_120), .B1(n_102), .B2(n_103), .C(n_127), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_141), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_129), .B(n_125), .Y(n_202) );
INVxp67_ASAP7_75t_SL g203 ( .A(n_161), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_129), .B(n_116), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_129), .B(n_125), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_145), .B(n_128), .Y(n_206) );
OAI21xp33_ASAP7_75t_L g207 ( .A1(n_151), .A2(n_127), .B(n_118), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_151), .A2(n_112), .B1(n_110), .B2(n_108), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_154), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_171), .B(n_96), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_172), .B(n_99), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_141), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_156), .B(n_105), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_156), .B(n_172), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_168), .B(n_101), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_168), .B(n_106), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_137), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_132), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_141), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_141), .Y(n_224) );
INVxp67_ASAP7_75t_SL g225 ( .A(n_142), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_140), .B(n_107), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_164), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_132), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_152), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
NAND2xp33_ASAP7_75t_SL g232 ( .A(n_146), .B(n_11), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_140), .B(n_113), .Y(n_233) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_131), .B(n_12), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_141), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_153), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_225), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_185), .B(n_146), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_194), .B(n_170), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_177), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_197), .B(n_144), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_195), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_189), .A2(n_157), .B1(n_148), .B2(n_150), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_188), .B(n_170), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_195), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_188), .A2(n_137), .B(n_153), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_189), .A2(n_157), .B1(n_148), .B2(n_150), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_193), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_174), .B(n_142), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_220), .B(n_140), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_188), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_190), .Y(n_253) );
NOR2x1p5_ASAP7_75t_L g254 ( .A(n_183), .B(n_136), .Y(n_254) );
NAND2xp33_ASAP7_75t_L g255 ( .A(n_186), .B(n_170), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_195), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_203), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_214), .B(n_140), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_186), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_191), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_214), .B(n_143), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_204), .Y(n_262) );
AO21x1_ASAP7_75t_L g263 ( .A1(n_221), .A2(n_158), .B(n_153), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_186), .A2(n_162), .B1(n_158), .B2(n_170), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g265 ( .A(n_191), .B(n_143), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_186), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_183), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_175), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_184), .B(n_143), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_186), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_226), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_181), .B(n_143), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_178), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_226), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_214), .Y(n_276) );
AND2x6_ASAP7_75t_L g277 ( .A(n_180), .B(n_162), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g278 ( .A(n_180), .B(n_159), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_230), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_182), .A2(n_162), .B1(n_158), .B2(n_163), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_179), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_221), .A2(n_137), .B(n_130), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_210), .B(n_170), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_181), .B(n_159), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_211), .B(n_170), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_208), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_231), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_196), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_202), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_232), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_202), .A2(n_159), .B1(n_163), .B2(n_137), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_236), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_219), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_202), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_181), .B(n_159), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_202), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_205), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_205), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_212), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_216), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_205), .A2(n_228), .B1(n_187), .B2(n_234), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_221), .B(n_163), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_208), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_215), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_238), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_294), .B(n_234), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_240), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_272), .A2(n_200), .B1(n_232), .B2(n_213), .C(n_206), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_278), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_241), .A2(n_199), .B(n_192), .C(n_207), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_282), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_237), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_257), .B(n_213), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_303), .A2(n_173), .B(n_192), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_276), .A2(n_205), .B1(n_257), .B2(n_262), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_276), .Y(n_317) );
BUFx4f_ASAP7_75t_L g318 ( .A(n_285), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_303), .A2(n_173), .B(n_218), .Y(n_319) );
INVx5_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_250), .A2(n_218), .B(n_217), .C(n_206), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_292), .B(n_209), .C(n_227), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_259), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_253), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_300), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_250), .B(n_205), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_243), .B(n_217), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_272), .A2(n_213), .B1(n_209), .B2(n_227), .C(n_199), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_248), .A2(n_302), .B1(n_291), .B2(n_269), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_289), .B(n_233), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_251), .B(n_163), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_258), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_267), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_281), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_259), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_252), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_261), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_269), .B(n_137), .C(n_163), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g341 ( .A(n_252), .B(n_215), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_266), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_268), .B(n_163), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_279), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g345 ( .A(n_297), .B(n_235), .C(n_224), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_266), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_296), .B(n_12), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_270), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_279), .B(n_13), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_247), .A2(n_235), .B(n_201), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_260), .B(n_13), .Y(n_351) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_273), .A2(n_130), .B(n_134), .C(n_133), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g353 ( .A1(n_296), .A2(n_135), .B(n_133), .C(n_134), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_277), .A2(n_201), .B1(n_224), .B2(n_223), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_278), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_297), .B(n_14), .Y(n_356) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_254), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_260), .A2(n_135), .B(n_134), .C(n_133), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_270), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_340), .A2(n_283), .B(n_263), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_340), .A2(n_239), .B(n_286), .Y(n_361) );
AO32x2_ASAP7_75t_L g362 ( .A1(n_306), .A2(n_290), .A3(n_299), .B1(n_298), .B2(n_280), .Y(n_362) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_323), .A2(n_239), .B(n_284), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_307), .B(n_293), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_323), .A2(n_321), .B(n_319), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_324), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_308), .A2(n_295), .B1(n_277), .B2(n_242), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_312), .B(n_295), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_350), .A2(n_286), .B(n_284), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_309), .A2(n_280), .B1(n_249), .B2(n_244), .C(n_288), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_349), .A2(n_264), .B(n_245), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_346), .Y(n_375) );
NAND3xp33_ASAP7_75t_SL g376 ( .A(n_335), .B(n_265), .C(n_264), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_SL g377 ( .A1(n_352), .A2(n_245), .B(n_256), .C(n_246), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_315), .A2(n_265), .B(n_223), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_355), .B(n_242), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_322), .B(n_277), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_333), .A2(n_274), .B(n_271), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_351), .B(n_358), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_326), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_329), .Y(n_384) );
AOI21xp33_ASAP7_75t_SL g385 ( .A1(n_331), .A2(n_14), .B(n_275), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_313), .B(n_277), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_331), .A2(n_304), .B1(n_287), .B2(n_305), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_SL g390 ( .A1(n_328), .A2(n_327), .B(n_330), .C(n_339), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_135), .B(n_130), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_327), .A2(n_255), .B(n_304), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g393 ( .A1(n_311), .A2(n_304), .B(n_287), .C(n_132), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_364), .B(n_328), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_387), .A2(n_347), .B1(n_325), .B2(n_332), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_387), .B(n_344), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_387), .A2(n_316), .B1(n_314), .B2(n_336), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_383), .B(n_310), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_357), .B1(n_317), .B2(n_356), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_385), .A2(n_318), .B1(n_338), .B2(n_345), .C(n_341), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_385), .A2(n_366), .B(n_365), .C(n_371), .Y(n_401) );
AOI221xp5_ASAP7_75t_SL g402 ( .A1(n_366), .A2(n_359), .B1(n_348), .B2(n_342), .C(n_337), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_369), .A2(n_338), .B(n_320), .C(n_132), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_375), .A2(n_318), .B1(n_320), .B2(n_342), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_383), .A2(n_320), .B1(n_359), .B2(n_342), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_384), .A2(n_359), .B1(n_348), .B2(n_337), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_390), .A2(n_341), .B(n_287), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_384), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_365), .A2(n_348), .B1(n_337), .B2(n_304), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_365), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_377), .A2(n_287), .B(n_229), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_371), .A2(n_229), .B1(n_222), .B2(n_198), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_376), .A2(n_229), .B1(n_222), .B2(n_198), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_371), .B(n_19), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_229), .B1(n_222), .B2(n_198), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_222), .B(n_198), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_389), .A2(n_176), .B1(n_21), .B2(n_25), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_360), .A2(n_176), .B(n_27), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_386), .Y(n_422) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_410), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_408), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_394), .B(n_360), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_397), .B(n_379), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_396), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_395), .B(n_379), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_415), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_398), .B(n_379), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_398), .B(n_386), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_415), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_401), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_401), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_421), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_399), .B(n_373), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_421), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_418), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_396), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_414), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_419), .B(n_380), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_419), .A2(n_422), .B1(n_400), .B2(n_380), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_422), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_414), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_404), .B(n_380), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_409), .B(n_380), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_406), .B(n_363), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_402), .B(n_363), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_407), .B(n_370), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_421), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_403), .A2(n_370), .B1(n_367), .B2(n_388), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_405), .B(n_368), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_417), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_363), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_420), .B(n_367), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_423), .B(n_362), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_427), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_452), .B(n_451), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_437), .B(n_367), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_425), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_424), .B(n_362), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_424), .B(n_381), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_429), .B(n_362), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_441), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_434), .A2(n_392), .B1(n_416), .B2(n_412), .C(n_367), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_440), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_429), .B(n_362), .Y(n_471) );
OAI22x1_ASAP7_75t_L g472 ( .A1(n_446), .A2(n_362), .B1(n_381), .B2(n_31), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_440), .B(n_362), .Y(n_473) );
INVx4_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_451), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_430), .B(n_388), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_430), .B(n_382), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_434), .B(n_388), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_435), .B(n_388), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_442), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_435), .B(n_388), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_433), .B(n_361), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_442), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_433), .B(n_382), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_438), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_426), .B(n_361), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_443), .B(n_391), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_443), .B(n_391), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_447), .B(n_378), .Y(n_491) );
AND2x4_ASAP7_75t_SL g492 ( .A(n_448), .B(n_378), .Y(n_492) );
OAI322xp33_ASAP7_75t_L g493 ( .A1(n_428), .A2(n_411), .A3(n_176), .B1(n_36), .B2(n_37), .C1(n_42), .C2(n_43), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_446), .B(n_374), .Y(n_494) );
OR2x6_ASAP7_75t_L g495 ( .A(n_449), .B(n_372), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_447), .B(n_374), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_431), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_431), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_452), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_432), .B(n_372), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_436), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_444), .A2(n_176), .B1(n_28), .B2(n_46), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_452), .B(n_20), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_432), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_436), .Y(n_506) );
INVx6_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_450), .B(n_49), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_439), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_497), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_475), .B(n_450), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_470), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_475), .B(n_453), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_475), .B(n_453), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_462), .A2(n_455), .B1(n_458), .B2(n_454), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_465), .B(n_457), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_465), .B(n_457), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_468), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_474), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_474), .B(n_456), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_502), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_461), .B(n_456), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_481), .Y(n_524) );
INVx4_ASAP7_75t_L g525 ( .A(n_474), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_465), .B(n_439), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_502), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_481), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_484), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_484), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_498), .B(n_449), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_463), .B(n_51), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_461), .B(n_52), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_460), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_497), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_463), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_474), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_502), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_466), .Y(n_539) );
AOI31xp33_ASAP7_75t_L g540 ( .A1(n_503), .A2(n_53), .A3(n_54), .B(n_57), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_499), .B(n_60), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_497), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_506), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_499), .B(n_61), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_466), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_501), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_505), .A2(n_63), .B1(n_64), .B2(n_79), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_501), .B(n_488), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_483), .B(n_473), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_505), .B(n_473), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_483), .B(n_461), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_461), .B(n_489), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_464), .B(n_487), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_464), .B(n_487), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_478), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_478), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_489), .B(n_490), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_490), .B(n_467), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_486), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_467), .B(n_471), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_506), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_471), .B(n_496), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_496), .B(n_491), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_477), .B(n_500), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_491), .B(n_495), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_495), .B(n_488), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_486), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_495), .B(n_492), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_534), .B(n_507), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_512), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_558), .B(n_507), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_512), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_518), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_549), .B(n_485), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_547), .B(n_459), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_520), .B(n_500), .Y(n_577) );
NOR2xp67_ASAP7_75t_L g578 ( .A(n_520), .B(n_472), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_537), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_547), .B(n_536), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_558), .B(n_507), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_536), .B(n_459), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_518), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_549), .B(n_485), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_524), .Y(n_586) );
NAND2xp67_ASAP7_75t_L g587 ( .A(n_569), .B(n_492), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_515), .A2(n_507), .B1(n_503), .B2(n_508), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_528), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_528), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_529), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_564), .B(n_552), .Y(n_592) );
BUFx2_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_556), .B(n_507), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_529), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_522), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_510), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_519), .B(n_485), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_520), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_564), .B(n_492), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_552), .B(n_508), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_551), .B(n_494), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_550), .B(n_494), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_513), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_538), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_550), .B(n_495), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_553), .B(n_500), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_553), .B(n_500), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_520), .Y(n_610) );
NOR2x1_ASAP7_75t_R g611 ( .A(n_525), .B(n_504), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_563), .B(n_477), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_515), .A2(n_504), .B1(n_477), .B2(n_495), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_535), .A2(n_504), .B(n_493), .C(n_477), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_530), .Y(n_616) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_525), .B(n_504), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_525), .B(n_476), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_530), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_559), .B(n_509), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_548), .B(n_469), .C(n_480), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_559), .B(n_509), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_588), .A2(n_567), .B1(n_542), .B2(n_523), .Y(n_623) );
OA21x2_ASAP7_75t_L g624 ( .A1(n_614), .A2(n_556), .B(n_557), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_578), .A2(n_540), .B(n_548), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_598), .B(n_557), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_617), .A2(n_525), .B1(n_521), .B2(n_533), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_570), .A2(n_567), .B1(n_566), .B2(n_523), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_607), .A2(n_566), .B1(n_531), .B2(n_511), .C(n_569), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_580), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_600), .B(n_533), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_599), .B(n_568), .Y(n_633) );
OAI222xp33_ASAP7_75t_L g634 ( .A1(n_600), .A2(n_533), .B1(n_561), .B2(n_511), .C1(n_523), .C2(n_563), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_571), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_570), .A2(n_545), .B(n_541), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_573), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_592), .B(n_561), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_617), .A2(n_533), .B(n_565), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_605), .B(n_568), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_574), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_594), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_583), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_593), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_610), .A2(n_521), .B(n_532), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_611), .A2(n_472), .B(n_493), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_575), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g648 ( .A1(n_615), .A2(n_523), .A3(n_532), .B1(n_565), .B2(n_513), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_585), .Y(n_649) );
OAI222xp33_ASAP7_75t_L g650 ( .A1(n_579), .A2(n_565), .B1(n_546), .B2(n_539), .C1(n_560), .C2(n_554), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_572), .B(n_565), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_594), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_586), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_589), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_621), .A2(n_560), .B1(n_517), .B2(n_516), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_605), .B(n_514), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_584), .Y(n_657) );
INVxp33_ASAP7_75t_L g658 ( .A(n_618), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_618), .A2(n_517), .B1(n_516), .B2(n_539), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_590), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_655), .B(n_582), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_626), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_647), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_657), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_631), .B(n_579), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_638), .B(n_612), .Y(n_666) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_655), .A2(n_595), .B1(n_582), .B2(n_576), .C1(n_602), .C2(n_581), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g668 ( .A1(n_623), .A2(n_609), .A3(n_608), .B1(n_576), .B2(n_595), .C1(n_601), .C2(n_619), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_640), .B(n_604), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_656), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_623), .A2(n_639), .B1(n_625), .B2(n_640), .Y(n_671) );
OAI22xp33_ASAP7_75t_SL g672 ( .A1(n_630), .A2(n_587), .B1(n_577), .B2(n_620), .Y(n_672) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_627), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_635), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_637), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_644), .B(n_622), .Y(n_676) );
OAI222xp33_ASAP7_75t_L g677 ( .A1(n_648), .A2(n_577), .B1(n_603), .B2(n_596), .C1(n_591), .C2(n_616), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_641), .Y(n_678) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_646), .A2(n_606), .B(n_546), .C(n_555), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_642), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_643), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_634), .A2(n_606), .B(n_597), .C(n_613), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_642), .Y(n_683) );
AOI21xp33_ASAP7_75t_SL g684 ( .A1(n_628), .A2(n_597), .B(n_514), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_671), .A2(n_658), .B1(n_659), .B2(n_629), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_679), .A2(n_627), .B1(n_633), .B2(n_659), .Y(n_686) );
NAND5xp2_ASAP7_75t_L g687 ( .A(n_667), .B(n_632), .C(n_645), .D(n_636), .E(n_633), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_662), .Y(n_688) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_661), .A2(n_651), .A3(n_654), .B1(n_653), .B2(n_660), .C1(n_649), .C2(n_652), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_684), .A2(n_624), .B(n_652), .C(n_469), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_682), .A2(n_650), .B(n_632), .C(n_624), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_663), .Y(n_692) );
OAI211xp5_ASAP7_75t_SL g693 ( .A1(n_668), .A2(n_527), .B(n_544), .C(n_562), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_673), .A2(n_624), .B1(n_527), .B2(n_544), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_672), .A2(n_526), .B1(n_544), .B2(n_527), .C(n_562), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_674), .Y(n_696) );
NAND2xp33_ASAP7_75t_SL g697 ( .A(n_669), .B(n_543), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_664), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_698), .B(n_670), .Y(n_699) );
OAI22xp33_ASAP7_75t_SL g700 ( .A1(n_685), .A2(n_665), .B1(n_681), .B2(n_678), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g701 ( .A1(n_695), .A2(n_677), .B1(n_665), .B2(n_675), .C1(n_680), .C2(n_666), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_689), .B(n_666), .Y(n_702) );
XOR2xp5_ASAP7_75t_L g703 ( .A(n_686), .B(n_676), .Y(n_703) );
AOI32xp33_ASAP7_75t_L g704 ( .A1(n_693), .A2(n_680), .A3(n_676), .B1(n_683), .B2(n_526), .Y(n_704) );
AND4x1_ASAP7_75t_L g705 ( .A(n_691), .B(n_476), .C(n_479), .D(n_480), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_697), .Y(n_706) );
NAND3xp33_ASAP7_75t_SL g707 ( .A(n_701), .B(n_691), .C(n_692), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_700), .A2(n_687), .B(n_694), .Y(n_708) );
NAND4xp75_ASAP7_75t_L g709 ( .A(n_702), .B(n_696), .C(n_688), .D(n_690), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_703), .B(n_683), .Y(n_710) );
NOR2x1p5_ASAP7_75t_L g711 ( .A(n_705), .B(n_538), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_707), .Y(n_713) );
NOR3xp33_ASAP7_75t_SL g714 ( .A(n_709), .B(n_699), .C(n_706), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_712), .Y(n_715) );
BUFx2_ASAP7_75t_SL g716 ( .A(n_713), .Y(n_716) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_715), .A2(n_714), .B1(n_708), .B2(n_711), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_717), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_716), .B(n_704), .Y(n_719) );
AOI22xp5_ASAP7_75t_SL g720 ( .A1(n_719), .A2(n_479), .B1(n_482), .B2(n_543), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_509), .B(n_482), .Y(n_721) );
endmodule