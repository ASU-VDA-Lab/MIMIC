module fake_netlist_5_1842_n_1446 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1446);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1446;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_370;
wire n_976;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

INVx1_ASAP7_75t_L g366 ( 
.A(n_76),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_35),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_47),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_176),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_304),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_129),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_360),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_91),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_184),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_46),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_225),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_268),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_69),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_201),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_353),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_205),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_83),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_58),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_1),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_87),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_166),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_237),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_104),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_44),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_16),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_31),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_249),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_291),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_136),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_98),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_28),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_150),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_280),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_295),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_224),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_239),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_209),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_233),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_327),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_306),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_352),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_0),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_349),
.Y(n_411)
);

BUFx8_ASAP7_75t_SL g412 ( 
.A(n_174),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_118),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_51),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_271),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_214),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_298),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_193),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_269),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_11),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_194),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_57),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_216),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_191),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_278),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_198),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_259),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_330),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_77),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_153),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_339),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_133),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_23),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_138),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_345),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_134),
.Y(n_438)
);

BUFx2_ASAP7_75t_SL g439 ( 
.A(n_88),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_192),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_263),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_12),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_253),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_354),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_283),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_50),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_169),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_165),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_59),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_247),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_9),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_163),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_343),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_135),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_15),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_63),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_234),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_66),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_105),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_185),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_96),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_270),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_74),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_261),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_127),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_211),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_52),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_128),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_14),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_294),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_85),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g474 ( 
.A(n_203),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_199),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_71),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_337),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_358),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_189),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_36),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_3),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_260),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_362),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_48),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_273),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_97),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_267),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_38),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_255),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_266),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_152),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_335),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_332),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_320),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_148),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_137),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_61),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_86),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_226),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_361),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_334),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_93),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_28),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_318),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_236),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_52),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_17),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_218),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_336),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_340),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_212),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_50),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_139),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_65),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_103),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_81),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_309),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_238),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_302),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_24),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_142),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_110),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_7),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_124),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_125),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_262),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_62),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_299),
.Y(n_528)
);

HB1xp67_ASAP7_75t_SL g529 ( 
.A(n_229),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_82),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_257),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_235),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_54),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_145),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_70),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_202),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_180),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_122),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_279),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_210),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_301),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_364),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_344),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_231),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_33),
.Y(n_545)
);

BUFx8_ASAP7_75t_SL g546 ( 
.A(n_217),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_341),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_42),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_140),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_325),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_346),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_44),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_200),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_250),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_221),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_305),
.Y(n_556)
);

CKINVDCx14_ASAP7_75t_R g557 ( 
.A(n_351),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_40),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_365),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_42),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_25),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_92),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_47),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_222),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_156),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_38),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_272),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_73),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_53),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_72),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_144),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_258),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_316),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_9),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_230),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_244),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_323),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_506),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_367),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_420),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_406),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_425),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_523),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_523),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_370),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_569),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_373),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_441),
.Y(n_589)
);

INVxp67_ASAP7_75t_SL g590 ( 
.A(n_459),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_377),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_541),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_375),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_551),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_384),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_393),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_418),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_383),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_399),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_564),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_368),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_443),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_478),
.B(n_0),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_452),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_389),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_450),
.Y(n_606)
);

INVxp67_ASAP7_75t_SL g607 ( 
.A(n_376),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_469),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_394),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_480),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_397),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_520),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_395),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_561),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_396),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_402),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_436),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_378),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_450),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_569),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_398),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_367),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_402),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_378),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_463),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_484),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_468),
.B(n_1),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_463),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_401),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_467),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_474),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_461),
.Y(n_635)
);

INVxp33_ASAP7_75t_SL g636 ( 
.A(n_391),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_467),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_412),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_403),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_461),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_498),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_380),
.B(n_2),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_366),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_392),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_369),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_409),
.B(n_2),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_404),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_407),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_413),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_422),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_423),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_371),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_372),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_498),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_410),
.Y(n_655)
);

NOR2xp67_ASAP7_75t_L g656 ( 
.A(n_387),
.B(n_3),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_387),
.B(n_4),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_381),
.B(n_411),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_374),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_424),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_379),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_382),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_412),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_414),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_426),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_428),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_385),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_435),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_386),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_546),
.Y(n_670)
);

NOR2xp67_ASAP7_75t_L g671 ( 
.A(n_390),
.B(n_4),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_390),
.B(n_5),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_432),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_546),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_388),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_405),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_438),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_447),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_408),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_416),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_417),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_421),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_456),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_607),
.A2(n_474),
.B1(n_557),
.B2(n_503),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_643),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_619),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_645),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_652),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_581),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_668),
.B(n_557),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_586),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_583),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_653),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_588),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_659),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_SL g696 ( 
.A(n_638),
.B(n_488),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_591),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_661),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_601),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_593),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_662),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_667),
.Y(n_702)
);

AND2x2_ASAP7_75t_SL g703 ( 
.A(n_597),
.B(n_400),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_613),
.A2(n_512),
.B1(n_533),
.B2(n_507),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_587),
.B(n_466),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_619),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_626),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_626),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_SL g709 ( 
.A1(n_579),
.A2(n_548),
.B1(n_552),
.B2(n_545),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_630),
.B(n_558),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_598),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_669),
.Y(n_712)
);

BUFx8_ASAP7_75t_L g713 ( 
.A(n_621),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_593),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_596),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_596),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_605),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_634),
.B(n_555),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_609),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_592),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_587),
.B(n_554),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_636),
.B(n_555),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_644),
.B(n_664),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_675),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_578),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_658),
.B(n_483),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_595),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_615),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_618),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_599),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_602),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_604),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_676),
.Y(n_733)
);

NOR2x1_ASAP7_75t_L g734 ( 
.A(n_656),
.B(n_439),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_579),
.A2(n_566),
.B1(n_574),
.B2(n_563),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_624),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_679),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_680),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_681),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_682),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_589),
.B(n_400),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_582),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_590),
.B(n_415),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_584),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_655),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_632),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_578),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_678),
.Y(n_748)
);

XOR2xp5_ASAP7_75t_L g749 ( 
.A(n_594),
.B(n_440),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_639),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_647),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_608),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_585),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_600),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_610),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_606),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_611),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_612),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_614),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_622),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_616),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_617),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_627),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_SL g764 ( 
.A(n_638),
.B(n_415),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_628),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_631),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_633),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_637),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_657),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_690),
.B(n_683),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_710),
.B(n_648),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_726),
.B(n_649),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_710),
.B(n_650),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_691),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_745),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_763),
.B(n_765),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_699),
.B(n_651),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_707),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_766),
.B(n_767),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_694),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_757),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_704),
.B(n_580),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_748),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_723),
.B(n_660),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_714),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_697),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_741),
.B(n_419),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_686),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_703),
.B(n_665),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_759),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_725),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_723),
.B(n_623),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_734),
.B(n_666),
.Y(n_793)
);

AND2x6_ASAP7_75t_L g794 ( 
.A(n_741),
.B(n_419),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_686),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_686),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_762),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_705),
.B(n_620),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_706),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_685),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_706),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_684),
.B(n_673),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_705),
.B(n_677),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_687),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_706),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_769),
.A2(n_630),
.B1(n_603),
.B2(n_642),
.Y(n_806)
);

AND2x6_ASAP7_75t_L g807 ( 
.A(n_743),
.B(n_538),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_718),
.B(n_603),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_721),
.B(n_553),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_711),
.B(n_642),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_688),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_714),
.Y(n_812)
);

INVx4_ASAP7_75t_SL g813 ( 
.A(n_709),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_768),
.B(n_671),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_721),
.B(n_571),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_714),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_743),
.B(n_646),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_708),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_708),
.B(n_442),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_708),
.B(n_448),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_756),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_727),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_727),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_693),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_725),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_695),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_R g827 ( 
.A(n_717),
.B(n_646),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_698),
.Y(n_828)
);

OAI21xp33_ASAP7_75t_L g829 ( 
.A1(n_722),
.A2(n_702),
.B(n_701),
.Y(n_829)
);

BUFx4f_ASAP7_75t_L g830 ( 
.A(n_727),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_712),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_747),
.B(n_672),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_732),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_719),
.B(n_635),
.Y(n_834)
);

BUFx6f_ASAP7_75t_SL g835 ( 
.A(n_724),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_747),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_733),
.A2(n_577),
.B1(n_538),
.B2(n_445),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_764),
.B(n_427),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_760),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_728),
.B(n_451),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_737),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_738),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_739),
.B(n_429),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_740),
.B(n_742),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_744),
.B(n_453),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_689),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_729),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_753),
.B(n_716),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_732),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_736),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_746),
.A2(n_529),
.B1(n_455),
.B2(n_457),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_730),
.B(n_577),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_732),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_731),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_750),
.B(n_640),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_752),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_755),
.B(n_430),
.Y(n_857)
);

AND2x6_ASAP7_75t_L g858 ( 
.A(n_758),
.B(n_402),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_751),
.B(n_454),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_761),
.B(n_460),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_700),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_700),
.Y(n_862)
);

AND3x1_ASAP7_75t_L g863 ( 
.A(n_802),
.B(n_735),
.C(n_709),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_770),
.B(n_641),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_772),
.B(n_431),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_828),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_817),
.B(n_787),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_828),
.Y(n_868)
);

BUFx8_ASAP7_75t_L g869 ( 
.A(n_835),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_806),
.A2(n_433),
.B1(n_437),
.B2(n_434),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_771),
.B(n_735),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_773),
.B(n_696),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_784),
.B(n_462),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_830),
.B(n_464),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_787),
.A2(n_444),
.B1(n_449),
.B2(n_446),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_862),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_822),
.B(n_465),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_832),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_787),
.B(n_794),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_777),
.B(n_749),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_831),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_822),
.B(n_472),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_831),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_783),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_791),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_794),
.B(n_458),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_856),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_794),
.B(n_470),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_783),
.B(n_715),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_775),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_832),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_803),
.B(n_475),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_807),
.B(n_473),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_807),
.B(n_477),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_851),
.B(n_654),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_782),
.A2(n_485),
.B1(n_489),
.B2(n_479),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_807),
.B(n_490),
.Y(n_897)
);

OR2x6_ASAP7_75t_L g898 ( 
.A(n_847),
.B(n_692),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_825),
.B(n_715),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_781),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_790),
.A2(n_495),
.B1(n_501),
.B2(n_491),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_853),
.B(n_508),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_778),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_L g904 ( 
.A(n_829),
.B(n_482),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_797),
.B(n_509),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_836),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_778),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_789),
.B(n_810),
.Y(n_908)
);

NOR2x1p5_ASAP7_75t_L g909 ( 
.A(n_774),
.B(n_663),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_798),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_800),
.B(n_510),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_838),
.A2(n_519),
.B(n_521),
.C(n_517),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_804),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_786),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_809),
.B(n_486),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_840),
.B(n_670),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_811),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_780),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_815),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_824),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_826),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_841),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_842),
.B(n_528),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_823),
.B(n_531),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_854),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_SL g926 ( 
.A1(n_808),
.A2(n_625),
.B1(n_629),
.B2(n_720),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_854),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_848),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_799),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_819),
.A2(n_542),
.B(n_537),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_792),
.B(n_625),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_799),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_823),
.B(n_549),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_792),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_776),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_849),
.B(n_55),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_776),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_785),
.B(n_550),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_814),
.B(n_487),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_859),
.B(n_674),
.Y(n_940)
);

AND2x6_ASAP7_75t_SL g941 ( 
.A(n_834),
.B(n_556),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_812),
.B(n_562),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_779),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_779),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_816),
.B(n_567),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_850),
.B(n_786),
.Y(n_946)
);

INVx8_ASAP7_75t_L g947 ( 
.A(n_808),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_857),
.B(n_572),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_855),
.B(n_754),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_844),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_788),
.B(n_492),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_795),
.B(n_493),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_796),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_857),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_845),
.B(n_629),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_860),
.B(n_494),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_801),
.B(n_402),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_805),
.B(n_496),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_L g959 ( 
.A(n_821),
.B(n_499),
.C(n_497),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_818),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_908),
.A2(n_843),
.B(n_814),
.C(n_793),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_918),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_866),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_889),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_919),
.B(n_839),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_949),
.B(n_827),
.Y(n_966)
);

AND2x6_ASAP7_75t_L g967 ( 
.A(n_879),
.B(n_846),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_950),
.B(n_833),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_928),
.B(n_837),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_914),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_865),
.B(n_820),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_903),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_884),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_868),
.B(n_861),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_881),
.Y(n_975)
);

NOR2x1p5_ASAP7_75t_L g976 ( 
.A(n_931),
.B(n_813),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_960),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_910),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_898),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_880),
.B(n_713),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_960),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_L g982 ( 
.A(n_867),
.B(n_852),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_890),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_883),
.B(n_852),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_898),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_937),
.B(n_813),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_871),
.A2(n_852),
.B1(n_502),
.B2(n_504),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_922),
.B(n_861),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_872),
.B(n_861),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_929),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_899),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_907),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_917),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_900),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_864),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_934),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_929),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_899),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_870),
.B(n_500),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_913),
.B(n_505),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_921),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_929),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_925),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_920),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_887),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_946),
.B(n_511),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_955),
.B(n_513),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_954),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_863),
.A2(n_515),
.B1(n_516),
.B2(n_514),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_956),
.B(n_518),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_SL g1011 ( 
.A(n_926),
.B(n_524),
.C(n_522),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_896),
.A2(n_476),
.B1(n_445),
.B2(n_858),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_935),
.B(n_525),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_885),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_885),
.B(n_445),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_932),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_906),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_943),
.B(n_56),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_944),
.B(n_526),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_876),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_927),
.B(n_60),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_898),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_948),
.Y(n_1023)
);

NOR2x2_ASAP7_75t_L g1024 ( 
.A(n_926),
.B(n_713),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_953),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_905),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_878),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_911),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_923),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_947),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_902),
.B(n_527),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_891),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_984),
.A2(n_888),
.B(n_886),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1026),
.B(n_948),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_962),
.B(n_909),
.Y(n_1035)
);

AO31x2_ASAP7_75t_L g1036 ( 
.A1(n_961),
.A2(n_912),
.A3(n_893),
.B(n_897),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_SL g1037 ( 
.A1(n_971),
.A2(n_894),
.B(n_875),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_966),
.B(n_916),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_971),
.A2(n_952),
.B(n_951),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_973),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_989),
.A2(n_933),
.B(n_924),
.Y(n_1041)
);

OA21x2_ASAP7_75t_L g1042 ( 
.A1(n_984),
.A2(n_930),
.B(n_938),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_969),
.A2(n_875),
.B1(n_895),
.B2(n_947),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_SL g1044 ( 
.A1(n_968),
.A2(n_945),
.B(n_942),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1028),
.B(n_873),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_977),
.A2(n_958),
.B(n_936),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_977),
.A2(n_981),
.B(n_1015),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1029),
.B(n_915),
.Y(n_1048)
);

AO31x2_ASAP7_75t_L g1049 ( 
.A1(n_1010),
.A2(n_940),
.A3(n_936),
.B(n_904),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_999),
.A2(n_874),
.B(n_892),
.C(n_939),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1007),
.B(n_959),
.Y(n_1051)
);

INVx3_ASAP7_75t_SL g1052 ( 
.A(n_985),
.Y(n_1052)
);

BUFx12f_ASAP7_75t_L g1053 ( 
.A(n_1030),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_1017),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_995),
.B(n_947),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_969),
.A2(n_901),
.B1(n_882),
.B2(n_877),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_SL g1057 ( 
.A1(n_968),
.A2(n_67),
.B(n_64),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_1010),
.A2(n_957),
.A3(n_858),
.B(n_941),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_981),
.A2(n_957),
.B(n_75),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_963),
.B(n_530),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_972),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_982),
.A2(n_476),
.B(n_445),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_1015),
.A2(n_957),
.B(n_78),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1014),
.A2(n_476),
.B(n_532),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_975),
.A2(n_957),
.B(n_535),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_1021),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_994),
.B(n_534),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1031),
.A2(n_476),
.B(n_536),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1001),
.B(n_539),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_998),
.B(n_68),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_992),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_974),
.A2(n_858),
.B(n_543),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1025),
.A2(n_80),
.B(n_79),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_991),
.B(n_84),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1031),
.B(n_540),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_995),
.B(n_544),
.Y(n_1076)
);

AO31x2_ASAP7_75t_L g1077 ( 
.A1(n_999),
.A2(n_7),
.A3(n_5),
.B(n_6),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1020),
.A2(n_90),
.B(n_89),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1005),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_973),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_965),
.B(n_869),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_993),
.A2(n_95),
.B(n_94),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1004),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1000),
.A2(n_559),
.B(n_547),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1013),
.A2(n_568),
.B(n_565),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_1017),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1008),
.A2(n_570),
.B(n_573),
.C(n_575),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1018),
.A2(n_576),
.B1(n_869),
.B2(n_182),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1017),
.B(n_99),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_1000),
.A2(n_101),
.B(n_100),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1018),
.A2(n_183),
.B1(n_356),
.B2(n_355),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1019),
.A2(n_106),
.B(n_102),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_991),
.B(n_6),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1040),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_1080),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_1033),
.A2(n_1019),
.B(n_1012),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1054),
.B(n_986),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1079),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1046),
.A2(n_988),
.B(n_1027),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1066),
.A2(n_1009),
.B1(n_1021),
.B2(n_987),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_1066),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1086),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1079),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_1053),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1047),
.A2(n_997),
.B(n_1006),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1073),
.A2(n_1022),
.B(n_978),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1034),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1061),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1071),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1078),
.A2(n_976),
.B(n_967),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1083),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1093),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1070),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1082),
.A2(n_967),
.B(n_996),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1074),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1059),
.A2(n_967),
.B(n_1016),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1070),
.Y(n_1117)
);

OAI211xp5_ASAP7_75t_L g1118 ( 
.A1(n_1088),
.A2(n_980),
.B(n_964),
.C(n_1011),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_1074),
.B(n_990),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1039),
.A2(n_1023),
.B(n_1016),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_1052),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1062),
.A2(n_967),
.B(n_1003),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1050),
.A2(n_986),
.B(n_979),
.C(n_1032),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1041),
.A2(n_983),
.B(n_990),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1076),
.B(n_1032),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1038),
.B(n_1032),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1037),
.A2(n_1056),
.B(n_1092),
.Y(n_1127)
);

CKINVDCx11_ASAP7_75t_R g1128 ( 
.A(n_1043),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1055),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1048),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1045),
.B(n_990),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1042),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1042),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1044),
.A2(n_1002),
.B(n_108),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_1091),
.Y(n_1135)
);

NAND2x1p5_ASAP7_75t_L g1136 ( 
.A(n_1089),
.B(n_1002),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1051),
.B(n_1002),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1068),
.A2(n_970),
.B(n_109),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_1081),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1035),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_1057),
.B(n_1024),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1063),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1060),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1088),
.B(n_363),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1075),
.A2(n_111),
.B(n_107),
.Y(n_1145)
);

NOR2x1_ASAP7_75t_SL g1146 ( 
.A(n_1135),
.B(n_1072),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1098),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1127),
.A2(n_1087),
.B(n_1084),
.C(n_1069),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1144),
.A2(n_1128),
.B1(n_1135),
.B2(n_1127),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1135),
.A2(n_1091),
.B(n_1065),
.C(n_1067),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1143),
.A2(n_1064),
.B(n_1085),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1103),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1132),
.A2(n_1049),
.A3(n_1036),
.B(n_1090),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1138),
.B(n_1090),
.C(n_1049),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_SL g1155 ( 
.A(n_1138),
.B(n_1049),
.C(n_1058),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1129),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1094),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_1101),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1097),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1107),
.B(n_1077),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1108),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1101),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1094),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_L g1164 ( 
.A(n_1135),
.B(n_1058),
.Y(n_1164)
);

OAI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_1145),
.A2(n_1036),
.B1(n_1058),
.B2(n_1077),
.C(n_12),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1130),
.B(n_1107),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1095),
.B(n_1137),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1144),
.A2(n_1077),
.B1(n_1036),
.B2(n_11),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1109),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1111),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1115),
.B(n_112),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1097),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1095),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1115),
.B(n_113),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1112),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1125),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_1176)
);

CKINVDCx16_ASAP7_75t_R g1177 ( 
.A(n_1139),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1124),
.Y(n_1178)
);

INVx5_ASAP7_75t_L g1179 ( 
.A(n_1101),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1113),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1126),
.B(n_114),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1145),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_SL g1183 ( 
.A(n_1140),
.B(n_18),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1117),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1131),
.B(n_19),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1102),
.B(n_20),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1118),
.A2(n_1100),
.B1(n_1121),
.B2(n_1141),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1099),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1123),
.B(n_20),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1118),
.B(n_115),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1119),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1101),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1105),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1100),
.B(n_21),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1141),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1141),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1119),
.B(n_26),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1136),
.A2(n_1104),
.B1(n_1120),
.B2(n_1096),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1110),
.B(n_1120),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1136),
.A2(n_1134),
.B1(n_1096),
.B2(n_1116),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1106),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1133),
.B(n_26),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1194),
.A2(n_1142),
.B1(n_1114),
.B2(n_1122),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1156),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1161),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1196),
.A2(n_1195),
.B1(n_1149),
.B2(n_1177),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1182),
.A2(n_1142),
.B1(n_29),
.B2(n_30),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1185),
.B(n_116),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1167),
.B(n_117),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1163),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1190),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1197),
.B(n_119),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1183),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_1213)
);

OAI211xp5_ASAP7_75t_L g1214 ( 
.A1(n_1175),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1150),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1215)
);

AOI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_1176),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_1216)
);

OAI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1148),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.C(n_43),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1189),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1187),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1168),
.A2(n_1181),
.B1(n_1180),
.B2(n_1171),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1157),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1171),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1174),
.A2(n_54),
.B1(n_120),
.B2(n_121),
.Y(n_1223)
);

AOI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1166),
.A2(n_1173),
.B1(n_1165),
.B2(n_1186),
.C1(n_1174),
.C2(n_1170),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1154),
.A2(n_1155),
.B(n_1151),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1191),
.B(n_123),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1202),
.A2(n_1169),
.B1(n_1184),
.B2(n_1147),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1172),
.Y(n_1228)
);

OAI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1198),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.C(n_132),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1164),
.A2(n_141),
.B1(n_143),
.B2(n_146),
.Y(n_1230)
);

OAI211xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1159),
.A2(n_147),
.B(n_149),
.C(n_151),
.Y(n_1231)
);

AOI221xp5_ASAP7_75t_L g1232 ( 
.A1(n_1160),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.C(n_158),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1158),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1172),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_1234)
);

AOI211xp5_ASAP7_75t_L g1235 ( 
.A1(n_1172),
.A2(n_162),
.B(n_164),
.C(n_167),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1152),
.B(n_168),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1199),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1199),
.A2(n_173),
.B1(n_175),
.B2(n_177),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1179),
.A2(n_1192),
.B1(n_1158),
.B2(n_1162),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1200),
.A2(n_1193),
.B(n_1201),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1162),
.B(n_178),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1179),
.A2(n_179),
.B1(n_181),
.B2(n_186),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1179),
.B(n_187),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1178),
.B(n_188),
.C(n_190),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1188),
.A2(n_195),
.B(n_196),
.Y(n_1245)
);

INVx5_ASAP7_75t_SL g1246 ( 
.A(n_1146),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1153),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1153),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1192),
.A2(n_197),
.B1(n_204),
.B2(n_206),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1153),
.A2(n_207),
.B(n_208),
.Y(n_1250)
);

CKINVDCx10_ASAP7_75t_R g1251 ( 
.A(n_1177),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1156),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1167),
.B(n_213),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1149),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_1254)
);

OAI21xp33_ASAP7_75t_L g1255 ( 
.A1(n_1194),
.A2(n_223),
.B(n_227),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1187),
.A2(n_228),
.B1(n_232),
.B2(n_240),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1233),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1225),
.B(n_1240),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1225),
.B(n_241),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1240),
.B(n_242),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1221),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1205),
.B(n_1247),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1248),
.B(n_243),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1210),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1250),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1246),
.B(n_245),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1224),
.B(n_246),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1233),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1227),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1250),
.B(n_1203),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1246),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1239),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1251),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1253),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1246),
.B(n_248),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1228),
.B(n_251),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1217),
.A2(n_252),
.B1(n_254),
.B2(n_256),
.C(n_264),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1209),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1236),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1226),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1245),
.B(n_265),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1245),
.B(n_274),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1244),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1208),
.B(n_275),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1226),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1215),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1212),
.B(n_276),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1243),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1241),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1220),
.B(n_277),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1235),
.A2(n_281),
.B(n_282),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1229),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1231),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1207),
.B(n_284),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1256),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1230),
.B(n_285),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1206),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1204),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1261),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1262),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1297),
.A2(n_1216),
.B1(n_1232),
.B2(n_1242),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1261),
.B(n_1218),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1271),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1257),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1258),
.B(n_1211),
.C(n_1213),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1269),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1264),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1262),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1258),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1274),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1265),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1265),
.A2(n_1214),
.B(n_1255),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1264),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1267),
.A2(n_1219),
.B(n_1249),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1277),
.B(n_1222),
.C(n_1223),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1270),
.B(n_1289),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1271),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1268),
.Y(n_1318)
);

AOI211xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1291),
.A2(n_1252),
.B(n_1254),
.C(n_1238),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1268),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1273),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1268),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1270),
.B(n_1237),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1309),
.B(n_1289),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1316),
.B(n_1283),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1304),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1321),
.B(n_1298),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1310),
.B(n_1298),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1303),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1316),
.B(n_1278),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1308),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1306),
.B(n_1283),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1307),
.B(n_1278),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1300),
.B(n_1279),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1321),
.B(n_1279),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1313),
.B(n_1278),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1299),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1320),
.B(n_1272),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1303),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1317),
.B(n_1272),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1318),
.Y(n_1341)
);

OAI31xp33_ASAP7_75t_L g1342 ( 
.A1(n_1332),
.A2(n_1297),
.A3(n_1305),
.B(n_1301),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1340),
.B(n_1320),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1340),
.B(n_1322),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1329),
.Y(n_1345)
);

NOR2x1_ASAP7_75t_L g1346 ( 
.A(n_1332),
.B(n_1272),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1333),
.B(n_1322),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1338),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1339),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1334),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1328),
.B(n_1304),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1325),
.A2(n_1315),
.B(n_1314),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1326),
.B(n_1304),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1343),
.B(n_1344),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1353),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1348),
.B(n_1325),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1350),
.B(n_1324),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1345),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1346),
.B(n_1342),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1351),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1352),
.Y(n_1361)
);

AND2x4_ASAP7_75t_SL g1362 ( 
.A(n_1347),
.B(n_1327),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1352),
.B(n_1324),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1345),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1349),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1353),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1342),
.B(n_1330),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1358),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1359),
.A2(n_1319),
.B(n_1273),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1362),
.Y(n_1370)
);

OAI222xp33_ASAP7_75t_L g1371 ( 
.A1(n_1361),
.A2(n_1323),
.B1(n_1295),
.B2(n_1259),
.C1(n_1302),
.C2(n_1282),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1355),
.Y(n_1372)
);

OAI322xp33_ASAP7_75t_L g1373 ( 
.A1(n_1363),
.A2(n_1334),
.A3(n_1323),
.B1(n_1286),
.B2(n_1337),
.C1(n_1331),
.C2(n_1302),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1367),
.A2(n_1259),
.B(n_1281),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1365),
.B(n_1335),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1354),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1368),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1369),
.B(n_1360),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1371),
.A2(n_1355),
.B(n_1366),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1372),
.B(n_1356),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1370),
.B(n_1364),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1374),
.A2(n_1372),
.B1(n_1375),
.B2(n_1295),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1376),
.B(n_1358),
.Y(n_1383)
);

INVxp33_ASAP7_75t_L g1384 ( 
.A(n_1373),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1377),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1383),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1381),
.B(n_1357),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_R g1388 ( 
.A(n_1380),
.B(n_1266),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1378),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1384),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1382),
.B(n_1379),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1391),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1390),
.A2(n_1382),
.B1(n_1281),
.B2(n_1290),
.Y(n_1393)
);

OAI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1389),
.A2(n_1286),
.B1(n_1292),
.B2(n_1290),
.C(n_1326),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1386),
.B(n_1341),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1387),
.B(n_1336),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1385),
.A2(n_1281),
.B1(n_1282),
.B2(n_1292),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1388),
.A2(n_1281),
.B(n_1260),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1388),
.B(n_1326),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1392),
.B(n_1284),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1399),
.B(n_1284),
.C(n_1294),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1397),
.A2(n_1292),
.B1(n_1266),
.B2(n_1275),
.Y(n_1402)
);

AOI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1393),
.A2(n_1260),
.B1(n_1294),
.B2(n_1293),
.C(n_1296),
.Y(n_1403)
);

NAND4xp25_ASAP7_75t_L g1404 ( 
.A(n_1395),
.B(n_1394),
.C(n_1396),
.D(n_1398),
.Y(n_1404)
);

AOI211xp5_ASAP7_75t_L g1405 ( 
.A1(n_1392),
.A2(n_1296),
.B(n_1275),
.C(n_1293),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1392),
.A2(n_1276),
.B(n_1287),
.C(n_1312),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1400),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1404),
.B(n_1311),
.Y(n_1408)
);

AOI321xp33_ASAP7_75t_L g1409 ( 
.A1(n_1401),
.A2(n_1287),
.A3(n_1276),
.B1(n_1234),
.B2(n_1288),
.C(n_1263),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1402),
.Y(n_1410)
);

NOR4xp25_ASAP7_75t_L g1411 ( 
.A(n_1406),
.B(n_1263),
.C(n_1288),
.D(n_1311),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1405),
.Y(n_1412)
);

AOI322xp5_ASAP7_75t_L g1413 ( 
.A1(n_1403),
.A2(n_1287),
.A3(n_1276),
.B1(n_1280),
.B2(n_1285),
.C1(n_1312),
.C2(n_1257),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1400),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1400),
.B(n_1287),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1410),
.B(n_1312),
.Y(n_1416)
);

OAI21xp33_ASAP7_75t_L g1417 ( 
.A1(n_1412),
.A2(n_1276),
.B(n_1280),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1414),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1407),
.B(n_1280),
.Y(n_1419)
);

NOR3x1_ASAP7_75t_L g1420 ( 
.A(n_1408),
.B(n_286),
.C(n_287),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1408),
.B(n_1285),
.Y(n_1421)
);

NAND4xp75_ASAP7_75t_L g1422 ( 
.A(n_1415),
.B(n_1411),
.C(n_1413),
.D(n_1409),
.Y(n_1422)
);

NOR3xp33_ASAP7_75t_L g1423 ( 
.A(n_1414),
.B(n_1285),
.C(n_1257),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1407),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1418),
.Y(n_1425)
);

NOR3xp33_ASAP7_75t_SL g1426 ( 
.A(n_1424),
.B(n_288),
.C(n_289),
.Y(n_1426)
);

NOR4xp25_ASAP7_75t_L g1427 ( 
.A(n_1416),
.B(n_1285),
.C(n_292),
.D(n_293),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1419),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1419),
.B(n_1257),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1422),
.A2(n_290),
.B1(n_296),
.B2(n_297),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1425),
.B(n_1420),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1428),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1430),
.Y(n_1433)
);

XOR2xp5_ASAP7_75t_L g1434 ( 
.A(n_1429),
.B(n_1421),
.Y(n_1434)
);

AOI22x1_ASAP7_75t_L g1435 ( 
.A1(n_1432),
.A2(n_1427),
.B1(n_1426),
.B2(n_1423),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1431),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1436),
.A2(n_1433),
.B1(n_1417),
.B2(n_1434),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1435),
.B(n_300),
.Y(n_1438)
);

OR3x1_ASAP7_75t_L g1439 ( 
.A(n_1437),
.B(n_303),
.C(n_307),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1438),
.B(n_350),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1439),
.B(n_308),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1440),
.A2(n_311),
.B(n_312),
.Y(n_1442)
);

AOI222xp33_ASAP7_75t_L g1443 ( 
.A1(n_1441),
.A2(n_1442),
.B1(n_314),
.B2(n_315),
.C1(n_317),
.C2(n_319),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1443),
.A2(n_1442),
.B1(n_321),
.B2(n_322),
.Y(n_1444)
);

OAI221xp5_ASAP7_75t_R g1445 ( 
.A1(n_1444),
.A2(n_313),
.B1(n_324),
.B2(n_326),
.C(n_328),
.Y(n_1445)
);

AOI211xp5_ASAP7_75t_L g1446 ( 
.A1(n_1445),
.A2(n_329),
.B(n_331),
.C(n_333),
.Y(n_1446)
);


endmodule