module fake_jpeg_86_n_320 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_48),
.B(n_50),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_0),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_1),
.CON(n_50),
.SN(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_30),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_30),
.Y(n_99)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_24),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_60),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_55),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_29),
.B1(n_30),
.B2(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_61),
.A2(n_75),
.B1(n_84),
.B2(n_88),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_18),
.B1(n_35),
.B2(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_36),
.B1(n_49),
.B2(n_31),
.Y(n_112)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_71),
.Y(n_120)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_35),
.B1(n_25),
.B2(n_27),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_38),
.B1(n_22),
.B2(n_20),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_76),
.A2(n_39),
.B1(n_34),
.B2(n_28),
.Y(n_119)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_40),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_25),
.B1(n_27),
.B2(n_37),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_96),
.Y(n_133)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_103),
.B1(n_26),
.B2(n_31),
.Y(n_130)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_49),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_30),
.Y(n_107)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_36),
.Y(n_134)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_19),
.B1(n_39),
.B2(n_34),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_134),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_79),
.C(n_72),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_77),
.C(n_80),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_98),
.B1(n_82),
.B2(n_66),
.Y(n_147)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_62),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_28),
.B1(n_26),
.B2(n_19),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_124),
.Y(n_143)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_81),
.B1(n_23),
.B2(n_36),
.Y(n_161)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_141),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_139),
.B(n_145),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_69),
.B1(n_103),
.B2(n_88),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_147),
.B1(n_113),
.B2(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_63),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_58),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_142),
.B(n_164),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_146),
.C(n_136),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_61),
.C(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_65),
.A3(n_75),
.B1(n_23),
.B2(n_16),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_83),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_162),
.C(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_62),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_134),
.B1(n_108),
.B2(n_132),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_126),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_112),
.A2(n_23),
.B1(n_5),
.B2(n_6),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_23),
.B(n_5),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_3),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_200),
.B1(n_201),
.B2(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_181),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_126),
.B(n_136),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_178),
.A2(n_148),
.B(n_163),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_183),
.C(n_153),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_128),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_184),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_186),
.B1(n_203),
.B2(n_147),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_122),
.B1(n_108),
.B2(n_115),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_197),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_125),
.B(n_132),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_169),
.B(n_152),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_196),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_122),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_125),
.B1(n_137),
.B2(n_127),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_151),
.A2(n_113),
.B1(n_114),
.B2(n_127),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_111),
.B1(n_131),
.B2(n_129),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_206),
.A2(n_218),
.B(n_222),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_212),
.B1(n_189),
.B2(n_197),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_148),
.B1(n_152),
.B2(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_169),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_224),
.C(n_227),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_175),
.A2(n_171),
.B(n_162),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_143),
.B(n_154),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_189),
.B(n_174),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_166),
.B1(n_158),
.B2(n_111),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_226),
.A2(n_229),
.B1(n_186),
.B2(n_202),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_158),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_185),
.A2(n_166),
.B1(n_111),
.B2(n_6),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_15),
.C(n_5),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_182),
.C(n_176),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_222),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_203),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_236),
.B(n_238),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_237),
.B1(n_224),
.B2(n_216),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_235),
.A2(n_246),
.B1(n_220),
.B2(n_215),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_205),
.B(n_200),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_187),
.B1(n_174),
.B2(n_194),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_208),
.B(n_177),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_242),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_247),
.Y(n_263)
);

A2O1A1O1Ixp25_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_195),
.B(n_198),
.C(n_180),
.D(n_188),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_210),
.A2(n_184),
.B1(n_7),
.B2(n_8),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_209),
.B1(n_217),
.B2(n_11),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_3),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_262),
.B1(n_265),
.B2(n_7),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_227),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_11),
.C(n_12),
.Y(n_282)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_266),
.B1(n_250),
.B2(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_210),
.B1(n_229),
.B2(n_226),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_230),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_268),
.C(n_239),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_221),
.B1(n_217),
.B2(n_209),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_217),
.C(n_8),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_231),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_236),
.B1(n_249),
.B2(n_233),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_271),
.A2(n_272),
.B1(n_275),
.B2(n_256),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_233),
.B1(n_231),
.B2(n_239),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_263),
.B(n_243),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_279),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_235),
.B1(n_252),
.B2(n_248),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_266),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_246),
.C(n_11),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_282),
.C(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_275),
.B1(n_278),
.B2(n_274),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_270),
.A2(n_268),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_288),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_270),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_264),
.CI(n_255),
.CON(n_288),
.SN(n_288)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_278),
.C(n_282),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_285),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_258),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_261),
.B1(n_13),
.B2(n_14),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_296),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_307),
.B(n_292),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_300),
.B(n_295),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_311),
.B(n_290),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_284),
.B(n_302),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_306),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_313),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_314),
.B(n_303),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_303),
.B(n_301),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_288),
.B(n_13),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_15),
.C(n_12),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_12),
.B(n_14),
.Y(n_320)
);


endmodule