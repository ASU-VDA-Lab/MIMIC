module fake_jpeg_193_n_682 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_682);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_682;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_650;
wire n_344;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_64),
.Y(n_188)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_66),
.Y(n_191)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_68),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_69),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_70),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_73),
.Y(n_186)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_11),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_78),
.A2(n_84),
.B(n_121),
.Y(n_226)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_80),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_11),
.C(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_83),
.B(n_108),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_11),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_89),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_90),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

CKINVDCx6p67_ASAP7_75t_R g152 ( 
.A(n_94),
.Y(n_152)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_98),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_27),
.B(n_10),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_31),
.B(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_124),
.Y(n_144)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

CKINVDCx6p67_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_132),
.Y(n_174)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_116),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_12),
.B1(n_18),
.B2(n_17),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_29),
.B1(n_25),
.B2(n_41),
.Y(n_161)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_27),
.B(n_8),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_122),
.Y(n_229)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_25),
.B(n_19),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_26),
.Y(n_125)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_39),
.B(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_41),
.Y(n_168)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_31),
.Y(n_128)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_129),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_33),
.A2(n_12),
.B(n_17),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_1),
.Y(n_140)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_32),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_80),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_135),
.B(n_198),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_53),
.B1(n_32),
.B2(n_39),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_139),
.A2(n_146),
.B1(n_150),
.B2(n_154),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_140),
.B(n_168),
.C(n_176),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_78),
.A2(n_53),
.B1(n_39),
.B2(n_26),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_58),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_147),
.B(n_165),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_53),
.B1(n_36),
.B2(n_42),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_42),
.B1(n_36),
.B2(n_54),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_61),
.A2(n_129),
.B1(n_118),
.B2(n_117),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_158),
.A2(n_183),
.B1(n_1),
.B2(n_2),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_79),
.A2(n_42),
.B1(n_36),
.B2(n_54),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_159),
.A2(n_184),
.B1(n_194),
.B2(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_161),
.A2(n_177),
.B1(n_185),
.B2(n_210),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_94),
.A2(n_58),
.A3(n_57),
.B1(n_43),
.B2(n_52),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_163),
.B(n_1),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_62),
.B(n_43),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_57),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_122),
.A2(n_40),
.B1(n_56),
.B2(n_54),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_64),
.A2(n_73),
.B1(n_69),
.B2(n_111),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_81),
.A2(n_42),
.B1(n_36),
.B2(n_54),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_70),
.A2(n_56),
.B1(n_51),
.B2(n_29),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_71),
.A2(n_49),
.B1(n_52),
.B2(n_56),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_189),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_113),
.A2(n_49),
.B(n_59),
.C(n_24),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_192),
.B(n_220),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_81),
.A2(n_56),
.B1(n_59),
.B2(n_24),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_82),
.B(n_40),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_195),
.B(n_196),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_89),
.B(n_59),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_82),
.B(n_40),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_66),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_100),
.A2(n_44),
.B1(n_34),
.B2(n_55),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_91),
.Y(n_214)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_93),
.A2(n_55),
.B1(n_12),
.B2(n_13),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_99),
.B(n_12),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_219),
.B(n_200),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_116),
.B(n_17),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_104),
.Y(n_224)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_105),
.A2(n_55),
.B1(n_7),
.B2(n_14),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_151),
.B(n_103),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_231),
.Y(n_317)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_162),
.B(n_103),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_235),
.B(n_253),
.Y(n_332)
);

INVx3_ASAP7_75t_SL g236 ( 
.A(n_142),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_236),
.Y(n_324)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_237),
.Y(n_316)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_239),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_185),
.A2(n_106),
.B1(n_55),
.B2(n_14),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_240),
.A2(n_271),
.B1(n_204),
.B2(n_202),
.Y(n_318)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_241),
.Y(n_342)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_134),
.Y(n_243)
);

INVx4_ASAP7_75t_SL g353 ( 
.A(n_243),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_152),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_245),
.B(n_281),
.Y(n_315)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_247),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_152),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_248),
.B(n_277),
.Y(n_325)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_157),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_250),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_174),
.A2(n_102),
.B1(n_55),
.B2(n_7),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_252),
.A2(n_257),
.B1(n_261),
.B2(n_273),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_160),
.B(n_102),
.Y(n_253)
);

OA22x2_ASAP7_75t_SL g254 ( 
.A1(n_150),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g327 ( 
.A1(n_254),
.A2(n_312),
.B1(n_145),
.B2(n_223),
.Y(n_327)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_255),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_174),
.A2(n_7),
.B1(n_17),
.B2(n_4),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_258),
.Y(n_361)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_157),
.Y(n_259)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_259),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_171),
.B(n_4),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_260),
.B(n_270),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_138),
.Y(n_262)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_134),
.Y(n_264)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_268),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_199),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_193),
.B(n_4),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_6),
.B1(n_7),
.B2(n_15),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_176),
.A2(n_142),
.B1(n_146),
.B2(n_164),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_274),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_227),
.A2(n_6),
.B1(n_15),
.B2(n_19),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_275),
.A2(n_278),
.B1(n_279),
.B2(n_305),
.Y(n_339)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_178),
.Y(n_276)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_153),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_181),
.A2(n_6),
.B1(n_19),
.B2(n_2),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_167),
.A2(n_2),
.B1(n_172),
.B2(n_136),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_179),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_154),
.A2(n_2),
.B1(n_183),
.B2(n_158),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_282),
.A2(n_217),
.B1(n_188),
.B2(n_209),
.Y(n_348)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_166),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_287),
.Y(n_328)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_137),
.Y(n_286)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_286),
.Y(n_365)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_144),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_288),
.B(n_298),
.Y(n_347)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_289),
.B(n_290),
.Y(n_360)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_148),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_192),
.B(n_149),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_175),
.Y(n_321)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_292),
.B(n_293),
.Y(n_368)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_215),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_159),
.A2(n_184),
.B1(n_139),
.B2(n_194),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_294),
.A2(n_256),
.B1(n_242),
.B2(n_308),
.Y(n_376)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_167),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_173),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_297),
.Y(n_372)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_156),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_300),
.Y(n_337)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_222),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_136),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_304),
.Y(n_352)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_191),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_198),
.A2(n_199),
.B1(n_143),
.B2(n_141),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_169),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_309),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_207),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_191),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_311),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_141),
.Y(n_311)
);

AO22x1_ASAP7_75t_SL g312 ( 
.A1(n_190),
.A2(n_202),
.B1(n_170),
.B2(n_209),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_190),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_314),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_207),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_318),
.B(n_320),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_321),
.A2(n_322),
.B(n_236),
.Y(n_409)
);

OR2x2_ASAP7_75t_SL g322 ( 
.A(n_307),
.B(n_143),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_327),
.B(n_336),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_280),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_351),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g336 ( 
.A(n_244),
.B(n_267),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_294),
.A2(n_221),
.B1(n_223),
.B2(n_170),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_282),
.A2(n_261),
.B1(n_234),
.B2(n_254),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_346),
.A2(n_366),
.B1(n_369),
.B2(n_317),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_348),
.A2(n_375),
.B1(n_376),
.B2(n_292),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_231),
.B(n_155),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_231),
.B(n_155),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_359),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_269),
.B(n_225),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_269),
.B(n_225),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_371),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_254),
.A2(n_221),
.B1(n_170),
.B2(n_212),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_308),
.A2(n_212),
.B1(n_188),
.B2(n_217),
.Y(n_369)
);

CKINVDCx12_ASAP7_75t_R g370 ( 
.A(n_258),
.Y(n_370)
);

INVx3_ASAP7_75t_SL g402 ( 
.A(n_370),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_250),
.B(n_182),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_285),
.B(n_186),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_262),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_284),
.A2(n_186),
.B1(n_197),
.B2(n_246),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_245),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_378),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_375),
.A2(n_284),
.B1(n_308),
.B2(n_312),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_379),
.A2(n_393),
.B1(n_397),
.B2(n_424),
.Y(n_450)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_308),
.C(n_276),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_391),
.C(n_401),
.Y(n_433)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_326),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_389),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_376),
.A2(n_312),
.B1(n_310),
.B2(n_304),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_387),
.A2(n_423),
.B1(n_411),
.B2(n_412),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_352),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_232),
.C(n_286),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_347),
.B(n_290),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_392),
.B(n_400),
.Y(n_452)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_321),
.A2(n_251),
.B1(n_265),
.B2(n_266),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_337),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_406),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_317),
.A2(n_233),
.B1(n_259),
.B2(n_243),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_L g445 ( 
.A1(n_399),
.A2(n_409),
.B(n_388),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_347),
.B(n_299),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_336),
.B(n_322),
.C(n_358),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_320),
.A2(n_264),
.B1(n_293),
.B2(n_289),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_404),
.B1(n_422),
.B2(n_324),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_323),
.Y(n_405)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_332),
.B(n_311),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_241),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_371),
.C(n_350),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_419),
.Y(n_430)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_414),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_338),
.B(n_325),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_421),
.Y(n_443)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_420),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_338),
.B(n_301),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_417),
.B(n_371),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_418),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_359),
.B(n_237),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_362),
.A2(n_274),
.B1(n_249),
.B2(n_297),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_348),
.A2(n_238),
.B1(n_247),
.B2(n_263),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_351),
.A2(n_255),
.B1(n_268),
.B2(n_272),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_327),
.A2(n_333),
.B1(n_372),
.B2(n_364),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_339),
.Y(n_457)
);

BUFx12_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_429),
.A2(n_435),
.B1(n_446),
.B2(n_451),
.Y(n_478)
);

AO22x1_ASAP7_75t_L g432 ( 
.A1(n_408),
.A2(n_388),
.B1(n_387),
.B2(n_377),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_444),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_379),
.A2(n_327),
.B1(n_372),
.B2(n_357),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_417),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_440),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_397),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_433),
.C(n_459),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_445),
.A2(n_457),
.B1(n_396),
.B2(n_416),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_386),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_447),
.B(n_365),
.Y(n_498)
);

AOI32xp33_ASAP7_75t_L g449 ( 
.A1(n_382),
.A2(n_315),
.A3(n_327),
.B1(n_363),
.B2(n_328),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_408),
.A2(n_328),
.B1(n_373),
.B2(n_355),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_389),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_454),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_410),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_329),
.B1(n_373),
.B2(n_353),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_458),
.A2(n_402),
.B1(n_415),
.B2(n_421),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_408),
.A2(n_315),
.B(n_367),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_459),
.A2(n_354),
.B(n_370),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_380),
.A2(n_329),
.B1(n_355),
.B2(n_356),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_462),
.A2(n_390),
.B1(n_384),
.B2(n_413),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_380),
.B(n_365),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_464),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_381),
.B(n_367),
.Y(n_464)
);

AO21x2_ASAP7_75t_L g468 ( 
.A1(n_435),
.A2(n_423),
.B(n_424),
.Y(n_468)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_468),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_454),
.A2(n_388),
.B1(n_385),
.B2(n_395),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_469),
.A2(n_476),
.B1(n_467),
.B2(n_490),
.Y(n_519)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_470),
.Y(n_512)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_437),
.Y(n_471)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_471),
.Y(n_523)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_456),
.Y(n_473)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_473),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_440),
.A2(n_385),
.B1(n_395),
.B2(n_394),
.Y(n_476)
);

OAI21xp33_ASAP7_75t_SL g536 ( 
.A1(n_477),
.A2(n_500),
.B(n_503),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_484),
.C(n_494),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_457),
.A2(n_396),
.B(n_409),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_480),
.A2(n_496),
.B(n_444),
.Y(n_528)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_456),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_481),
.Y(n_517)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_448),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_433),
.B(n_401),
.C(n_391),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_453),
.B(n_407),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_485),
.B(n_432),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_448),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_486),
.B(n_489),
.Y(n_518)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_488),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_491),
.A2(n_431),
.B1(n_437),
.B2(n_441),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_450),
.A2(n_419),
.B1(n_420),
.B2(n_418),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_492),
.A2(n_429),
.B1(n_451),
.B2(n_461),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_465),
.B(n_402),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_498),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_340),
.C(n_349),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_443),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_497),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_457),
.A2(n_450),
.B(n_458),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_349),
.C(n_335),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_502),
.C(n_441),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_443),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_434),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_436),
.B(n_335),
.C(n_342),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_438),
.A2(n_418),
.B1(n_405),
.B2(n_383),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_426),
.B(n_354),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_504),
.B(n_324),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_507),
.A2(n_508),
.B1(n_514),
.B2(n_539),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_483),
.A2(n_436),
.B1(n_430),
.B2(n_449),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_427),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_509),
.B(n_510),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_483),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_511),
.B(n_522),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_427),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_513),
.B(n_515),
.C(n_516),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_483),
.A2(n_430),
.B1(n_432),
.B2(n_466),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_464),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_434),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_519),
.B(n_467),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_487),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g524 ( 
.A(n_487),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_524),
.B(n_531),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_525),
.B(n_532),
.C(n_499),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_527),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_528),
.A2(n_480),
.B(n_500),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_426),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_475),
.B(n_476),
.C(n_469),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_478),
.A2(n_462),
.B1(n_466),
.B2(n_461),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_534),
.A2(n_540),
.B1(n_468),
.B2(n_495),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_537),
.A2(n_468),
.B1(n_492),
.B2(n_496),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_501),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_538),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_468),
.A2(n_441),
.B1(n_431),
.B2(n_460),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_468),
.A2(n_452),
.B1(n_441),
.B2(n_460),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_490),
.B(n_452),
.Y(n_541)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_541),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_542),
.B(n_550),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_547),
.A2(n_563),
.B(n_569),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_548),
.A2(n_573),
.B1(n_539),
.B2(n_507),
.Y(n_577)
);

NOR3xp33_ASAP7_75t_SL g550 ( 
.A(n_541),
.B(n_470),
.C(n_472),
.Y(n_550)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_551),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_571),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_473),
.Y(n_553)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_553),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_505),
.B(n_481),
.Y(n_555)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_555),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_508),
.A2(n_474),
.B1(n_486),
.B2(n_497),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_556),
.A2(n_560),
.B1(n_565),
.B2(n_568),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_530),
.B(n_486),
.Y(n_558)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_558),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_502),
.Y(n_559)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_559),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_517),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_562),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_528),
.A2(n_488),
.B(n_482),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_521),
.Y(n_564)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_564),
.Y(n_590)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_533),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_519),
.B(n_474),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_566),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_514),
.B(n_526),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_567),
.Y(n_586)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_533),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_512),
.B(n_471),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_489),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_529),
.B(n_405),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_537),
.Y(n_583)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_535),
.Y(n_573)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_577),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_SL g580 ( 
.A(n_570),
.B(n_515),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_580),
.B(n_588),
.Y(n_609)
);

FAx1_ASAP7_75t_SL g581 ( 
.A(n_561),
.B(n_532),
.CI(n_510),
.CON(n_581),
.SN(n_581)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_581),
.B(n_593),
.Y(n_608)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_583),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_570),
.B(n_509),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_552),
.B(n_506),
.C(n_513),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_543),
.C(n_559),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_551),
.A2(n_520),
.B1(n_540),
.B2(n_536),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_592),
.A2(n_594),
.B1(n_595),
.B2(n_549),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_SL g593 ( 
.A1(n_548),
.A2(n_520),
.B(n_518),
.C(n_535),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_562),
.A2(n_534),
.B1(n_516),
.B2(n_525),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_564),
.A2(n_506),
.B1(n_523),
.B2(n_329),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_549),
.A2(n_523),
.B1(n_341),
.B2(n_428),
.Y(n_596)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_596),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_SL g597 ( 
.A(n_543),
.B(n_428),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_563),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_589),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_599),
.B(n_601),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_600),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_589),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_556),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_603),
.B(n_610),
.Y(n_627)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_578),
.Y(n_605)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_605),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_575),
.A2(n_546),
.B(n_547),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_606),
.A2(n_617),
.B(n_583),
.Y(n_623)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_611),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_582),
.B(n_555),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_612),
.B(n_616),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_566),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_613),
.B(n_618),
.C(n_588),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_598),
.B(n_560),
.Y(n_614)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_614),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_615),
.A2(n_576),
.B1(n_596),
.B2(n_567),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_582),
.B(n_542),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_575),
.A2(n_592),
.B(n_587),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_595),
.B(n_568),
.C(n_565),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_586),
.B(n_544),
.Y(n_619)
);

OAI321xp33_ASAP7_75t_L g621 ( 
.A1(n_619),
.A2(n_611),
.A3(n_561),
.B1(n_585),
.B2(n_590),
.C(n_554),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_619),
.A2(n_545),
.B1(n_544),
.B2(n_587),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_620),
.B(n_629),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_621),
.A2(n_631),
.B(n_633),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_623),
.B(n_626),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_625),
.B(n_603),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_600),
.B(n_584),
.C(n_594),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_602),
.A2(n_579),
.B1(n_554),
.B2(n_577),
.Y(n_630)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_630),
.Y(n_646)
);

OAI321xp33_ASAP7_75t_L g631 ( 
.A1(n_614),
.A2(n_545),
.A3(n_550),
.B1(n_553),
.B2(n_571),
.C(n_558),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_580),
.C(n_557),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_632),
.B(n_616),
.C(n_613),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_606),
.A2(n_593),
.B(n_557),
.Y(n_633)
);

FAx1_ASAP7_75t_SL g635 ( 
.A(n_608),
.B(n_581),
.CI(n_593),
.CON(n_635),
.SN(n_635)
);

AOI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_635),
.A2(n_608),
.B1(n_604),
.B2(n_581),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_638),
.B(n_649),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_639),
.B(n_642),
.Y(n_657)
);

AO21x1_ASAP7_75t_L g654 ( 
.A1(n_640),
.A2(n_645),
.B(n_637),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_629),
.B(n_614),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_641),
.B(n_647),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g642 ( 
.A(n_633),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_636),
.B(n_602),
.C(n_607),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_643),
.B(n_644),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_622),
.B(n_617),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_607),
.C(n_610),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_625),
.B(n_609),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_623),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_651),
.B(n_652),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_627),
.B(n_626),
.C(n_630),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_SL g670 ( 
.A1(n_654),
.A2(n_660),
.B(n_428),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_650),
.A2(n_628),
.B1(n_624),
.B2(n_593),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_656),
.B(n_662),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_650),
.A2(n_635),
.B(n_634),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_646),
.A2(n_635),
.B(n_627),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_661),
.A2(n_640),
.B(n_647),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_648),
.A2(n_573),
.B1(n_569),
.B2(n_572),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_643),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_663),
.B(n_341),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g664 ( 
.A(n_655),
.B(n_638),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_664),
.B(n_668),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_659),
.B(n_652),
.Y(n_665)
);

NAND3xp33_ASAP7_75t_SL g672 ( 
.A(n_665),
.B(n_667),
.C(n_669),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_653),
.A2(n_639),
.B1(n_649),
.B2(n_609),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_670),
.A2(n_661),
.B(n_660),
.Y(n_674)
);

OAI21xp33_ASAP7_75t_L g671 ( 
.A1(n_666),
.A2(n_657),
.B(n_654),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_671),
.B(n_674),
.C(n_655),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_673),
.B(n_665),
.C(n_658),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_675),
.A2(n_676),
.B(n_672),
.Y(n_677)
);

AOI322xp5_ASAP7_75t_L g678 ( 
.A1(n_677),
.A2(n_361),
.A3(n_330),
.B1(n_324),
.B2(n_345),
.C1(n_342),
.C2(n_319),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_678),
.B(n_330),
.C(n_345),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_SL g680 ( 
.A1(n_679),
.A2(n_361),
.B(n_319),
.C(n_316),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_680),
.A2(n_361),
.B1(n_344),
.B2(n_316),
.Y(n_681)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_681),
.B(n_344),
.Y(n_682)
);


endmodule