module fake_jpeg_30739_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_20),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_1),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_59),
.B(n_74),
.Y(n_166)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_63),
.Y(n_127)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_31),
.B(n_1),
.CON(n_74),
.SN(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_1),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_95),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_23),
.B(n_2),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_51),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_3),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_25),
.B(n_4),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_106),
.Y(n_153)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_4),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_36),
.C(n_26),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_28),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_111),
.B(n_128),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_46),
.B1(n_32),
.B2(n_34),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_115),
.A2(n_140),
.B1(n_27),
.B2(n_26),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_67),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_59),
.B(n_28),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_142),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_56),
.A2(n_46),
.B1(n_32),
.B2(n_34),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_58),
.B(n_42),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_84),
.B(n_42),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_48),
.Y(n_184)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_54),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_74),
.B1(n_48),
.B2(n_43),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_174),
.Y(n_260)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_176),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_63),
.B(n_36),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_177),
.A2(n_153),
.B(n_50),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_178),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_43),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_179),
.B(n_214),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_184),
.B(n_201),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_109),
.A2(n_105),
.B1(n_107),
.B2(n_71),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_188),
.A2(n_212),
.B1(n_218),
.B2(n_224),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_189),
.Y(n_264)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_57),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_191),
.B(n_197),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_193),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_130),
.A2(n_86),
.B1(n_83),
.B2(n_76),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_194),
.A2(n_208),
.B1(n_227),
.B2(n_228),
.Y(n_265)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_120),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_199),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_49),
.C(n_27),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_127),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_114),
.B(n_33),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_202),
.B(n_217),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_124),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_213),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_135),
.A2(n_60),
.B1(n_75),
.B2(n_58),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_155),
.A2(n_99),
.B1(n_69),
.B2(n_102),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_125),
.B(n_37),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_216),
.Y(n_242)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_136),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_118),
.A2(n_98),
.B1(n_92),
.B2(n_90),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_220),
.Y(n_255)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_108),
.B(n_33),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_49),
.Y(n_235)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_108),
.B(n_22),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_155),
.A2(n_87),
.B1(n_78),
.B2(n_72),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_129),
.Y(n_275)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_115),
.A2(n_68),
.B1(n_66),
.B2(n_61),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_146),
.A2(n_70),
.B1(n_46),
.B2(n_34),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_230),
.A2(n_165),
.B1(n_150),
.B2(n_123),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_161),
.B1(n_147),
.B2(n_163),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_232),
.A2(n_237),
.B1(n_224),
.B2(n_245),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_127),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_234),
.A2(n_238),
.B(n_75),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_235),
.B(n_204),
.C(n_5),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_161),
.B1(n_147),
.B2(n_156),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_188),
.A2(n_146),
.B1(n_165),
.B2(n_152),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_243),
.A2(n_277),
.B1(n_164),
.B2(n_172),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_140),
.B1(n_152),
.B2(n_150),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_245),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_201),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_131),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_170),
.B(n_154),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_22),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_266),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_198),
.B(n_50),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_203),
.B(n_37),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_271),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_180),
.B(n_153),
.C(n_129),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_276),
.C(n_196),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_191),
.B(n_202),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_194),
.A2(n_208),
.B(n_205),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

BUFx16f_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_282),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_206),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_283),
.B(n_296),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_286),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_241),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_123),
.B1(n_156),
.B2(n_164),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_304),
.B1(n_239),
.B2(n_277),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_197),
.B1(n_215),
.B2(n_211),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_212),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_249),
.C(n_259),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_240),
.B(n_193),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_185),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_234),
.B(n_192),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_254),
.B(n_271),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_298),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_181),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_182),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_307),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_242),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_303),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_181),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_238),
.A2(n_29),
.B(n_216),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_305),
.A2(n_279),
.B(n_272),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_306),
.B(n_276),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_53),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_263),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_312),
.Y(n_355)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_255),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_268),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_288),
.Y(n_330)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_320),
.Y(n_341)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_204),
.Y(n_315)
);

AOI32xp33_ASAP7_75t_L g338 ( 
.A1(n_315),
.A2(n_249),
.A3(n_270),
.B1(n_274),
.B2(n_267),
.Y(n_338)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_316),
.Y(n_334)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_233),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_317),
.A2(n_322),
.B1(n_256),
.B2(n_264),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_29),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_318),
.Y(n_342)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_261),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_319),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_257),
.B(n_53),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_272),
.B(n_270),
.Y(n_326)
);

CKINVDCx12_ASAP7_75t_R g322 ( 
.A(n_263),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_290),
.B1(n_292),
.B2(n_313),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_323),
.A2(n_324),
.B1(n_347),
.B2(n_349),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_309),
.A2(n_243),
.B1(n_239),
.B2(n_245),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_325),
.A2(n_357),
.B1(n_337),
.B2(n_359),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_326),
.B(n_339),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_SL g392 ( 
.A(n_327),
.B(n_338),
.C(n_319),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_279),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_353),
.C(n_358),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_343),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_331),
.A2(n_351),
.B(n_333),
.C(n_327),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_306),
.A2(n_279),
.B(n_274),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_333),
.A2(n_351),
.B(n_289),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_280),
.B(n_273),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_311),
.A2(n_245),
.B1(n_189),
.B2(n_126),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_287),
.A2(n_126),
.B1(n_256),
.B2(n_267),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_305),
.A2(n_236),
.B(n_278),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_304),
.A2(n_278),
.B1(n_264),
.B2(n_259),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_357),
.A2(n_359),
.B1(n_322),
.B2(n_284),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_258),
.C(n_251),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_291),
.A2(n_258),
.B1(n_251),
.B2(n_149),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_288),
.B(n_53),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_282),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_332),
.B(n_299),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_362),
.B(n_369),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_363),
.A2(n_377),
.B1(n_381),
.B2(n_396),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_315),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_366),
.Y(n_400)
);

AO21x1_ASAP7_75t_L g406 ( 
.A1(n_365),
.A2(n_392),
.B(n_393),
.Y(n_406)
);

AOI32xp33_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_303),
.A3(n_298),
.B1(n_296),
.B2(n_302),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_332),
.B(n_297),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_330),
.B(n_286),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_372),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_348),
.C(n_343),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_371),
.B(n_337),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_301),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_373),
.A2(n_344),
.B(n_334),
.Y(n_427)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_334),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_345),
.B(n_312),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_379),
.B(n_344),
.Y(n_426)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_325),
.A2(n_284),
.B1(n_283),
.B2(n_320),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_307),
.C(n_314),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_367),
.C(n_353),
.Y(n_405)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_282),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_387),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_319),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_354),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_388),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_330),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_390),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_354),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_336),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_336),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_331),
.B(n_300),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_329),
.A2(n_324),
.B1(n_323),
.B2(n_347),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_367),
.B(n_327),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_407),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_341),
.Y(n_403)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_412),
.C(n_415),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_335),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_341),
.Y(n_409)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_335),
.Y(n_410)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_410),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_346),
.C(n_342),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_342),
.C(n_361),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_416),
.B(n_365),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_294),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_373),
.A2(n_337),
.B(n_338),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_418),
.A2(n_427),
.B(n_365),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_316),
.Y(n_420)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_316),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_423),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_337),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_425),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_349),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_426),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_427),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_445),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_402),
.A2(n_384),
.B1(n_364),
.B2(n_385),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_432),
.A2(n_426),
.B1(n_408),
.B2(n_421),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_393),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_433),
.A2(n_436),
.B(n_439),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_434),
.B(n_450),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_402),
.A2(n_384),
.B1(n_395),
.B2(n_368),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_443),
.B1(n_449),
.B2(n_428),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_365),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_441),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_406),
.A2(n_365),
.B(n_378),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_377),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_404),
.A2(n_394),
.B1(n_375),
.B2(n_380),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_376),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_456),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_424),
.A2(n_390),
.B1(n_388),
.B2(n_383),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_446),
.A2(n_442),
.B1(n_431),
.B2(n_421),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_356),
.Y(n_447)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_448),
.B(n_452),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_404),
.A2(n_317),
.B1(n_310),
.B2(n_46),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_416),
.B(n_149),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_401),
.B(n_4),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_415),
.B(n_137),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_400),
.C(n_412),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_465),
.C(n_466),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_406),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_462),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_433),
.B1(n_440),
.B2(n_436),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_406),
.C(n_409),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_425),
.C(n_398),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_398),
.C(n_418),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_467),
.A2(n_468),
.B1(n_473),
.B2(n_474),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_432),
.A2(n_428),
.B1(n_422),
.B2(n_419),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_403),
.C(n_422),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_477),
.C(n_434),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_455),
.A2(n_453),
.B1(n_454),
.B2(n_429),
.Y(n_470)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_413),
.C(n_419),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_479),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_447),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_472),
.B(n_476),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_441),
.A2(n_397),
.B1(n_411),
.B2(n_413),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_397),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_413),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_475),
.Y(n_480)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_480),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_439),
.B1(n_446),
.B2(n_433),
.Y(n_486)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_488),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_460),
.B(n_479),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_489),
.B(n_464),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_490),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_29),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_459),
.A2(n_478),
.B1(n_466),
.B2(n_465),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_496),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_450),
.C(n_411),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_497),
.C(n_53),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_458),
.A2(n_137),
.B1(n_136),
.B2(n_122),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_495),
.A2(n_469),
.B1(n_464),
.B2(n_458),
.Y(n_501)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_462),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_463),
.B(n_45),
.C(n_126),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_513),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_494),
.B1(n_495),
.B2(n_8),
.Y(n_524)
);

INVx6_ASAP7_75t_L g502 ( 
.A(n_481),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_511),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_484),
.A2(n_480),
.B1(n_492),
.B2(n_487),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_505),
.A2(n_506),
.B1(n_512),
.B2(n_488),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_485),
.A2(n_477),
.B1(n_122),
.B2(n_7),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_73),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_509),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_29),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_483),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_499),
.B(n_502),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_518),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_482),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_521),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_504),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_510),
.A2(n_489),
.B(n_491),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_522),
.A2(n_513),
.B1(n_9),
.B2(n_10),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_507),
.B(n_497),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_525),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_524),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_506),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_503),
.B(n_53),
.C(n_7),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_6),
.Y(n_533)
);

OAI21xp33_ASAP7_75t_L g530 ( 
.A1(n_516),
.A2(n_512),
.B(n_509),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_530),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_526),
.C(n_525),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_533),
.B(n_535),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_519),
.B(n_6),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_537),
.B(n_540),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_529),
.B(n_528),
.C(n_527),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_538),
.A2(n_53),
.B(n_11),
.Y(n_544)
);

NOR2x1_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_517),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_519),
.C(n_514),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_541),
.A2(n_530),
.B(n_514),
.Y(n_542)
);

AOI322xp5_ASAP7_75t_L g546 ( 
.A1(n_542),
.A2(n_544),
.A3(n_536),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_16),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_543),
.B(n_539),
.Y(n_545)
);

O2A1O1Ixp33_ASAP7_75t_L g547 ( 
.A1(n_545),
.A2(n_546),
.B(n_536),
.C(n_12),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_9),
.C(n_12),
.Y(n_548)
);

AO21x1_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_9),
.B(n_13),
.Y(n_549)
);

MAJx2_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_13),
.C(n_14),
.Y(n_550)
);

O2A1O1Ixp33_ASAP7_75t_SL g551 ( 
.A1(n_550),
.A2(n_14),
.B(n_16),
.C(n_549),
.Y(n_551)
);


endmodule