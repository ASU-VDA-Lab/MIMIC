module fake_jpeg_2825_n_192 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_22),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_2),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_76),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_4),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_66),
.Y(n_90)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_50),
.B1(n_62),
.B2(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_89),
.B1(n_56),
.B2(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_51),
.B1(n_66),
.B2(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_56),
.B1(n_49),
.B2(n_59),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_99),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_89),
.B1(n_65),
.B2(n_62),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_58),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_107),
.Y(n_122)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_53),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_49),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_124),
.B1(n_128),
.B2(n_5),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_57),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_86),
.B(n_57),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_121),
.B(n_6),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_86),
.B(n_69),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_61),
.B1(n_68),
.B2(n_54),
.Y(n_124)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_4),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_131),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_25),
.B1(n_45),
.B2(n_44),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_135),
.B1(n_137),
.B2(n_113),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_7),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_23),
.B1(n_41),
.B2(n_36),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_121),
.B1(n_120),
.B2(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_8),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_143),
.B(n_149),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_48),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_35),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_34),
.C(n_31),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_30),
.C(n_29),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_8),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_148),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_9),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_157),
.B1(n_13),
.B2(n_15),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_146),
.C(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_28),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_27),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_161),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_19),
.B(n_12),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_165),
.B(n_147),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_11),
.B(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_175),
.B1(n_165),
.B2(n_157),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_145),
.C(n_134),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_155),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_145),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_156),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_144),
.B1(n_132),
.B2(n_16),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_158),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_179),
.C(n_181),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_180),
.B1(n_171),
.B2(n_173),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_166),
.A3(n_163),
.B1(n_151),
.B2(n_162),
.C(n_159),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_172),
.B(n_170),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_184),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

AOI21x1_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_154),
.B(n_16),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_182),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_187),
.B(n_183),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_13),
.B(n_17),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_17),
.C(n_18),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_18),
.Y(n_192)
);


endmodule