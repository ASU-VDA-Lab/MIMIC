module fake_jpeg_14439_n_590 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_590);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_590;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_7),
.B(n_14),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_65),
.Y(n_115)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_63),
.A2(n_46),
.B1(n_53),
.B2(n_29),
.Y(n_159)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_67),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_79),
.Y(n_134)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_77),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

NAND2x1_ASAP7_75t_SL g81 ( 
.A(n_30),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_81),
.B(n_87),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_16),
.Y(n_87)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_16),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_90),
.B(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_37),
.B(n_16),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_0),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_93),
.B(n_98),
.Y(n_167)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_23),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_37),
.B(n_0),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_111),
.Y(n_177)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_23),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_38),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_122),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_60),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_118),
.B(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_99),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_61),
.B(n_35),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_70),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_123),
.B(n_149),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_60),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_35),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_160),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_32),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_88),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_153),
.B(n_157),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_62),
.B(n_21),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_39),
.B1(n_29),
.B2(n_52),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_81),
.B(n_53),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_77),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_166),
.B(n_97),
.Y(n_235)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_68),
.B(n_46),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_99),
.Y(n_202)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_180),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_67),
.B1(n_82),
.B2(n_41),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_181),
.A2(n_51),
.B(n_45),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g266 ( 
.A(n_186),
.Y(n_266)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

BUFx2_ASAP7_75t_SL g252 ( 
.A(n_188),
.Y(n_252)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_190),
.B(n_198),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx3_ASAP7_75t_SL g286 ( 
.A(n_192),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_115),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_209),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_195),
.A2(n_234),
.B1(n_27),
.B2(n_25),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_124),
.A2(n_33),
.B1(n_75),
.B2(n_71),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_196),
.A2(n_229),
.B1(n_170),
.B2(n_119),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_SL g197 ( 
.A(n_161),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_197),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_111),
.Y(n_198)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_202),
.B(n_205),
.Y(n_264)
);

CKINVDCx12_ASAP7_75t_R g203 ( 
.A(n_161),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_203),
.Y(n_294)
);

CKINVDCx12_ASAP7_75t_R g204 ( 
.A(n_135),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_204),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_134),
.B(n_39),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_175),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_115),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_111),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

CKINVDCx12_ASAP7_75t_R g213 ( 
.A(n_133),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_214),
.Y(n_271)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_27),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_236),
.Y(n_273)
);

CKINVDCx12_ASAP7_75t_R g222 ( 
.A(n_139),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_126),
.Y(n_227)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_227),
.Y(n_291)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_154),
.A2(n_33),
.B1(n_57),
.B2(n_97),
.Y(n_229)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_231),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_134),
.B(n_52),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_232),
.B(n_117),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_177),
.A2(n_109),
.B1(n_103),
.B2(n_101),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_128),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_152),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_240),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_125),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_131),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_181),
.B1(n_229),
.B2(n_172),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_132),
.Y(n_242)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_144),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_113),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_196),
.A2(n_177),
.B1(n_131),
.B2(n_152),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_253),
.A2(n_254),
.B1(n_156),
.B2(n_199),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_193),
.B(n_176),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_261),
.A2(n_295),
.B(n_241),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_283),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_183),
.B(n_127),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_276),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_274),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_208),
.B(n_148),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_278),
.A2(n_298),
.B1(n_197),
.B2(n_180),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_230),
.B(n_113),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_216),
.B(n_162),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_292),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_216),
.B(n_140),
.C(n_141),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_274),
.C(n_260),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_200),
.B(n_145),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_234),
.A2(n_113),
.B1(n_145),
.B2(n_44),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_188),
.A2(n_172),
.B1(n_156),
.B2(n_45),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_302),
.B(n_318),
.C(n_313),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_304),
.A2(n_282),
.B1(n_262),
.B2(n_256),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_187),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_305),
.B(n_306),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_185),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_309),
.A2(n_345),
.B1(n_284),
.B2(n_286),
.Y(n_359)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_310),
.Y(n_370)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_184),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_319),
.Y(n_357)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_224),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_323),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_182),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_317),
.B(n_320),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_207),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_325),
.Y(n_355)
);

AND2x6_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_128),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_227),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_243),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_321),
.B(n_322),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_206),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_201),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_246),
.B(n_215),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_329),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_257),
.B(n_231),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_326),
.B(n_328),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_290),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_330),
.C(n_339),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_257),
.B(n_214),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_225),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_217),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_189),
.B(n_212),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_331),
.A2(n_343),
.B(n_251),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_281),
.A2(n_132),
.B1(n_136),
.B2(n_146),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_347),
.B1(n_263),
.B2(n_266),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_270),
.B(n_214),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_333),
.B(n_337),
.Y(n_374)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_334),
.Y(n_394)
);

BUFx12f_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

BUFx8_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_191),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_250),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_344),
.Y(n_368)
);

CKINVDCx12_ASAP7_75t_R g339 ( 
.A(n_274),
.Y(n_339)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_248),
.Y(n_341)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_248),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_350),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_287),
.A2(n_51),
.B(n_220),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_263),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_249),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_349),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_249),
.A2(n_136),
.B1(n_146),
.B2(n_86),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_247),
.B(n_226),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_348),
.B(n_297),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g349 ( 
.A(n_252),
.B(n_51),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_301),
.A2(n_282),
.B1(n_286),
.B2(n_266),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_364),
.B1(n_369),
.B2(n_377),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_301),
.B(n_284),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_361),
.C(n_367),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_339),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_308),
.A2(n_262),
.B1(n_299),
.B2(n_256),
.Y(n_366)
);

OA22x2_ASAP7_75t_L g419 ( 
.A1(n_366),
.A2(n_385),
.B1(n_344),
.B2(n_311),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_293),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_316),
.A2(n_299),
.B1(n_192),
.B2(n_186),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_343),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_318),
.B(n_251),
.C(n_291),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_376),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_305),
.B(n_293),
.C(n_291),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_308),
.A2(n_242),
.B1(n_238),
.B2(n_78),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_306),
.B(n_297),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_391),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_308),
.A2(n_331),
.B1(n_323),
.B2(n_330),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_382),
.A2(n_383),
.B1(n_390),
.B2(n_347),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_303),
.A2(n_25),
.B1(n_50),
.B2(n_55),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_332),
.A2(n_84),
.B1(n_73),
.B2(n_247),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_387),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_319),
.A2(n_25),
.B1(n_233),
.B2(n_226),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_313),
.B(n_269),
.C(n_271),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_315),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_395),
.B(n_400),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_SL g441 ( 
.A1(n_396),
.A2(n_394),
.B(n_365),
.Y(n_441)
);

OAI32xp33_ASAP7_75t_L g398 ( 
.A1(n_371),
.A2(n_324),
.A3(n_329),
.B1(n_349),
.B2(n_325),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_415),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_338),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_335),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_401),
.B(n_410),
.Y(n_447)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_368),
.Y(n_402)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_404),
.A2(n_424),
.B1(n_425),
.B2(n_431),
.Y(n_466)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_389),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_414),
.A2(n_372),
.B(n_390),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_358),
.B(n_350),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_416),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_341),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_419),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_363),
.B(n_342),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_421),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_300),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_374),
.B(n_346),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_428),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_382),
.A2(n_312),
.B1(n_340),
.B2(n_345),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_371),
.A2(n_314),
.B1(n_269),
.B2(n_275),
.Y(n_425)
);

INVx13_ASAP7_75t_L g426 ( 
.A(n_370),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_426),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_310),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_429),
.Y(n_461)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_307),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_430),
.B(n_394),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_355),
.A2(n_275),
.B1(n_336),
.B2(n_55),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_386),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_335),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_367),
.C(n_361),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_406),
.C(n_425),
.Y(n_472)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_403),
.B(n_353),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_442),
.B(n_449),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_355),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_445),
.Y(n_478)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_355),
.Y(n_445)
);

AOI21xp33_ASAP7_75t_L g477 ( 
.A1(n_448),
.A2(n_452),
.B(n_419),
.Y(n_477)
);

XNOR2x1_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_373),
.Y(n_449)
);

NOR4xp25_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_357),
.C(n_378),
.D(n_376),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_455),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_420),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_377),
.B(n_380),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_456),
.B(n_465),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_424),
.A2(n_354),
.B1(n_366),
.B2(n_385),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_397),
.B1(n_407),
.B2(n_417),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_414),
.A2(n_380),
.B(n_375),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_460),
.A2(n_334),
.B(n_362),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_397),
.A2(n_351),
.B1(n_392),
.B2(n_375),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_462),
.A2(n_399),
.B1(n_409),
.B2(n_419),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_392),
.Y(n_463)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_463),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_415),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_468),
.A2(n_479),
.B1(n_487),
.B2(n_464),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_473),
.C(n_480),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_431),
.C(n_404),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_474),
.A2(n_482),
.B1(n_484),
.B2(n_490),
.Y(n_499)
);

A2O1A1O1Ixp25_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_398),
.B(n_427),
.C(n_409),
.D(n_426),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_476),
.A2(n_451),
.B(n_434),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_477),
.B(n_486),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_466),
.A2(n_419),
.B1(n_399),
.B2(n_416),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_443),
.C(n_445),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_440),
.A2(n_423),
.B1(n_408),
.B2(n_432),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_335),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_488),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_440),
.A2(n_233),
.B1(n_240),
.B2(n_336),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_51),
.C(n_240),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_492),
.C(n_446),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_439),
.B(n_336),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_459),
.A2(n_55),
.B1(n_50),
.B2(n_44),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_44),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_461),
.A2(n_0),
.B(n_1),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_489),
.B(n_494),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_465),
.A2(n_50),
.B1(n_41),
.B2(n_28),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_447),
.B(n_457),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_450),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_49),
.C(n_41),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_463),
.Y(n_494)
);

NAND2x1_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_0),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_495),
.A2(n_433),
.B(n_435),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_471),
.A2(n_437),
.B1(n_438),
.B2(n_462),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_496),
.A2(n_509),
.B1(n_484),
.B2(n_490),
.Y(n_525)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_472),
.B(n_457),
.CI(n_448),
.CON(n_500),
.SN(n_500)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_500),
.B(n_504),
.Y(n_521)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_437),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_510),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_474),
.A2(n_456),
.B1(n_438),
.B2(n_444),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_506),
.A2(n_511),
.B1(n_479),
.B2(n_495),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_508),
.B(n_513),
.Y(n_537)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_482),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_475),
.A2(n_433),
.B1(n_446),
.B2(n_464),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_518),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_469),
.B(n_454),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_454),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_514),
.B(n_516),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_478),
.Y(n_522)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_480),
.B(n_450),
.C(n_435),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_478),
.C(n_492),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_435),
.Y(n_518)
);

FAx1_ASAP7_75t_SL g519 ( 
.A(n_470),
.B(n_2),
.CI(n_3),
.CON(n_519),
.SN(n_519)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_519),
.A2(n_473),
.B1(n_476),
.B2(n_495),
.Y(n_526)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_520),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_522),
.B(n_499),
.Y(n_551)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_508),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_523),
.B(n_528),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_525),
.A2(n_531),
.B1(n_512),
.B2(n_501),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_526),
.A2(n_533),
.B1(n_524),
.B2(n_527),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_499),
.A2(n_487),
.B1(n_488),
.B2(n_485),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_529),
.B(n_507),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_470),
.C(n_483),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_530),
.B(n_534),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_509),
.A2(n_28),
.B1(n_22),
.B2(n_5),
.Y(n_531)
);

OA21x2_ASAP7_75t_SL g532 ( 
.A1(n_505),
.A2(n_28),
.B(n_23),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_532),
.B(n_511),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_3),
.C(n_4),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_497),
.B(n_4),
.C(n_5),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_536),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_507),
.B(n_515),
.C(n_498),
.Y(n_536)
);

MAJx2_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_500),
.C(n_498),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_539),
.B(n_530),
.C(n_526),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_540),
.B(n_543),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_542),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_510),
.C(n_506),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_523),
.A2(n_501),
.B(n_518),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_545),
.A2(n_533),
.B(n_524),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_546),
.A2(n_549),
.B1(n_552),
.B2(n_527),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_537),
.B(n_502),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_550),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_504),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g567 ( 
.A(n_551),
.B(n_555),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_525),
.A2(n_500),
.B1(n_519),
.B2(n_8),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_554),
.B(n_4),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_522),
.B(n_519),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_556),
.A2(n_558),
.B(n_565),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_557),
.B(n_550),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_542),
.A2(n_534),
.B(n_535),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_559),
.A2(n_564),
.B1(n_9),
.B2(n_10),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_553),
.A2(n_531),
.B1(n_6),
.B2(n_8),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_552),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_551),
.B(n_555),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_546),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_547),
.A2(n_4),
.B(n_6),
.Y(n_565)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_568),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_569),
.B(n_572),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_561),
.A2(n_541),
.B1(n_545),
.B2(n_543),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_570),
.A2(n_573),
.B1(n_575),
.B2(n_564),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_563),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_562),
.B(n_544),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_539),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_576),
.B(n_577),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_574),
.B(n_567),
.C(n_564),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_579),
.B(n_575),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_582),
.B(n_583),
.C(n_581),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_578),
.B(n_564),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_584),
.Y(n_586)
);

AOI322xp5_ASAP7_75t_L g585 ( 
.A1(n_583),
.A2(n_580),
.A3(n_579),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_11),
.Y(n_585)
);

INVxp33_ASAP7_75t_L g587 ( 
.A(n_586),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_585),
.Y(n_588)
);

OAI221xp5_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_589),
.A2(n_10),
.B(n_12),
.Y(n_590)
);


endmodule