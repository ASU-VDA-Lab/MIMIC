module fake_jpeg_492_n_609 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_609);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_609;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_82),
.Y(n_136)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_61),
.Y(n_192)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_62),
.Y(n_150)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_64),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_65),
.B(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_67),
.B(n_70),
.Y(n_153)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_71),
.B(n_74),
.Y(n_154)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_73),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_19),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_76),
.Y(n_156)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_84),
.Y(n_221)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_18),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_90),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_45),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_100),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_43),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_97),
.B(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_25),
.B(n_1),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_17),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_33),
.B(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_27),
.B(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_118),
.B(n_124),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_33),
.B(n_2),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_120),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_37),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_56),
.B(n_28),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_51),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_128),
.Y(n_180)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_27),
.B(n_2),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_59),
.B1(n_78),
.B2(n_85),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_129),
.A2(n_146),
.B1(n_158),
.B2(n_163),
.Y(n_272)
);

OR2x4_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_40),
.Y(n_131)
);

OR2x2_ASAP7_75t_SL g252 ( 
.A(n_131),
.B(n_10),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_116),
.B1(n_51),
.B2(n_114),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_144),
.A2(n_174),
.B1(n_178),
.B2(n_158),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_53),
.B1(n_50),
.B2(n_48),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_58),
.A2(n_50),
.B1(n_48),
.B2(n_44),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_84),
.A2(n_52),
.B1(n_46),
.B2(n_30),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_80),
.A2(n_87),
.B1(n_125),
.B2(n_46),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_60),
.Y(n_175)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_91),
.A2(n_52),
.B1(n_30),
.B2(n_34),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_176),
.A2(n_178),
.B1(n_185),
.B2(n_187),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_109),
.A2(n_44),
.B1(n_36),
.B2(n_40),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_69),
.Y(n_179)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_179),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_62),
.B(n_34),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_206),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_66),
.A2(n_36),
.B1(n_28),
.B2(n_37),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_81),
.A2(n_37),
.B1(n_40),
.B2(n_32),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_188),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_89),
.A2(n_37),
.B1(n_40),
.B2(n_32),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_189),
.A2(n_198),
.B1(n_218),
.B2(n_156),
.Y(n_288)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_64),
.A2(n_37),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_63),
.Y(n_201)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_113),
.B(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_79),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_127),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_210),
.A2(n_198),
.B(n_146),
.C(n_186),
.Y(n_294)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_77),
.Y(n_213)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_64),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_112),
.B(n_3),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_216),
.B(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_106),
.B(n_3),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_72),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_61),
.Y(n_219)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_154),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g344 ( 
.A(n_222),
.B(n_255),
.C(n_274),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_224),
.Y(n_316)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_226),
.Y(n_351)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_137),
.Y(n_229)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_5),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_230),
.B(n_242),
.Y(n_306)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_231),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_140),
.B(n_106),
.C(n_101),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_232),
.B(n_274),
.CI(n_252),
.CON(n_334),
.SN(n_334)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_234),
.Y(n_327)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_156),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_239),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_131),
.A2(n_76),
.B1(n_73),
.B2(n_101),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_240),
.A2(n_238),
.B(n_272),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_7),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_151),
.B(n_8),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_254),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_172),
.B(n_9),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_246),
.B(n_247),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_172),
.B(n_10),
.Y(n_247)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_249),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_L g356 ( 
.A1(n_252),
.A2(n_283),
.B(n_293),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_131),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_253),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_173),
.B(n_11),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_141),
.Y(n_255)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_141),
.B(n_13),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_284),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_147),
.B(n_13),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_262),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_13),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_261),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_147),
.B(n_14),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_193),
.B(n_15),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_263),
.B(n_271),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_264),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_185),
.A2(n_15),
.B1(n_17),
.B2(n_189),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_265),
.A2(n_204),
.B1(n_207),
.B2(n_203),
.Y(n_309)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_139),
.Y(n_269)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_165),
.B(n_17),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_270),
.B(n_296),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_160),
.B(n_17),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_164),
.B(n_169),
.C(n_167),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_170),
.B(n_153),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_278),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_276),
.A2(n_261),
.B1(n_293),
.B2(n_235),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_165),
.B(n_181),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_190),
.Y(n_279)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_150),
.Y(n_280)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_142),
.Y(n_281)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_282),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_136),
.B(n_166),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_138),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_130),
.B(n_200),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_285),
.B(n_287),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_145),
.A2(n_157),
.B1(n_149),
.B2(n_148),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_152),
.B1(n_204),
.B2(n_207),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_135),
.B(n_209),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_288),
.A2(n_295),
.B1(n_265),
.B2(n_273),
.Y(n_314)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_162),
.Y(n_289)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_182),
.B(n_133),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_291),
.B(n_298),
.Y(n_333)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_197),
.Y(n_292)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_150),
.B(n_168),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_294),
.A2(n_228),
.B(n_256),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_192),
.A2(n_195),
.B1(n_220),
.B2(n_221),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_161),
.B(n_194),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_183),
.B(n_199),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_183),
.B(n_199),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_264),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_203),
.B(n_152),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_300),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_304),
.A2(n_310),
.B1(n_335),
.B2(n_280),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_240),
.B(n_186),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_307),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_309),
.A2(n_314),
.B1(n_329),
.B2(n_337),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_284),
.A2(n_186),
.B1(n_223),
.B2(n_283),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_312),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_283),
.B1(n_298),
.B2(n_299),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_SL g331 ( 
.A(n_236),
.B(n_245),
.C(n_243),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_331),
.B(n_338),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_358),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_261),
.A2(n_254),
.B1(n_291),
.B2(n_259),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_293),
.B(n_232),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_290),
.B(n_277),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_348),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_231),
.A2(n_239),
.B(n_237),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_346),
.A2(n_355),
.B(n_234),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_249),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_297),
.A2(n_237),
.B1(n_227),
.B2(n_229),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_350),
.A2(n_357),
.B1(n_226),
.B2(n_234),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_225),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_225),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_228),
.A2(n_279),
.B1(n_257),
.B2(n_241),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_360),
.A2(n_367),
.B1(n_388),
.B2(n_323),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_330),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_368),
.Y(n_414)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_352),
.Y(n_365)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_329),
.A2(n_250),
.B1(n_266),
.B2(n_281),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_366),
.A2(n_369),
.B1(n_377),
.B2(n_380),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_337),
.A2(n_269),
.B1(n_250),
.B2(n_244),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_248),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_310),
.A2(n_266),
.B1(n_244),
.B2(n_248),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_317),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_371),
.B(n_374),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_372),
.A2(n_391),
.B(n_398),
.Y(n_404)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_258),
.C(n_268),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_375),
.B(n_376),
.C(n_379),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_303),
.B(n_341),
.C(n_313),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_355),
.A2(n_358),
.B1(n_309),
.B2(n_335),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_303),
.B(n_268),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_267),
.B1(n_277),
.B2(n_289),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_381),
.B(n_382),
.Y(n_413)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_395),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_386),
.Y(n_407)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_305),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_387),
.B(n_389),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_312),
.A2(n_267),
.B1(n_282),
.B2(n_292),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_301),
.B(n_233),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_390),
.A2(n_327),
.B1(n_324),
.B2(n_332),
.Y(n_417)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_392),
.B(n_394),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_307),
.A2(n_251),
.B1(n_304),
.B2(n_302),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_393),
.A2(n_322),
.B1(n_347),
.B2(n_345),
.Y(n_430)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

INVx8_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_396),
.Y(n_421)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_399),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_326),
.A2(n_316),
.B(n_349),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_339),
.A2(n_346),
.B(n_302),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_400),
.A2(n_327),
.B(n_315),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_306),
.B(n_321),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_401),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_334),
.B(n_353),
.C(n_326),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_325),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_340),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_324),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_359),
.B(n_334),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_405),
.B(n_406),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_306),
.C(n_308),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_409),
.A2(n_410),
.B1(n_417),
.B2(n_424),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_384),
.A2(n_354),
.B1(n_336),
.B2(n_308),
.Y(n_410)
);

OAI32xp33_ASAP7_75t_L g411 ( 
.A1(n_361),
.A2(n_342),
.A3(n_343),
.B1(n_328),
.B2(n_331),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_373),
.A2(n_332),
.B(n_342),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_416),
.B(n_420),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_400),
.A2(n_315),
.B(n_323),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_377),
.A2(n_319),
.B1(n_324),
.B2(n_322),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_403),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_368),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_428),
.B(n_376),
.Y(n_451)
);

XOR2x2_ASAP7_75t_SL g429 ( 
.A(n_379),
.B(n_328),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_438),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_430),
.A2(n_436),
.B1(n_365),
.B2(n_364),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_385),
.A2(n_318),
.B1(n_345),
.B2(n_351),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_431),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_391),
.A2(n_351),
.B(n_318),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_433),
.A2(n_440),
.B(n_372),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_360),
.A2(n_325),
.B1(n_347),
.B2(n_397),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_398),
.A2(n_373),
.B(n_402),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_435),
.Y(n_441)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_441),
.Y(n_481)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_435),
.Y(n_443)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_444),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_445),
.A2(n_450),
.B1(n_466),
.B2(n_473),
.Y(n_486)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_446),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_439),
.B(n_375),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_449),
.B(n_454),
.C(n_464),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_436),
.A2(n_388),
.B1(n_367),
.B2(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_452),
.A2(n_404),
.B(n_412),
.Y(n_493)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_423),
.Y(n_453)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_453),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_413),
.B(n_378),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_428),
.A2(n_393),
.B1(n_369),
.B2(n_380),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_456),
.A2(n_408),
.B1(n_424),
.B2(n_407),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_395),
.C(n_394),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_461),
.C(n_469),
.Y(n_491)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_381),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_460),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_415),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_392),
.C(n_387),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_396),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_462),
.Y(n_487)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_467),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_362),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_410),
.A2(n_371),
.B1(n_399),
.B2(n_363),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_437),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_383),
.C(n_370),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_470),
.Y(n_498)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_472),
.Y(n_500)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_408),
.A2(n_374),
.B1(n_409),
.B2(n_430),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_418),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_418),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_429),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_475),
.B(n_478),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_476),
.A2(n_488),
.B1(n_492),
.B2(n_473),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_438),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_455),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_479),
.B(n_482),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_444),
.Y(n_480)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_406),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_406),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_484),
.B(n_495),
.C(n_496),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_440),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_499),
.C(n_471),
.Y(n_514)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_459),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_448),
.A2(n_414),
.B1(n_433),
.B2(n_416),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_493),
.A2(n_462),
.B(n_468),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_411),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_446),
.B(n_404),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_441),
.B(n_420),
.C(n_412),
.Y(n_499)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_502),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_453),
.B(n_413),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_504),
.B(n_442),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_448),
.B(n_443),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_513),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_486),
.A2(n_465),
.B1(n_442),
.B2(n_452),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_508),
.A2(n_521),
.B1(n_487),
.B2(n_526),
.Y(n_534)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_500),
.Y(n_509)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_514),
.Y(n_535)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_477),
.Y(n_513)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_499),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_516),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_491),
.B(n_458),
.C(n_470),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_517),
.B(n_529),
.C(n_478),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_487),
.A2(n_462),
.B1(n_468),
.B2(n_460),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_519),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_482),
.B(n_456),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_524),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_503),
.A2(n_497),
.B1(n_476),
.B2(n_498),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_498),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_522),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_530),
.Y(n_543)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_494),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_525),
.B(n_528),
.Y(n_545)
);

XNOR2x2_ASAP7_75t_SL g540 ( 
.A(n_526),
.B(n_527),
.Y(n_540)
);

FAx1_ASAP7_75t_SL g527 ( 
.A(n_484),
.B(n_407),
.CI(n_467),
.CON(n_527),
.SN(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_501),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_421),
.C(n_472),
.Y(n_529)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_493),
.A2(n_445),
.B(n_463),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_533),
.B(n_518),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_534),
.A2(n_508),
.B1(n_521),
.B2(n_492),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_495),
.C(n_475),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_537),
.B(n_539),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_485),
.C(n_479),
.Y(n_539)
);

BUFx12_ASAP7_75t_L g542 ( 
.A(n_519),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_542),
.Y(n_561)
);

INVxp33_ASAP7_75t_SL g544 ( 
.A(n_509),
.Y(n_544)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_544),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_L g546 ( 
.A1(n_510),
.A2(n_505),
.B(n_483),
.C(n_504),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_527),
.Y(n_554)
);

BUFx12_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_549),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_547),
.B(n_511),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_551),
.B(n_556),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_514),
.C(n_515),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_552),
.B(n_558),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_518),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_535),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_563),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_547),
.B(n_512),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_507),
.Y(n_557)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_545),
.B(n_515),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_562),
.B(n_564),
.C(n_566),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_538),
.B(n_483),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_537),
.B(n_531),
.C(n_520),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_565),
.A2(n_534),
.B1(n_543),
.B2(n_550),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_535),
.B(n_531),
.C(n_496),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_565),
.Y(n_567)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_567),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_569),
.B(n_572),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_571),
.A2(n_577),
.B1(n_563),
.B2(n_557),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_560),
.A2(n_532),
.B1(n_548),
.B2(n_555),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_543),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_573),
.B(n_559),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_541),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_574),
.B(n_576),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_552),
.B(n_536),
.C(n_546),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_554),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_562),
.B(n_421),
.C(n_548),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_580),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_570),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_585),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_568),
.B(n_579),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_577),
.A2(n_549),
.B(n_540),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_586),
.B(n_588),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_580),
.B(n_553),
.Y(n_588)
);

OAI211xp5_ASAP7_75t_SL g590 ( 
.A1(n_570),
.A2(n_549),
.B(n_540),
.C(n_542),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_590),
.A2(n_578),
.B(n_542),
.C(n_564),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_593),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_587),
.B(n_575),
.C(n_573),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_576),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_595),
.B(n_596),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_589),
.B(n_567),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_597),
.A2(n_590),
.B(n_586),
.Y(n_598)
);

OAI21xp33_ASAP7_75t_SL g604 ( 
.A1(n_598),
.A2(n_599),
.B(n_591),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_592),
.A2(n_584),
.B(n_582),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_601),
.B(n_600),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_602),
.A2(n_603),
.B1(n_604),
.B2(n_569),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_601),
.B(n_594),
.Y(n_603)
);

MAJx2_ASAP7_75t_L g607 ( 
.A(n_605),
.B(n_606),
.C(n_434),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_603),
.Y(n_606)
);

AOI221xp5_ASAP7_75t_L g608 ( 
.A1(n_607),
.A2(n_422),
.B1(n_426),
.B2(n_425),
.C(n_419),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_422),
.Y(n_609)
);


endmodule