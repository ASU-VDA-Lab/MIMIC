module fake_jpeg_13580_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_49),
.B(n_50),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_54),
.Y(n_106)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_68),
.Y(n_74)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_70),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_71),
.Y(n_78)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_23),
.B1(n_26),
.B2(n_20),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_77),
.A2(n_103),
.B(n_108),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_92),
.B1(n_110),
.B2(n_113),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_23),
.B1(n_26),
.B2(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_33),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_105),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_25),
.B1(n_50),
.B2(n_47),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_100),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_40),
.A2(n_24),
.B(n_20),
.C(n_19),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_32),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_30),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_28),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_21),
.B1(n_27),
.B2(n_22),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_39),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_55),
.A2(n_23),
.B1(n_26),
.B2(n_19),
.Y(n_113)
);

BUFx2_ASAP7_75t_SL g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_24),
.C(n_19),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_131),
.C(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_98),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_77),
.A2(n_43),
.B1(n_24),
.B2(n_47),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_126),
.A2(n_140),
.B1(n_154),
.B2(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_129),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_27),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_39),
.C(n_44),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_22),
.B1(n_21),
.B2(n_15),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_151),
.B(n_128),
.Y(n_175)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_143),
.Y(n_172)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_75),
.B(n_28),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_21),
.B1(n_22),
.B2(n_15),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_141),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_15),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_4),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_79),
.A2(n_28),
.B1(n_45),
.B2(n_44),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_150),
.B1(n_102),
.B2(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_14),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_3),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_85),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_153),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_91),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_82),
.A2(n_104),
.B1(n_76),
.B2(n_88),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_0),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_76),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_83),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_88),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_180),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_150),
.B1(n_122),
.B2(n_118),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_174),
.B1(n_175),
.B2(n_179),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_102),
.C(n_89),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_169),
.B(n_176),
.C(n_13),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_170),
.A2(n_183),
.B1(n_190),
.B2(n_141),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_129),
.A2(n_93),
.B1(n_84),
.B2(n_89),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_89),
.C(n_80),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_188),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_123),
.A2(n_84),
.B1(n_80),
.B2(n_73),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_127),
.B(n_0),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_120),
.A2(n_73),
.B1(n_83),
.B2(n_2),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_184),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_120),
.A2(n_83),
.B1(n_1),
.B2(n_3),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_157),
.Y(n_218)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_117),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_124),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_125),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_4),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_161),
.Y(n_198)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_124),
.B1(n_148),
.B2(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_201),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_139),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_145),
.B1(n_147),
.B2(n_140),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_203),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_139),
.B1(n_136),
.B2(n_138),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_172),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_154),
.B1(n_144),
.B2(n_130),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_206),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_171),
.A2(n_188),
.B1(n_197),
.B2(n_165),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_210),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_156),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_222),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_160),
.B(n_196),
.C(n_166),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

INVx6_ASAP7_75t_SL g212 ( 
.A(n_182),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_156),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_213),
.B(n_221),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_152),
.B1(n_132),
.B2(n_133),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_230),
.B1(n_173),
.B2(n_164),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_162),
.B(n_146),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

AOI211xp5_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_153),
.B(n_125),
.C(n_119),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_236),
.B(n_163),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_180),
.B(n_185),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_232),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_179),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_177),
.B(n_9),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_163),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_169),
.B(n_10),
.Y(n_235)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_173),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_241),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_170),
.B(n_174),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_243),
.A2(n_246),
.B(n_251),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_160),
.B(n_176),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_205),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_226),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_255),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_220),
.A2(n_189),
.B(n_195),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_216),
.A2(n_184),
.B1(n_189),
.B2(n_181),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_260),
.B1(n_266),
.B2(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_219),
.B(n_158),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_158),
.B(n_161),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.Y(n_279)
);

OAI22x1_ASAP7_75t_SL g266 ( 
.A1(n_216),
.A2(n_182),
.B1(n_194),
.B2(n_158),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_199),
.A2(n_164),
.B1(n_194),
.B2(n_13),
.Y(n_268)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_263),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_280),
.Y(n_318)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_283),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_207),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_284),
.B(n_299),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_236),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_215),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_291),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_202),
.B1(n_200),
.B2(n_230),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_300),
.B1(n_252),
.B2(n_266),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_210),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_208),
.C(n_213),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_294),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_215),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_209),
.B1(n_232),
.B2(n_203),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_247),
.B1(n_258),
.B2(n_259),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_201),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_255),
.C(n_254),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_296),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_234),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_301),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_212),
.C(n_224),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_254),
.C(n_242),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_233),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_256),
.A2(n_204),
.B1(n_228),
.B2(n_198),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_323),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_271),
.B(n_242),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_303),
.A2(n_295),
.B(n_297),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_240),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_309),
.C(n_310),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_275),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_261),
.C(n_262),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_261),
.C(n_266),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_281),
.A2(n_259),
.B1(n_239),
.B2(n_247),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_316),
.B1(n_300),
.B2(n_299),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_314),
.A2(n_322),
.B1(n_280),
.B2(n_276),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_274),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_321),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_281),
.A2(n_258),
.B1(n_272),
.B2(n_245),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_320),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_252),
.B1(n_243),
.B2(n_268),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_245),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_293),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_328),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_330),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_303),
.A2(n_279),
.B(n_273),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_284),
.C(n_279),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_332),
.B(n_341),
.Y(n_361)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_335),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_315),
.B(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_314),
.A2(n_296),
.B1(n_291),
.B2(n_286),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_337),
.A2(n_344),
.B1(n_312),
.B2(n_321),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_342),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_339),
.A2(n_345),
.B1(n_346),
.B2(n_322),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_301),
.C(n_282),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_309),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_260),
.B1(n_267),
.B2(n_265),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_323),
.A2(n_204),
.B(n_270),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_347),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_363),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_333),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_358),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_331),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_359),
.Y(n_364)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_355),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_334),
.A2(n_310),
.B1(n_304),
.B2(n_312),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_340),
.Y(n_360)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_353),
.A2(n_340),
.B(n_346),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_369),
.B(n_355),
.Y(n_380)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_362),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_367),
.Y(n_378)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_336),
.C(n_330),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_342),
.C(n_331),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_370),
.Y(n_379)
);

AO221x1_ASAP7_75t_L g370 ( 
.A1(n_354),
.A2(n_338),
.B1(n_328),
.B2(n_335),
.C(n_329),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_332),
.C(n_339),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_372),
.B(n_375),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_307),
.C(n_344),
.Y(n_375)
);

OAI221xp5_ASAP7_75t_L g376 ( 
.A1(n_351),
.A2(n_313),
.B1(n_347),
.B2(n_308),
.C(n_337),
.Y(n_376)
);

NAND4xp25_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_308),
.C(n_319),
.D(n_270),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_374),
.A2(n_348),
.B1(n_357),
.B2(n_358),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

A2O1A1Ixp33_ASAP7_75t_SL g388 ( 
.A1(n_380),
.A2(n_384),
.B(n_375),
.C(n_373),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_356),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_381),
.A2(n_237),
.B(n_211),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_349),
.C(n_345),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_383),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_365),
.A2(n_313),
.B1(n_356),
.B2(n_319),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_371),
.A2(n_229),
.B1(n_237),
.B2(n_214),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_381),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_214),
.C(n_270),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_373),
.C(n_229),
.Y(n_391)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_378),
.A2(n_372),
.B(n_364),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_389),
.A2(n_383),
.B(n_385),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_390),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_386),
.Y(n_399)
);

AOI31xp67_ASAP7_75t_L g398 ( 
.A1(n_393),
.A2(n_394),
.A3(n_396),
.B(n_380),
.Y(n_398)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_379),
.A2(n_211),
.B(n_11),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_387),
.B(n_211),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_382),
.C(n_377),
.Y(n_397)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_397),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_398),
.B(n_388),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_402),
.B(n_392),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_403),
.Y(n_406)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_405),
.A2(n_400),
.B(n_401),
.Y(n_407)
);

AO21x1_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_404),
.B(n_11),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_406),
.C(n_12),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_12),
.Y(n_410)
);


endmodule