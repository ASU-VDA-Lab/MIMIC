module real_aes_2724_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_0), .B(n_115), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_1), .A2(n_124), .B(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_2), .A2(n_102), .B1(n_743), .B2(n_747), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_3), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_4), .B(n_115), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_5), .B(n_131), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_6), .B(n_131), .Y(n_501) );
INVx1_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_8), .B(n_131), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g775 ( .A(n_9), .Y(n_775) );
NAND2xp33_ASAP7_75t_L g482 ( .A(n_10), .B(n_133), .Y(n_482) );
AND2x2_ASAP7_75t_L g151 ( .A(n_11), .B(n_140), .Y(n_151) );
AND2x2_ASAP7_75t_L g160 ( .A(n_12), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g137 ( .A(n_13), .Y(n_137) );
AOI221x1_ASAP7_75t_L g523 ( .A1(n_14), .A2(n_25), .B1(n_115), .B2(n_124), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_15), .B(n_131), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_16), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_17), .B(n_115), .Y(n_478) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_18), .A2(n_140), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_19), .B(n_135), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_20), .B(n_131), .Y(n_461) );
AO21x1_ASAP7_75t_L g496 ( .A1(n_21), .A2(n_115), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_22), .B(n_115), .Y(n_185) );
INVx1_ASAP7_75t_L g448 ( .A(n_23), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_24), .A2(n_87), .B1(n_115), .B2(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_26), .Y(n_759) );
NAND2x1_ASAP7_75t_L g510 ( .A(n_27), .B(n_131), .Y(n_510) );
NAND2x1_ASAP7_75t_L g471 ( .A(n_28), .B(n_133), .Y(n_471) );
OR2x2_ASAP7_75t_L g138 ( .A(n_29), .B(n_84), .Y(n_138) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_29), .A2(n_84), .B(n_137), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_30), .B(n_133), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_31), .B(n_131), .Y(n_481) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_32), .A2(n_161), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_33), .B(n_133), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_34), .A2(n_124), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_35), .B(n_131), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_36), .A2(n_124), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g121 ( .A(n_37), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g125 ( .A(n_37), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g232 ( .A(n_37), .Y(n_232) );
OR2x6_ASAP7_75t_L g446 ( .A(n_38), .B(n_447), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g773 ( .A(n_38), .B(n_445), .C(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_39), .B(n_115), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_40), .B(n_115), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_41), .B(n_131), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_42), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_43), .B(n_133), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_44), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_45), .A2(n_124), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_46), .A2(n_124), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_47), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_48), .B(n_133), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_49), .B(n_115), .Y(n_167) );
INVx1_ASAP7_75t_L g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g128 ( .A(n_50), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_51), .A2(n_106), .B1(n_765), .B2(n_766), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_51), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_52), .B(n_131), .Y(n_158) );
AND2x2_ASAP7_75t_L g196 ( .A(n_53), .B(n_135), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_54), .B(n_133), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_55), .B(n_131), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_56), .B(n_133), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_57), .A2(n_124), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_58), .B(n_115), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_59), .B(n_115), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_60), .A2(n_124), .B(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g191 ( .A(n_61), .B(n_136), .Y(n_191) );
AO21x1_ASAP7_75t_L g498 ( .A1(n_62), .A2(n_124), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_63), .B(n_115), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_64), .B(n_133), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_65), .B(n_115), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_66), .B(n_133), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_67), .A2(n_93), .B1(n_124), .B2(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_68), .B(n_131), .Y(n_188) );
AND2x2_ASAP7_75t_L g546 ( .A(n_69), .B(n_136), .Y(n_546) );
INVx1_ASAP7_75t_L g120 ( .A(n_70), .Y(n_120) );
INVx1_ASAP7_75t_L g126 ( .A(n_70), .Y(n_126) );
AND2x2_ASAP7_75t_L g474 ( .A(n_71), .B(n_161), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_72), .B(n_133), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_73), .A2(n_124), .B(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_74), .A2(n_124), .B(n_129), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_75), .A2(n_124), .B(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g182 ( .A(n_76), .B(n_136), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_77), .B(n_135), .Y(n_221) );
INVx1_ASAP7_75t_L g449 ( .A(n_78), .Y(n_449) );
INVx1_ASAP7_75t_L g102 ( .A(n_79), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_80), .B(n_115), .Y(n_463) );
AND2x2_ASAP7_75t_L g484 ( .A(n_81), .B(n_161), .Y(n_484) );
AND2x2_ASAP7_75t_L g139 ( .A(n_82), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g497 ( .A(n_83), .B(n_172), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_85), .B(n_133), .Y(n_462) );
AND2x2_ASAP7_75t_L g513 ( .A(n_86), .B(n_161), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_88), .B(n_131), .Y(n_544) );
INVxp33_ASAP7_75t_L g777 ( .A(n_89), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_90), .A2(n_124), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_91), .B(n_133), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_92), .A2(n_124), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_94), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_95), .B(n_131), .Y(n_489) );
BUFx2_ASAP7_75t_L g190 ( .A(n_96), .Y(n_190) );
BUFx2_ASAP7_75t_L g753 ( .A(n_97), .Y(n_753) );
BUFx2_ASAP7_75t_SL g762 ( .A(n_97), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_98), .A2(n_124), .B(n_480), .Y(n_479) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_770), .B(n_776), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_750), .B(n_760), .Y(n_100) );
OAI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_103), .B(n_742), .Y(n_101) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_441), .B1(n_450), .B2(n_740), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_106), .A2(n_443), .B1(n_744), .B2(n_745), .Y(n_743) );
INVx5_ASAP7_75t_L g765 ( .A(n_106), .Y(n_765) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_345), .Y(n_106) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_270), .C(n_306), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_244), .Y(n_108) );
AOI211xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_162), .B(n_192), .C(n_217), .Y(n_109) );
AND2x2_ASAP7_75t_L g335 ( .A(n_110), .B(n_194), .Y(n_335) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_142), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_111), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g368 ( .A(n_111), .B(n_250), .Y(n_368) );
AND2x2_ASAP7_75t_L g384 ( .A(n_111), .B(n_209), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_111), .B(n_394), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_111), .B(n_418), .Y(n_417) );
INVx4_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_SL g204 ( .A(n_112), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g239 ( .A(n_112), .Y(n_239) );
AND2x2_ASAP7_75t_L g286 ( .A(n_112), .B(n_219), .Y(n_286) );
AND2x2_ASAP7_75t_L g305 ( .A(n_112), .B(n_142), .Y(n_305) );
BUFx2_ASAP7_75t_L g310 ( .A(n_112), .Y(n_310) );
AND2x2_ASAP7_75t_L g354 ( .A(n_112), .B(n_152), .Y(n_354) );
AND2x4_ASAP7_75t_L g426 ( .A(n_112), .B(n_427), .Y(n_426) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_112), .B(n_208), .Y(n_438) );
OR2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_139), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_123), .B(n_135), .Y(n_113) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_121), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
AND2x6_ASAP7_75t_L g133 ( .A(n_117), .B(n_126), .Y(n_133) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g131 ( .A(n_119), .B(n_128), .Y(n_131) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx5_ASAP7_75t_L g134 ( .A(n_121), .Y(n_134) );
AND2x2_ASAP7_75t_L g127 ( .A(n_122), .B(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_122), .Y(n_227) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx3_ASAP7_75t_L g228 ( .A(n_125), .Y(n_228) );
INVx2_ASAP7_75t_L g234 ( .A(n_126), .Y(n_234) );
AND2x4_ASAP7_75t_L g230 ( .A(n_127), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g226 ( .A(n_128), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_132), .B(n_134), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_133), .B(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_134), .A2(n_148), .B(n_149), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_134), .A2(n_157), .B(n_158), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_134), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_134), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_134), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_134), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_134), .A2(n_461), .B(n_462), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_134), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_134), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_134), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_134), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_134), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_134), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_134), .A2(n_543), .B(n_544), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_135), .Y(n_144) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_135), .A2(n_223), .B(n_229), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_135), .A2(n_486), .B(n_487), .Y(n_485) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_135), .A2(n_523), .B(n_527), .Y(n_522) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_135), .A2(n_523), .B(n_527), .Y(n_534) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x4_ASAP7_75t_L g172 ( .A(n_137), .B(n_138), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_140), .A2(n_185), .B(n_186), .Y(n_184) );
BUFx4f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_142), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g357 ( .A(n_142), .Y(n_357) );
BUFx2_ASAP7_75t_L g406 ( .A(n_142), .Y(n_406) );
INVx1_ASAP7_75t_L g428 ( .A(n_142), .Y(n_428) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_152), .Y(n_142) );
INVx3_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_143), .Y(n_394) );
AOI21x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_151), .Y(n_143) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_144), .A2(n_468), .B(n_474), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
INVx2_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_152), .B(n_205), .Y(n_209) );
INVx2_ASAP7_75t_L g294 ( .A(n_152), .Y(n_294) );
OR2x2_ASAP7_75t_L g301 ( .A(n_152), .B(n_250), .Y(n_301) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_160), .Y(n_152) );
INVx4_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_159), .Y(n_154) );
INVx3_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
AND2x2_ASAP7_75t_L g256 ( .A(n_162), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g290 ( .A(n_162), .B(n_253), .Y(n_290) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_173), .Y(n_162) );
AND2x2_ASAP7_75t_L g326 ( .A(n_163), .B(n_215), .Y(n_326) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g283 ( .A(n_164), .B(n_174), .Y(n_283) );
AND2x2_ASAP7_75t_L g402 ( .A(n_164), .B(n_183), .Y(n_402) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
INVx1_ASAP7_75t_L g242 ( .A(n_165), .Y(n_242) );
AND2x2_ASAP7_75t_L g298 ( .A(n_165), .B(n_174), .Y(n_298) );
AND2x2_ASAP7_75t_L g303 ( .A(n_165), .B(n_195), .Y(n_303) );
OR2x2_ASAP7_75t_L g366 ( .A(n_165), .B(n_183), .Y(n_366) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_165), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_172), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_172), .A2(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_SL g457 ( .A(n_172), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_172), .A2(n_478), .B(n_479), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_172), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g194 ( .A(n_173), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g243 ( .A(n_173), .Y(n_243) );
NOR2x1_ASAP7_75t_SL g173 ( .A(n_174), .B(n_183), .Y(n_173) );
AO21x1_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_182), .Y(n_174) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_175), .A2(n_176), .B(n_182), .Y(n_216) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_175), .A2(n_507), .B(n_513), .Y(n_506) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_175), .A2(n_540), .B(n_546), .Y(n_539) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_175), .A2(n_540), .B(n_546), .Y(n_575) );
AO21x2_ASAP7_75t_L g578 ( .A1(n_175), .A2(n_507), .B(n_513), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_181), .Y(n_176) );
AND2x2_ASAP7_75t_L g211 ( .A(n_183), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_SL g269 ( .A(n_183), .Y(n_269) );
NAND2x1_ASAP7_75t_L g279 ( .A(n_183), .B(n_195), .Y(n_279) );
OR2x2_ASAP7_75t_L g284 ( .A(n_183), .B(n_212), .Y(n_284) );
BUFx2_ASAP7_75t_L g340 ( .A(n_183), .Y(n_340) );
AND2x2_ASAP7_75t_L g376 ( .A(n_183), .B(n_255), .Y(n_376) );
AND2x2_ASAP7_75t_L g387 ( .A(n_183), .B(n_215), .Y(n_387) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_191), .Y(n_183) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_203), .B1(n_209), .B2(n_210), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_194), .A2(n_384), .B1(n_434), .B2(n_439), .Y(n_433) );
INVx4_ASAP7_75t_L g212 ( .A(n_195), .Y(n_212) );
INVx2_ASAP7_75t_L g253 ( .A(n_195), .Y(n_253) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_195), .Y(n_324) );
OR2x2_ASAP7_75t_L g339 ( .A(n_195), .B(n_215), .Y(n_339) );
OR2x2_ASAP7_75t_SL g365 ( .A(n_195), .B(n_366), .Y(n_365) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AND2x2_ASAP7_75t_SL g203 ( .A(n_204), .B(n_206), .Y(n_203) );
INVx2_ASAP7_75t_SL g246 ( .A(n_204), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_204), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g314 ( .A(n_204), .B(n_262), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_204), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_205), .Y(n_261) );
AND2x2_ASAP7_75t_L g317 ( .A(n_205), .B(n_294), .Y(n_317) );
INVx1_ASAP7_75t_L g427 ( .A(n_205), .Y(n_427) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_207), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_207), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g235 ( .A(n_208), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_209), .B(n_368), .Y(n_367) );
AOI321xp33_ASAP7_75t_L g389 ( .A1(n_210), .A2(n_291), .A3(n_359), .B1(n_390), .B2(n_391), .C(n_395), .Y(n_389) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_213), .Y(n_210) );
INVxp67_ASAP7_75t_SL g288 ( .A(n_211), .Y(n_288) );
AND2x2_ASAP7_75t_L g313 ( .A(n_211), .B(n_242), .Y(n_313) );
AND2x2_ASAP7_75t_L g388 ( .A(n_211), .B(n_298), .Y(n_388) );
INVx1_ASAP7_75t_L g257 ( .A(n_212), .Y(n_257) );
BUFx2_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g374 ( .A(n_212), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g312 ( .A(n_213), .Y(n_312) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
BUFx2_ASAP7_75t_L g319 ( .A(n_214), .Y(n_319) );
INVx2_ASAP7_75t_L g255 ( .A(n_215), .Y(n_255) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_215), .Y(n_278) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AOI21xp33_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_237), .B(n_240), .Y(n_217) );
NOR2xp67_ASAP7_75t_L g371 ( .A(n_218), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_235), .Y(n_219) );
INVx3_ASAP7_75t_L g262 ( .A(n_220), .Y(n_262) );
AND2x2_ASAP7_75t_L g293 ( .A(n_220), .B(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
AND2x4_ASAP7_75t_L g250 ( .A(n_221), .B(n_222), .Y(n_250) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_228), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2x1p5_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g333 ( .A(n_235), .Y(n_333) );
INVx1_ASAP7_75t_SL g418 ( .A(n_236), .Y(n_418) );
INVxp33_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_239), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g344 ( .A(n_239), .B(n_301), .Y(n_344) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
AND2x2_ASAP7_75t_L g348 ( .A(n_241), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_241), .B(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_242), .B(n_279), .Y(n_334) );
NOR4xp25_ASAP7_75t_L g429 ( .A(n_242), .B(n_273), .C(n_430), .D(n_431), .Y(n_429) );
OR2x2_ASAP7_75t_L g397 ( .A(n_243), .B(n_398), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_251), .B1(n_256), .B2(n_258), .C(n_263), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g272 ( .A(n_247), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g309 ( .A(n_248), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g329 ( .A(n_249), .Y(n_329) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
BUFx3_ASAP7_75t_L g352 ( .A(n_250), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_250), .B(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
OR2x2_ASAP7_75t_L g296 ( .A(n_253), .B(n_297), .Y(n_296) );
INVxp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_255), .B(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx2_ASAP7_75t_L g273 ( .A(n_260), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_260), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g265 ( .A(n_262), .Y(n_265) );
OAI321xp33_ASAP7_75t_L g377 ( .A1(n_262), .A2(n_370), .A3(n_378), .B1(n_383), .B2(n_385), .C(n_389), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
OR2x2_ASAP7_75t_L g332 ( .A(n_265), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g432 ( .A(n_268), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_269), .B(n_312), .Y(n_311) );
NAND2xp33_ASAP7_75t_SL g412 ( .A(n_269), .B(n_283), .Y(n_412) );
OAI211xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .B(n_285), .C(n_289), .Y(n_270) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_280), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g381 ( .A(n_278), .Y(n_381) );
INVx3_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
OR2x2_ASAP7_75t_L g423 ( .A(n_279), .B(n_297), .Y(n_423) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_281), .A2(n_365), .B1(n_367), .B2(n_369), .Y(n_364) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_SL g363 ( .A(n_284), .Y(n_363) );
OR2x2_ASAP7_75t_L g440 ( .A(n_284), .B(n_297), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_291), .B(n_295), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_293), .B(n_310), .Y(n_409) );
AND2x2_ASAP7_75t_L g415 ( .A(n_293), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_302), .B2(n_304), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_297), .A2(n_340), .B(n_342), .C(n_344), .Y(n_341) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_300), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_300), .B(n_392), .Y(n_414) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g386 ( .A(n_303), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_305), .A2(n_337), .B(n_340), .C(n_341), .Y(n_336) );
NAND3xp33_ASAP7_75t_SL g306 ( .A(n_307), .B(n_321), .C(n_336), .Y(n_306) );
AOI222xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_313), .B2(n_314), .C1(n_315), .C2(n_318), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g370 ( .A(n_310), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_310), .B(n_343), .Y(n_396) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g330 ( .A(n_317), .Y(n_330) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OR2x2_ASAP7_75t_L g435 ( .A(n_319), .B(n_352), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_320), .A2(n_411), .B1(n_413), .B2(n_415), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_327), .B1(n_331), .B2(n_334), .C(n_335), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI21xp5_ASAP7_75t_SL g395 ( .A1(n_328), .A2(n_396), .B(n_397), .Y(n_395) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g343 ( .A(n_329), .Y(n_343) );
AND2x2_ASAP7_75t_L g437 ( .A(n_329), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g421 ( .A(n_333), .Y(n_421) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g350 ( .A(n_339), .B(n_340), .Y(n_350) );
INVx1_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
NOR3xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_377), .C(n_399), .Y(n_345) );
OAI211xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_351), .B(n_353), .C(n_358), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_348), .A2(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_364), .C(n_371), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g382 ( .A(n_365), .Y(n_382) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_366), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_368), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g430 ( .A(n_368), .Y(n_430) );
AND2x2_ASAP7_75t_L g420 ( .A(n_370), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g390 ( .A(n_372), .Y(n_390) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g398 ( .A(n_374), .Y(n_398) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_386), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_429), .Y(n_419) );
OAI21xp33_ASAP7_75t_SL g434 ( .A1(n_391), .A2(n_435), .B(n_436), .Y(n_434) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g399 ( .A(n_400), .B(n_410), .C(n_419), .D(n_433), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B1(n_407), .B2(n_408), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx6p67_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
AND2x6_ASAP7_75t_SL g444 ( .A(n_445), .B(n_446), .Y(n_444) );
OR2x6_ASAP7_75t_SL g740 ( .A(n_445), .B(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g749 ( .A(n_445), .B(n_446), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_445), .B(n_741), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_446), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_448), .B(n_449), .Y(n_772) );
INVx2_ASAP7_75t_L g744 ( .A(n_450), .Y(n_744) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_638), .Y(n_450) );
NAND3xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_550), .C(n_605), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_491), .B1(n_514), .B2(n_518), .C(n_528), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_475), .Y(n_453) );
AND2x2_ASAP7_75t_SL g516 ( .A(n_454), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g549 ( .A(n_454), .Y(n_549) );
AND2x2_ASAP7_75t_L g594 ( .A(n_454), .B(n_531), .Y(n_594) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_466), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g582 ( .A(n_456), .Y(n_582) );
INVx1_ASAP7_75t_L g592 ( .A(n_456), .Y(n_592) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_464), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_457), .B(n_465), .Y(n_464) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_457), .A2(n_458), .B(n_464), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_463), .Y(n_458) );
OR2x2_ASAP7_75t_L g571 ( .A(n_466), .B(n_476), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_466), .B(n_517), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_466), .B(n_483), .Y(n_615) );
INVx2_ASAP7_75t_L g624 ( .A(n_466), .Y(n_624) );
AND2x2_ASAP7_75t_L g645 ( .A(n_466), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g729 ( .A(n_466), .B(n_548), .Y(n_729) );
INVx4_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g557 ( .A(n_467), .B(n_483), .Y(n_557) );
AND2x2_ASAP7_75t_L g690 ( .A(n_467), .B(n_517), .Y(n_690) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_467), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
AND2x4_ASAP7_75t_L g644 ( .A(n_475), .B(n_645), .Y(n_644) );
AOI321xp33_ASAP7_75t_L g658 ( .A1(n_475), .A2(n_587), .A3(n_588), .B1(n_620), .B2(n_659), .C(n_662), .Y(n_658) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
BUFx3_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
INVx2_ASAP7_75t_L g548 ( .A(n_476), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_476), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g581 ( .A(n_476), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g614 ( .A(n_476), .Y(n_614) );
INVx5_ASAP7_75t_L g517 ( .A(n_483), .Y(n_517) );
NOR2x1_ASAP7_75t_SL g566 ( .A(n_483), .B(n_556), .Y(n_566) );
BUFx2_ASAP7_75t_L g661 ( .A(n_483), .Y(n_661) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVxp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_504), .Y(n_492) );
NOR2xp33_ASAP7_75t_SL g559 ( .A(n_493), .B(n_560), .Y(n_559) );
NOR4xp25_ASAP7_75t_L g662 ( .A(n_493), .B(n_656), .C(n_660), .D(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g700 ( .A(n_493), .Y(n_700) );
AND2x2_ASAP7_75t_L g734 ( .A(n_493), .B(n_674), .Y(n_734) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g589 ( .A(n_495), .Y(n_589) );
OAI21x1_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_498), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g503 ( .A(n_497), .Y(n_503) );
AOI33xp33_ASAP7_75t_L g730 ( .A1(n_504), .A2(n_532), .A3(n_563), .B1(n_579), .B2(n_685), .B3(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g520 ( .A(n_505), .B(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g530 ( .A(n_505), .B(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g537 ( .A(n_506), .Y(n_537) );
INVxp67_ASAP7_75t_L g618 ( .A(n_506), .Y(n_618) );
AND2x2_ASAP7_75t_L g674 ( .A(n_506), .B(n_539), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_514), .A2(n_696), .B(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_L g683 ( .A(n_515), .B(n_557), .Y(n_683) );
AND3x2_ASAP7_75t_L g685 ( .A(n_515), .B(n_569), .C(n_624), .Y(n_685) );
INVx3_ASAP7_75t_SL g637 ( .A(n_516), .Y(n_637) );
INVx4_ASAP7_75t_L g531 ( .A(n_517), .Y(n_531) );
AND2x2_ASAP7_75t_L g569 ( .A(n_517), .B(n_556), .Y(n_569) );
INVxp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g563 ( .A(n_521), .Y(n_563) );
AND2x4_ASAP7_75t_L g588 ( .A(n_521), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g651 ( .A(n_521), .B(n_539), .Y(n_651) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g621 ( .A(n_522), .Y(n_621) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_522), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_R g528 ( .A1(n_529), .A2(n_532), .B(n_536), .C(n_547), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g580 ( .A(n_531), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_531), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_531), .B(n_548), .Y(n_709) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g691 ( .A(n_533), .B(n_681), .Y(n_691) );
AND2x2_ASAP7_75t_SL g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g538 ( .A(n_534), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g560 ( .A(n_534), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g576 ( .A(n_534), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g609 ( .A(n_534), .B(n_589), .Y(n_609) );
AND2x4_ASAP7_75t_L g574 ( .A(n_535), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g598 ( .A(n_535), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g636 ( .A(n_535), .B(n_561), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g564 ( .A(n_537), .B(n_561), .Y(n_564) );
AND2x2_ASAP7_75t_L g579 ( .A(n_537), .B(n_539), .Y(n_579) );
BUFx2_ASAP7_75t_L g635 ( .A(n_537), .Y(n_635) );
AND2x2_ASAP7_75t_L g649 ( .A(n_537), .B(n_560), .Y(n_649) );
INVx2_ASAP7_75t_L g561 ( .A(n_539), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_545), .Y(n_540) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_547), .A2(n_598), .B1(n_600), .B2(n_604), .Y(n_597) );
INVx2_ASAP7_75t_SL g628 ( .A(n_547), .Y(n_628) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x2_ASAP7_75t_L g603 ( .A(n_548), .B(n_556), .Y(n_603) );
INVx1_ASAP7_75t_L g710 ( .A(n_549), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_583), .C(n_597), .Y(n_550) );
OAI221xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_558), .B1(n_562), .B2(n_565), .C(n_567), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
INVxp67_ASAP7_75t_SL g739 ( .A(n_555), .Y(n_739) );
INVx1_ASAP7_75t_L g702 ( .A(n_557), .Y(n_702) );
AND2x2_ASAP7_75t_SL g712 ( .A(n_557), .B(n_581), .Y(n_712) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_561), .B(n_589), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OR2x2_ASAP7_75t_L g595 ( .A(n_563), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g673 ( .A(n_563), .Y(n_673) );
AND2x2_ASAP7_75t_L g608 ( .A(n_564), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g654 ( .A(n_566), .B(n_614), .Y(n_654) );
AND2x2_ASAP7_75t_L g731 ( .A(n_566), .B(n_729), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_572), .B1(n_579), .B2(n_580), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g590 ( .A(n_571), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx2_ASAP7_75t_L g596 ( .A(n_574), .Y(n_596) );
AND2x4_ASAP7_75t_L g620 ( .A(n_574), .B(n_621), .Y(n_620) );
OAI21xp33_ASAP7_75t_SL g650 ( .A1(n_574), .A2(n_651), .B(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g677 ( .A(n_574), .B(n_635), .Y(n_677) );
INVx2_ASAP7_75t_L g599 ( .A(n_575), .Y(n_599) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_575), .Y(n_632) );
INVx1_ASAP7_75t_SL g656 ( .A(n_576), .Y(n_656) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g587 ( .A(n_578), .Y(n_587) );
AND2x4_ASAP7_75t_SL g681 ( .A(n_578), .B(n_599), .Y(n_681) );
AND2x2_ASAP7_75t_L g678 ( .A(n_581), .B(n_624), .Y(n_678) );
AND2x2_ASAP7_75t_L g704 ( .A(n_581), .B(n_690), .Y(n_704) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_582), .Y(n_626) );
INVx1_ASAP7_75t_L g646 ( .A(n_582), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_590), .B1(n_593), .B2(n_595), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_588), .B(n_599), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_588), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g727 ( .A(n_588), .Y(n_727) );
INVx2_ASAP7_75t_SL g652 ( .A(n_590), .Y(n_652) );
AND2x2_ASAP7_75t_L g664 ( .A(n_592), .B(n_624), .Y(n_664) );
INVx2_ASAP7_75t_L g670 ( .A(n_592), .Y(n_670) );
INVxp33_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g629 ( .A(n_595), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_598), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g720 ( .A(n_598), .Y(n_720) );
INVx1_ASAP7_75t_L g648 ( .A(n_600), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_601), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g659 ( .A(n_603), .B(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_603), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_627), .C(n_630), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_610), .B1(n_612), .B2(n_616), .C(n_619), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g725 ( .A(n_610), .Y(n_725) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g694 ( .A(n_611), .B(n_660), .Y(n_694) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g625 ( .A(n_614), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g696 ( .A(n_616), .Y(n_696) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g693 ( .A(n_617), .Y(n_693) );
INVx1_ASAP7_75t_L g699 ( .A(n_618), .Y(n_699) );
OR2x2_ASAP7_75t_L g722 ( .A(n_618), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_SL g631 ( .A(n_621), .Y(n_631) );
AND2x2_ASAP7_75t_L g701 ( .A(n_621), .B(n_681), .Y(n_701) );
AND2x2_ASAP7_75t_SL g733 ( .A(n_621), .B(n_634), .Y(n_733) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g738 ( .A(n_624), .Y(n_738) );
INVx1_ASAP7_75t_L g688 ( .A(n_626), .Y(n_688) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B(n_633), .C(n_637), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_631), .B(n_681), .Y(n_705) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_634), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g642 ( .A(n_636), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g723 ( .A(n_636), .Y(n_723) );
NAND4xp75_ASAP7_75t_L g638 ( .A(n_639), .B(n_695), .C(n_711), .D(n_732), .Y(n_638) );
NOR3x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_657), .C(n_679), .Y(n_639) );
NAND4xp75_ASAP7_75t_L g640 ( .A(n_641), .B(n_647), .C(n_650), .D(n_653), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_642), .B(n_644), .Y(n_641) );
AND2x2_ASAP7_75t_L g692 ( .A(n_643), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g717 ( .A(n_644), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_SL g706 ( .A(n_649), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_665), .Y(n_657) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_661), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_671), .B(n_675), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g697 ( .A1(n_669), .A2(n_698), .A3(n_702), .B1(n_703), .B2(n_705), .C1(n_706), .C2(n_707), .Y(n_697) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_670), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_673), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_674), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .B(n_684), .C(n_686), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_691), .B1(n_692), .B2(n_694), .Y(n_686) );
NOR2xp33_ASAP7_75t_SL g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_701), .Y(n_698) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_704), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g714 ( .A(n_709), .B(n_715), .Y(n_714) );
O2A1O1Ixp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B(n_718), .C(n_721), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_714), .B(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI221xp5_ASAP7_75t_SL g721 ( .A1(n_722), .A2(n_724), .B1(n_726), .B2(n_728), .C(n_730), .Y(n_721) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
CKINVDCx11_ASAP7_75t_R g746 ( .A(n_740), .Y(n_746) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
INVxp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_755), .A2(n_764), .B(n_767), .Y(n_763) );
NOR2xp33_ASAP7_75t_SL g755 ( .A(n_756), .B(n_759), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
BUFx2_ASAP7_75t_L g769 ( .A(n_758), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx3_ASAP7_75t_SL g779 ( .A(n_771), .Y(n_779) );
AND2x2_ASAP7_75t_SL g771 ( .A(n_772), .B(n_773), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
endmodule