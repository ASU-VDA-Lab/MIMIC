module fake_ariane_1805_n_2422 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2422);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2422;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2370;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_2415;
wire n_436;
wire n_324;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_261;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_348;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_374;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2394;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_2395;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_108),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_160),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_151),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_87),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_178),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_26),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_32),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_158),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_114),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_10),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_111),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_118),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_200),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_218),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_42),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_185),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_153),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_33),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_106),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_133),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_72),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_99),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_124),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_12),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_76),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_64),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_83),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_0),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g271 ( 
.A(n_202),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_208),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_177),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_105),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_181),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_138),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_168),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_1),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_57),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_197),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_213),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_80),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_205),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_46),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_146),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_11),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_6),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_206),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_65),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_84),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_16),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_42),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_98),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_176),
.Y(n_297)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_14),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_117),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_25),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_230),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_110),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_7),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_86),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_144),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_40),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_173),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_118),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_20),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_80),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_103),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_115),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_110),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_53),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_180),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_224),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_3),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_150),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_32),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_93),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_68),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_123),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_5),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_201),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_190),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_53),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_45),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_121),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_203),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_102),
.Y(n_334)
);

BUFx4f_ASAP7_75t_SL g335 ( 
.A(n_122),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_221),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_219),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_220),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_165),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_131),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_14),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_60),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_196),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_235),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_54),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_105),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_152),
.Y(n_347)
);

BUFx5_ASAP7_75t_L g348 ( 
.A(n_4),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_130),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_79),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_34),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_170),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_189),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_164),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_103),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_47),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_0),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_145),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_233),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_64),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_161),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_36),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_4),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_84),
.Y(n_364)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_60),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_96),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_36),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_184),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_112),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_129),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_223),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_232),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_227),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_34),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_75),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_111),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_44),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_207),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_135),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_211),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_169),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_215),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_91),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_225),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_75),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_157),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_24),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_35),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_20),
.Y(n_389)
);

BUFx2_ASAP7_75t_SL g390 ( 
.A(n_40),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_83),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_25),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_12),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_71),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_187),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_143),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_191),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_7),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_167),
.Y(n_399)
);

BUFx8_ASAP7_75t_SL g400 ( 
.A(n_13),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_43),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_106),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_69),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_62),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_116),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_9),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_41),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_86),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_198),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_35),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_120),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_94),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_222),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_69),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_214),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_102),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_71),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_47),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_59),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_179),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_117),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_182),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_112),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_156),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_174),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_166),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_114),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_132),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_104),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_5),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_67),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_52),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_24),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_101),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_210),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_101),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_195),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_38),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_97),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_48),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_51),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_62),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_23),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_92),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_51),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_15),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_147),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_172),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_109),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_78),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_79),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_72),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_142),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_127),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_2),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_57),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_52),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_192),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_107),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_89),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_91),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_134),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_305),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_298),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_298),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_400),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_272),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_298),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_298),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_311),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_305),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_298),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_298),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_458),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_298),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_239),
.B(n_243),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_298),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_277),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_315),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_311),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_278),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_298),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_349),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_359),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_386),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_315),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_422),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_348),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_256),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_256),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_348),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_374),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_348),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_374),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_401),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_401),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_236),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_348),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_348),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_458),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_348),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_417),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_348),
.B(n_2),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_252),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_417),
.Y(n_505)
);

BUFx6f_ASAP7_75t_SL g506 ( 
.A(n_328),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_295),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_452),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_452),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_279),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_339),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_238),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_241),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_348),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_320),
.B(n_6),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_348),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_365),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_301),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_365),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_365),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_253),
.B(n_8),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_239),
.B(n_243),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_245),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_365),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_365),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_328),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_307),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_285),
.B(n_430),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_390),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_308),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_365),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_390),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_365),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_364),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_247),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_251),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_276),
.Y(n_537)
);

INVxp33_ASAP7_75t_SL g538 ( 
.A(n_259),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_383),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_260),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_388),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_246),
.B(n_8),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_365),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_365),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_433),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_263),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_246),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_265),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_R g549 ( 
.A(n_462),
.B(n_119),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_434),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_258),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_258),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_266),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_267),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_439),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_266),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_286),
.B(n_299),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_286),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_328),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_268),
.Y(n_560)
);

INVxp33_ASAP7_75t_L g561 ( 
.A(n_276),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_270),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_280),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_283),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_287),
.Y(n_565)
);

INVxp33_ASAP7_75t_L g566 ( 
.A(n_288),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_299),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_282),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_291),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_294),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_296),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_316),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_306),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_306),
.B(n_9),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_288),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_317),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_292),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_253),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_309),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_443),
.B(n_10),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_445),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_451),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_322),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_R g584 ( 
.A(n_237),
.B(n_125),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_249),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_323),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_329),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_330),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_478),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_483),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_464),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_R g592 ( 
.A(n_512),
.B(n_240),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_470),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_467),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_481),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_464),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_521),
.B(n_253),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_465),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_497),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_470),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_547),
.B(n_367),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_470),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_484),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_468),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_465),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_476),
.B(n_309),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_469),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_469),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_472),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_485),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_473),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_473),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_475),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_487),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_475),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_466),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_489),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_470),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_474),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_468),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_470),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_528),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_513),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_477),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_523),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_477),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_482),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_482),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_535),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_488),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_488),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_491),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_491),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_547),
.B(n_367),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_551),
.B(n_367),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_R g639 ( 
.A(n_540),
.B(n_242),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_548),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_529),
.B(n_318),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_493),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_507),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_522),
.B(n_557),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_493),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_551),
.B(n_318),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_498),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_536),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_480),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_490),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_554),
.Y(n_652)
);

INVxp33_ASAP7_75t_SL g653 ( 
.A(n_560),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_498),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_562),
.B(n_244),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_480),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_518),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_499),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_563),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_552),
.B(n_327),
.Y(n_660)
);

BUFx6f_ASAP7_75t_SL g661 ( 
.A(n_568),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_511),
.B(n_526),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_499),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_501),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_552),
.B(n_553),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_564),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_480),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_480),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_480),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_501),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_527),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_480),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_570),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_514),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_514),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_516),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_553),
.B(n_405),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_546),
.Y(n_678)
);

OA21x2_ASAP7_75t_L g679 ( 
.A1(n_503),
.A2(n_340),
.B(n_327),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_516),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_517),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_517),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_519),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_556),
.B(n_340),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_R g685 ( 
.A(n_571),
.B(n_248),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_492),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_665),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_681),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_644),
.B(n_526),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_681),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_622),
.B(n_474),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_665),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_665),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_679),
.A2(n_521),
.B1(n_542),
.B2(n_506),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_606),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_625),
.B(n_559),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_625),
.B(n_500),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_681),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_606),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_644),
.B(n_500),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_606),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_593),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_674),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_674),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_674),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_603),
.B(n_559),
.Y(n_706)
);

NAND3x1_ASAP7_75t_L g707 ( 
.A(n_641),
.B(n_574),
.C(n_580),
.Y(n_707)
);

AND2x6_ASAP7_75t_L g708 ( 
.A(n_597),
.B(n_331),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_597),
.B(n_578),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_603),
.B(n_561),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_SL g711 ( 
.A(n_626),
.B(n_576),
.C(n_572),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_641),
.B(n_511),
.Y(n_712)
);

INVx5_ASAP7_75t_L g713 ( 
.A(n_593),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_601),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_679),
.A2(n_506),
.B1(n_471),
.B2(n_479),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_597),
.B(n_568),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_622),
.B(n_601),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_674),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_680),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_680),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_597),
.B(n_568),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_649),
.B(n_538),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_R g723 ( 
.A(n_619),
.B(n_586),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_675),
.B(n_587),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_675),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_675),
.B(n_588),
.Y(n_726)
);

INVx8_ASAP7_75t_L g727 ( 
.A(n_661),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_681),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_675),
.Y(n_730)
);

OR2x2_ASAP7_75t_SL g731 ( 
.A(n_620),
.B(n_486),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_680),
.Y(n_732)
);

AND3x2_ASAP7_75t_L g733 ( 
.A(n_620),
.B(n_463),
.C(n_504),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_649),
.A2(n_495),
.B1(n_496),
.B2(n_494),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_633),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_633),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_678),
.B(n_506),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_662),
.B(n_528),
.Y(n_738)
);

INVx5_ASAP7_75t_L g739 ( 
.A(n_593),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_592),
.B(n_347),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_681),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_603),
.B(n_566),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_633),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_678),
.A2(n_505),
.B1(n_509),
.B2(n_502),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_682),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_681),
.Y(n_747)
);

AND2x6_ASAP7_75t_L g748 ( 
.A(n_597),
.B(n_331),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_637),
.B(n_556),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_633),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_681),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_682),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_637),
.B(n_558),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_637),
.B(n_515),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_682),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_682),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_599),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_599),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_599),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_589),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_599),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_599),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_638),
.B(n_331),
.Y(n_763)
);

AND2x2_ASAP7_75t_SL g764 ( 
.A(n_679),
.B(n_285),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_600),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_681),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_623),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_623),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_623),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_590),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_594),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_662),
.B(n_515),
.Y(n_772)
);

OAI21xp33_ASAP7_75t_L g773 ( 
.A1(n_608),
.A2(n_567),
.B(n_558),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_608),
.B(n_532),
.C(n_565),
.Y(n_774)
);

INVx4_ASAP7_75t_SL g775 ( 
.A(n_661),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_592),
.B(n_347),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_638),
.B(n_537),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_623),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_653),
.B(n_506),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_591),
.B(n_568),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_679),
.A2(n_510),
.B1(n_585),
.B2(n_573),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_623),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_638),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_591),
.B(n_567),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_596),
.B(n_573),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_677),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_632),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_677),
.B(n_579),
.Y(n_788)
);

INVx4_ASAP7_75t_SL g789 ( 
.A(n_661),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_677),
.B(n_575),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_633),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_596),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_653),
.B(n_569),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_598),
.Y(n_794)
);

OAI21xp33_ASAP7_75t_L g795 ( 
.A1(n_647),
.A2(n_579),
.B(n_405),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_640),
.B(n_583),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_634),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_651),
.B(n_577),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_598),
.B(n_519),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_647),
.B(n_405),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_652),
.B(n_520),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_607),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_659),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_607),
.B(n_520),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_651),
.B(n_250),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_609),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_686),
.B(n_666),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_673),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_L g809 ( 
.A(n_609),
.B(n_610),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_610),
.B(n_303),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_660),
.B(n_684),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_660),
.B(n_684),
.Y(n_812)
);

INVxp33_ASAP7_75t_L g813 ( 
.A(n_686),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_634),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_634),
.B(n_320),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_634),
.B(n_375),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_595),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_605),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_593),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_611),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_634),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_661),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_611),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_SL g824 ( 
.A(n_661),
.B(n_549),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_R g825 ( 
.A(n_613),
.B(n_584),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_639),
.B(n_292),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_612),
.B(n_375),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_612),
.B(n_353),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_614),
.B(n_524),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_614),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_615),
.B(n_524),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_615),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_617),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_616),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_616),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_639),
.B(n_353),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_SL g837 ( 
.A(n_600),
.B(n_328),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_618),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_618),
.B(n_525),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_627),
.Y(n_840)
);

BUFx4f_ASAP7_75t_L g841 ( 
.A(n_679),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_627),
.B(n_300),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_629),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_629),
.B(n_300),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_679),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_630),
.B(n_304),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_630),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_631),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_643),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_655),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_847),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_764),
.A2(n_580),
.B1(n_413),
.B2(n_343),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_689),
.A2(n_262),
.B1(n_361),
.B2(n_354),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_850),
.B(n_655),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_744),
.A2(n_635),
.B(n_631),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_722),
.B(n_530),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_812),
.B(n_811),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_798),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_812),
.B(n_685),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_764),
.A2(n_413),
.B1(n_343),
.B2(n_269),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_709),
.B(n_304),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_811),
.B(n_685),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_730),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_850),
.B(n_683),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_781),
.A2(n_413),
.B1(n_343),
.B2(n_290),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_847),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_811),
.B(n_635),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_841),
.A2(n_642),
.B(n_636),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_801),
.B(n_636),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_696),
.B(n_642),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_712),
.B(n_534),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_709),
.B(n_783),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_710),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_708),
.A2(n_361),
.B1(n_373),
.B2(n_354),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_696),
.B(n_645),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_SL g876 ( 
.A1(n_730),
.A2(n_831),
.B(n_802),
.C(n_806),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_749),
.B(n_645),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_798),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_809),
.A2(n_654),
.B(n_648),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_730),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_749),
.B(n_648),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_708),
.A2(n_379),
.B1(n_382),
.B2(n_373),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_848),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_708),
.A2(n_382),
.B1(n_409),
.B2(n_379),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_753),
.B(n_654),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_695),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_728),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_709),
.B(n_310),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_710),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_695),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_841),
.A2(n_663),
.B(n_664),
.C(n_658),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_SL g892 ( 
.A1(n_837),
.A2(n_541),
.B1(n_545),
.B2(n_539),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_743),
.B(n_310),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_708),
.A2(n_425),
.B1(n_435),
.B2(n_409),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_848),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_841),
.A2(n_663),
.B(n_658),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_753),
.B(n_664),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_779),
.B(n_670),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_694),
.A2(n_413),
.B1(n_343),
.B2(n_342),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_708),
.A2(n_435),
.B1(n_448),
.B2(n_425),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_788),
.B(n_670),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_826),
.B(n_737),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_715),
.A2(n_763),
.B1(n_708),
.B2(n_748),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_788),
.B(n_676),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_699),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_783),
.B(n_676),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_826),
.B(n_683),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_794),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_815),
.B(n_378),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_793),
.B(n_550),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_697),
.B(n_341),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_697),
.B(n_555),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_765),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_813),
.B(n_581),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_815),
.B(n_381),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_815),
.B(n_395),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_816),
.B(n_285),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_727),
.B(n_303),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_748),
.A2(n_448),
.B1(n_271),
.B2(n_424),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_763),
.A2(n_394),
.B1(n_407),
.B2(n_274),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_813),
.B(n_582),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_763),
.A2(n_441),
.B1(n_419),
.B2(n_430),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_748),
.A2(n_271),
.B1(n_424),
.B2(n_282),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_748),
.A2(n_763),
.B1(n_828),
.B2(n_706),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_823),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_699),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_701),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_816),
.B(n_430),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_816),
.B(n_442),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_701),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_763),
.A2(n_346),
.B1(n_440),
.B2(n_303),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_706),
.B(n_350),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_700),
.B(n_643),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_723),
.B(n_351),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_809),
.A2(n_604),
.B(n_602),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_754),
.B(n_442),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_703),
.Y(n_937)
);

NOR3x1_ASAP7_75t_L g938 ( 
.A(n_787),
.B(n_313),
.C(n_312),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_754),
.B(n_312),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_763),
.A2(n_346),
.B1(n_440),
.B2(n_303),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_825),
.B(n_355),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_796),
.B(n_356),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_717),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_777),
.B(n_357),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_827),
.B(n_313),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_754),
.B(n_314),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_748),
.A2(n_377),
.B1(n_389),
.B2(n_387),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_792),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_827),
.B(n_800),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_830),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_803),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_777),
.B(n_790),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_743),
.B(n_314),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_791),
.A2(n_531),
.B(n_525),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_792),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_808),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_827),
.B(n_324),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_800),
.B(n_324),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_748),
.A2(n_346),
.B1(n_440),
.B2(n_303),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_832),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_700),
.B(n_657),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_800),
.B(n_326),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_725),
.Y(n_963)
);

INVx8_ASAP7_75t_L g964 ( 
.A(n_727),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_773),
.B(n_326),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_772),
.B(n_727),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_842),
.B(n_334),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_842),
.B(n_334),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_687),
.B(n_345),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_703),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_834),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_717),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_842),
.B(n_345),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_844),
.B(n_846),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_844),
.B(n_360),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_727),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_688),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_828),
.A2(n_346),
.B1(n_440),
.B2(n_303),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_716),
.A2(n_721),
.B1(n_820),
.B2(n_780),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_844),
.B(n_360),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_828),
.A2(n_440),
.B1(n_346),
.B2(n_420),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_846),
.B(n_362),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_846),
.B(n_692),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_693),
.B(n_362),
.Y(n_984)
);

AND3x1_ASAP7_75t_L g985 ( 
.A(n_734),
.B(n_366),
.C(n_363),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_786),
.B(n_363),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_820),
.B(n_366),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_835),
.Y(n_988)
);

AND2x4_ASAP7_75t_SL g989 ( 
.A(n_833),
.B(n_657),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_777),
.B(n_369),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_725),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_838),
.Y(n_992)
);

NOR2x1p5_ASAP7_75t_L g993 ( 
.A(n_711),
.B(n_369),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_735),
.A2(n_403),
.B(n_404),
.C(n_406),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_828),
.A2(n_440),
.B1(n_346),
.B2(n_293),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_790),
.B(n_376),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_840),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_790),
.B(n_735),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_735),
.B(n_376),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_791),
.A2(n_533),
.B(n_531),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_688),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_736),
.B(n_385),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_745),
.B(n_392),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_718),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_736),
.B(n_750),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_SL g1006 ( 
.A(n_822),
.B(n_249),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_724),
.B(n_393),
.Y(n_1007)
);

NOR2x2_ASAP7_75t_L g1008 ( 
.A(n_772),
.B(n_671),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_736),
.B(n_385),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_724),
.B(n_398),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_750),
.B(n_843),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_750),
.B(n_391),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_767),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_718),
.Y(n_1014)
);

BUFx5_ASAP7_75t_L g1015 ( 
.A(n_828),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_726),
.B(n_402),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_726),
.B(n_738),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_784),
.B(n_391),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_760),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_704),
.Y(n_1020)
);

OAI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_772),
.A2(n_459),
.B1(n_444),
.B2(n_403),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_849),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_828),
.A2(n_249),
.B1(n_293),
.B2(n_420),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_785),
.B(n_404),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_845),
.A2(n_420),
.B1(n_293),
.B2(n_337),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_991),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_964),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_1019),
.B(n_760),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_859),
.B(n_738),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_SL g1030 ( 
.A(n_1019),
.B(n_770),
.C(n_771),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_857),
.B(n_770),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_989),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_872),
.B(n_772),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_L g1034 ( 
.A(n_910),
.B(n_807),
.C(n_771),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_943),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_872),
.B(n_775),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_872),
.B(n_775),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_908),
.Y(n_1038)
);

AND3x1_ASAP7_75t_SL g1039 ( 
.A(n_993),
.B(n_418),
.C(n_406),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_991),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_870),
.B(n_875),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_872),
.B(n_775),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_908),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_1015),
.B(n_688),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_869),
.B(n_740),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_1015),
.B(n_688),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_964),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_902),
.B(n_774),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_871),
.A2(n_740),
.B1(n_836),
.B2(n_776),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_925),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_SL g1051 ( 
.A(n_887),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_886),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_974),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_SL g1054 ( 
.A(n_966),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_L g1055 ( 
.A(n_862),
.B(n_807),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_989),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_873),
.B(n_776),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_913),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_SL g1059 ( 
.A(n_856),
.B(n_818),
.C(n_817),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_853),
.A2(n_818),
.B(n_817),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_1015),
.B(n_690),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_964),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1015),
.B(n_690),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_925),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_886),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_964),
.B(n_849),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_943),
.Y(n_1067)
);

AND2x6_ASAP7_75t_L g1068 ( 
.A(n_924),
.B(n_775),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_852),
.A2(n_899),
.B1(n_865),
.B2(n_860),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_950),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_890),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_873),
.B(n_836),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_890),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_887),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_951),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_858),
.B(n_805),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_951),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_889),
.B(n_805),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1022),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_889),
.B(n_714),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_956),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_983),
.B(n_762),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_R g1083 ( 
.A(n_956),
.B(n_671),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_867),
.B(n_762),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_SL g1085 ( 
.A(n_942),
.B(n_932),
.C(n_911),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_977),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_960),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_1022),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_914),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_921),
.Y(n_1090)
);

AND3x1_ASAP7_75t_L g1091 ( 
.A(n_853),
.B(n_691),
.C(n_421),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_952),
.B(n_731),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_878),
.B(n_767),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_948),
.A2(n_845),
.B1(n_814),
.B2(n_821),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_905),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_966),
.B(n_924),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_972),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_905),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_907),
.B(n_797),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_912),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_960),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_912),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1013),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_948),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_861),
.B(n_797),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_971),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_971),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1017),
.A2(n_824),
.B1(n_707),
.B2(n_767),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_933),
.B(n_757),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_861),
.B(n_833),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_861),
.B(n_888),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_961),
.B(n_758),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_888),
.B(n_814),
.Y(n_1113)
);

BUFx4f_ASAP7_75t_L g1114 ( 
.A(n_966),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_977),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_976),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_888),
.B(n_821),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_988),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1005),
.A2(n_804),
.B(n_799),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_998),
.B(n_767),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_948),
.Y(n_1121)
);

AND2x6_ASAP7_75t_SL g1122 ( 
.A(n_945),
.B(n_418),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_854),
.B(n_759),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_926),
.Y(n_1124)
);

AND2x6_ASAP7_75t_L g1125 ( 
.A(n_874),
.B(n_789),
.Y(n_1125)
);

NOR2x1_ASAP7_75t_L g1126 ( 
.A(n_941),
.B(n_729),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_949),
.B(n_761),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_966),
.B(n_789),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_977),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_868),
.A2(n_719),
.B(n_705),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_877),
.B(n_881),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_R g1132 ( 
.A(n_976),
.B(n_833),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_976),
.B(n_789),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1008),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1008),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_893),
.B(n_789),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_988),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_885),
.B(n_720),
.Y(n_1138)
);

AND2x6_ASAP7_75t_L g1139 ( 
.A(n_874),
.B(n_690),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_926),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_897),
.B(n_901),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_918),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_992),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_927),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_945),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_992),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_997),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_977),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_904),
.B(n_732),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_864),
.B(n_944),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_892),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_893),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_947),
.A2(n_824),
.B1(n_707),
.B2(n_795),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1015),
.B(n_955),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1015),
.B(n_690),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_997),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_896),
.A2(n_839),
.B(n_829),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_953),
.B(n_741),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_977),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_945),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_879),
.A2(n_752),
.B(n_746),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_851),
.Y(n_1162)
);

OR2x2_ASAP7_75t_SL g1163 ( 
.A(n_985),
.B(n_733),
.Y(n_1163)
);

INVx6_ASAP7_75t_L g1164 ( 
.A(n_1001),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_851),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_945),
.Y(n_1166)
);

INVx6_ASAP7_75t_L g1167 ( 
.A(n_1001),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1001),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_866),
.Y(n_1169)
);

NOR2x1p5_ASAP7_75t_L g1170 ( 
.A(n_990),
.B(n_822),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_953),
.B(n_755),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_955),
.B(n_909),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_927),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_866),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_883),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1013),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_955),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_1001),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_883),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1013),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_895),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_903),
.A2(n_782),
.B1(n_778),
.B2(n_769),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_895),
.Y(n_1183)
);

OR2x2_ASAP7_75t_SL g1184 ( 
.A(n_985),
.B(n_421),
.Y(n_1184)
);

AND2x6_ASAP7_75t_L g1185 ( 
.A(n_882),
.B(n_698),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1020),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_936),
.B(n_756),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_915),
.B(n_768),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_L g1189 ( 
.A(n_1001),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_916),
.B(n_729),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_930),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_996),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1020),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_930),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_937),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1011),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_906),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_863),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_937),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_919),
.A2(n_436),
.B(n_444),
.C(n_461),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_963),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_970),
.Y(n_1202)
);

OR2x2_ASAP7_75t_SL g1203 ( 
.A(n_957),
.B(n_436),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_929),
.B(n_729),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_SL g1205 ( 
.A(n_934),
.B(n_410),
.C(n_408),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_970),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_969),
.B(n_963),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_969),
.B(n_863),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1004),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_987),
.B(n_742),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_939),
.B(n_946),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_863),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_993),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_SL g1214 ( 
.A(n_947),
.B(n_414),
.C(n_412),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_880),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1004),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_969),
.Y(n_1217)
);

CKINVDCx16_ASAP7_75t_R g1218 ( 
.A(n_882),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_R g1219 ( 
.A(n_918),
.B(n_822),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1142),
.A2(n_923),
.B(n_894),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1041),
.A2(n_894),
.B1(n_900),
.B2(n_884),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1152),
.B(n_1021),
.Y(n_1222)
);

CKINVDCx11_ASAP7_75t_R g1223 ( 
.A(n_1032),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1161),
.A2(n_935),
.B(n_855),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1038),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1131),
.B(n_967),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1157),
.A2(n_1000),
.B(n_954),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1119),
.A2(n_1014),
.B(n_1002),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1141),
.A2(n_1006),
.B(n_898),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1138),
.A2(n_1006),
.B(n_876),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1218),
.B(n_1007),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1149),
.A2(n_1045),
.B(n_1094),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1043),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1027),
.Y(n_1234)
);

AOI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1044),
.A2(n_979),
.B(n_999),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1028),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1051),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1031),
.B(n_968),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1089),
.B(n_1010),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1089),
.B(n_1016),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1114),
.B(n_880),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1035),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1056),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1083),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1050),
.Y(n_1245)
);

BUFx2_ASAP7_75t_SL g1246 ( 
.A(n_1032),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1210),
.A2(n_891),
.B(n_880),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1127),
.A2(n_923),
.B(n_919),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1154),
.A2(n_1012),
.B(n_1009),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1154),
.A2(n_1014),
.B(n_742),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1044),
.A2(n_928),
.B(n_917),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1031),
.B(n_973),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1046),
.A2(n_742),
.B(n_975),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1064),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1029),
.A2(n_1049),
.B(n_1172),
.C(n_1048),
.Y(n_1255)
);

NAND2xp33_ASAP7_75t_L g1256 ( 
.A(n_1139),
.B(n_1015),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1029),
.B(n_1015),
.Y(n_1257)
);

O2A1O1Ixp5_ASAP7_75t_L g1258 ( 
.A1(n_1046),
.A2(n_1018),
.B(n_1024),
.C(n_984),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1067),
.B(n_1003),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1200),
.A2(n_994),
.A3(n_965),
.B(n_958),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1061),
.A2(n_986),
.B(n_962),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1061),
.A2(n_982),
.B(n_980),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1063),
.A2(n_1025),
.B(n_940),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1063),
.A2(n_1155),
.B(n_1158),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1195),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1197),
.B(n_920),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1076),
.B(n_922),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1070),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1195),
.Y(n_1269)
);

CKINVDCx8_ASAP7_75t_R g1270 ( 
.A(n_1122),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1192),
.B(n_1078),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1053),
.B(n_884),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1155),
.A2(n_931),
.B(n_959),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1200),
.A2(n_1182),
.A3(n_1172),
.B(n_1127),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1187),
.A2(n_1023),
.B(n_995),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1028),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1208),
.A2(n_1101),
.B1(n_1106),
.B2(n_1087),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1199),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1056),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1115),
.A2(n_981),
.B(n_978),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1052),
.A2(n_656),
.A3(n_650),
.B(n_621),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1048),
.B(n_900),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1115),
.A2(n_604),
.B(n_602),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1189),
.B(n_698),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1060),
.B(n_698),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1027),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1115),
.A2(n_604),
.B(n_602),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1189),
.A2(n_747),
.B(n_698),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1058),
.B(n_371),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1189),
.A2(n_751),
.B(n_747),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_L g1291 ( 
.A(n_1034),
.B(n_423),
.C(n_416),
.Y(n_1291)
);

NAND2x1_ASAP7_75t_L g1292 ( 
.A(n_1164),
.B(n_747),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1159),
.B(n_747),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1133),
.A2(n_766),
.B(n_751),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1052),
.A2(n_650),
.A3(n_656),
.B(n_621),
.Y(n_1295)
);

AO32x2_ASAP7_75t_L g1296 ( 
.A1(n_1178),
.A2(n_938),
.A3(n_810),
.B1(n_461),
.B2(n_459),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1148),
.A2(n_604),
.B(n_602),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1148),
.A2(n_667),
.B(n_621),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1080),
.B(n_938),
.Y(n_1299)
);

AOI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1190),
.A2(n_656),
.B(n_650),
.Y(n_1300)
);

AOI31xp67_ASAP7_75t_L g1301 ( 
.A1(n_1108),
.A2(n_1209),
.A3(n_1199),
.B(n_1071),
.Y(n_1301)
);

NAND2x1_ASAP7_75t_L g1302 ( 
.A(n_1164),
.B(n_751),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1090),
.A2(n_1092),
.B1(n_1097),
.B2(n_1091),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1204),
.A2(n_810),
.B(n_713),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1148),
.A2(n_667),
.B(n_621),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1128),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1080),
.B(n_751),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1100),
.B(n_427),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1116),
.A2(n_766),
.B(n_819),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1111),
.B(n_766),
.Y(n_1310)
);

BUFx2_ASAP7_75t_SL g1311 ( 
.A(n_1056),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1065),
.A2(n_667),
.A3(n_668),
.B(n_456),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1208),
.A2(n_766),
.B1(n_450),
.B2(n_455),
.Y(n_1313)
);

AOI211x1_ASAP7_75t_L g1314 ( 
.A1(n_1107),
.A2(n_455),
.B(n_456),
.C(n_450),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_1071),
.B(n_1065),
.Y(n_1315)
);

AO21x1_ASAP7_75t_L g1316 ( 
.A1(n_1120),
.A2(n_668),
.B(n_667),
.Y(n_1316)
);

AOI211x1_ASAP7_75t_L g1317 ( 
.A1(n_1118),
.A2(n_544),
.B(n_543),
.C(n_533),
.Y(n_1317)
);

NOR2x1_ASAP7_75t_SL g1318 ( 
.A(n_1047),
.B(n_819),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1073),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1096),
.B(n_819),
.Y(n_1320)
);

NAND3x1_ASAP7_75t_L g1321 ( 
.A(n_1055),
.B(n_431),
.C(n_429),
.Y(n_1321)
);

CKINVDCx9p33_ASAP7_75t_R g1322 ( 
.A(n_1074),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_SL g1323 ( 
.A1(n_1178),
.A2(n_668),
.B(n_544),
.Y(n_1323)
);

NOR2xp67_ASAP7_75t_L g1324 ( 
.A(n_1075),
.B(n_702),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1069),
.B(n_438),
.C(n_432),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_L g1326 ( 
.A(n_1160),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1211),
.B(n_446),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1073),
.A2(n_668),
.B(n_543),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1102),
.A2(n_449),
.B1(n_457),
.B2(n_460),
.C(n_337),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1095),
.A2(n_819),
.B(n_713),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1082),
.A2(n_1084),
.B(n_1099),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1027),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1095),
.A2(n_713),
.B(n_702),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1098),
.A2(n_713),
.B(n_702),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1137),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1116),
.A2(n_713),
.B(n_702),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1171),
.B(n_11),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1098),
.A2(n_739),
.B(n_702),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1162),
.A2(n_739),
.B(n_624),
.Y(n_1339)
);

NAND2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1114),
.B(n_739),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1027),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1083),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1171),
.B(n_15),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1093),
.B(n_16),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1159),
.B(n_1212),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1124),
.A2(n_739),
.B(n_337),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1124),
.A2(n_739),
.B(n_624),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1093),
.B(n_17),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1140),
.A2(n_672),
.A3(n_669),
.B(n_646),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1120),
.A2(n_255),
.B(n_254),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1140),
.A2(n_624),
.B(n_593),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1207),
.B(n_17),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1144),
.A2(n_672),
.B(n_669),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1159),
.B(n_311),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_L g1355 ( 
.A(n_1085),
.B(n_358),
.C(n_261),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1207),
.B(n_18),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1207),
.B(n_1143),
.Y(n_1357)
);

AND3x4_ASAP7_75t_L g1358 ( 
.A(n_1030),
.B(n_1059),
.C(n_1205),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1116),
.A2(n_368),
.B(n_264),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1116),
.A2(n_372),
.B(n_284),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1062),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1146),
.B(n_18),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_SL g1363 ( 
.A1(n_1178),
.A2(n_19),
.B(n_21),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1096),
.B(n_128),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1096),
.B(n_136),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1079),
.B(n_19),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1165),
.A2(n_672),
.B(n_669),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1144),
.A2(n_672),
.B(n_669),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1173),
.A2(n_672),
.B(n_669),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1088),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1173),
.Y(n_1371)
);

OA22x2_ASAP7_75t_L g1372 ( 
.A1(n_1217),
.A2(n_454),
.B1(n_453),
.B2(n_437),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1147),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1156),
.B(n_21),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1116),
.A2(n_302),
.B(n_257),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1196),
.A2(n_352),
.B(n_275),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_R g1377 ( 
.A(n_1047),
.B(n_273),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1110),
.B(n_1092),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1191),
.A2(n_672),
.B(n_669),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1191),
.A2(n_672),
.B(n_669),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1090),
.B(n_22),
.Y(n_1381)
);

INVx6_ASAP7_75t_L g1382 ( 
.A(n_1145),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1194),
.A2(n_672),
.B(n_669),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1153),
.A2(n_311),
.B(n_447),
.C(n_281),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1159),
.B(n_311),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1110),
.B(n_22),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1066),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1062),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1315),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1224),
.A2(n_1194),
.B(n_1174),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1224),
.A2(n_1175),
.B(n_1169),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1276),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1364),
.B(n_1365),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1364),
.B(n_1033),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1228),
.A2(n_1346),
.B(n_1351),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1282),
.A2(n_1151),
.B1(n_1135),
.B2(n_1134),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1228),
.A2(n_1181),
.B(n_1179),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1346),
.A2(n_1183),
.B(n_1202),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1306),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1364),
.B(n_1033),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1365),
.B(n_1033),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1365),
.B(n_1208),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1316),
.A2(n_1130),
.B(n_1186),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1306),
.B(n_1114),
.Y(n_1404)
);

NOR4xp25_ASAP7_75t_L g1405 ( 
.A(n_1255),
.B(n_1214),
.C(n_1193),
.D(n_1188),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1351),
.A2(n_1216),
.B(n_1206),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1221),
.A2(n_1185),
.B1(n_1139),
.B2(n_1166),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1353),
.A2(n_1215),
.B(n_1198),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1353),
.A2(n_1215),
.B(n_1198),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1384),
.A2(n_1130),
.B(n_1219),
.Y(n_1410)
);

CKINVDCx6p67_ASAP7_75t_R g1411 ( 
.A(n_1237),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1265),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1384),
.A2(n_1219),
.B(n_1123),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1230),
.A2(n_1072),
.B(n_1057),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1368),
.A2(n_1198),
.B(n_1215),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1368),
.A2(n_1126),
.B(n_1170),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1248),
.A2(n_1112),
.B(n_1109),
.Y(n_1417)
);

NAND2x1_ASAP7_75t_L g1418 ( 
.A(n_1294),
.B(n_1164),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1315),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1300),
.A2(n_1113),
.B(n_1105),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1306),
.B(n_1320),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1241),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1378),
.B(n_1320),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1255),
.A2(n_1117),
.B(n_1150),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1274),
.B(n_1203),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1229),
.A2(n_1150),
.B(n_1121),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1306),
.B(n_1159),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1265),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1269),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1238),
.A2(n_1081),
.B(n_1077),
.C(n_1104),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1236),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1235),
.A2(n_1136),
.B(n_1037),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1369),
.A2(n_1380),
.B(n_1379),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1369),
.A2(n_1380),
.B(n_1379),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1383),
.A2(n_1136),
.B(n_1068),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1320),
.B(n_1026),
.Y(n_1436)
);

AO32x2_ASAP7_75t_L g1437 ( 
.A1(n_1277),
.A2(n_1121),
.A3(n_1177),
.B1(n_1104),
.B2(n_1026),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1271),
.B(n_1145),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1232),
.A2(n_1037),
.B(n_1036),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1226),
.A2(n_1177),
.B(n_1139),
.Y(n_1440)
);

BUFx4_ASAP7_75t_SL g1441 ( 
.A(n_1236),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1241),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1252),
.B(n_1040),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1383),
.A2(n_1068),
.B(n_1086),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1269),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1303),
.B(n_1132),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1381),
.A2(n_1222),
.B1(n_1299),
.B2(n_1213),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1278),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1347),
.A2(n_1068),
.B(n_1086),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1347),
.A2(n_1068),
.B(n_1086),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1367),
.A2(n_1068),
.B(n_1086),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1381),
.A2(n_1213),
.B1(n_1184),
.B2(n_1039),
.C(n_1040),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1278),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1319),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1274),
.B(n_1103),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_R g1456 ( 
.A(n_1276),
.B(n_1160),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1319),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1242),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1333),
.A2(n_1338),
.B(n_1297),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1274),
.B(n_1103),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1333),
.A2(n_1068),
.B(n_1129),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1382),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1372),
.A2(n_1185),
.B1(n_1139),
.B2(n_1145),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1266),
.B(n_1166),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1258),
.A2(n_1139),
.B(n_1185),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1274),
.B(n_1176),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1371),
.Y(n_1467)
);

CKINVDCx16_ASAP7_75t_R g1468 ( 
.A(n_1237),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1312),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1338),
.A2(n_1129),
.B(n_1168),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1264),
.A2(n_1185),
.A3(n_1139),
.B(n_1125),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1283),
.A2(n_1298),
.B(n_1297),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1220),
.B(n_1128),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1283),
.A2(n_1129),
.B(n_1168),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_SL g1475 ( 
.A1(n_1247),
.A2(n_1132),
.B(n_1167),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1249),
.A2(n_1185),
.A3(n_1125),
.B(n_1054),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1312),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1231),
.B(n_1163),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1345),
.B(n_1128),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1281),
.Y(n_1480)
);

AND2x6_ASAP7_75t_L g1481 ( 
.A(n_1256),
.B(n_1036),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1298),
.A2(n_1129),
.B(n_1168),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1239),
.A2(n_1047),
.B1(n_1176),
.B2(n_1180),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1305),
.A2(n_1168),
.B(n_1167),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1312),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1267),
.A2(n_1185),
.B1(n_1125),
.B2(n_1066),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1340),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1312),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1382),
.B(n_1036),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1382),
.B(n_1037),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1370),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1305),
.A2(n_1167),
.B(n_1212),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1350),
.A2(n_1376),
.B(n_1348),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1334),
.A2(n_1212),
.B(n_1201),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1225),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1325),
.A2(n_1180),
.B(n_1042),
.C(n_1201),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1239),
.A2(n_1047),
.B1(n_1201),
.B2(n_1212),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1345),
.B(n_1201),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1308),
.B(n_1231),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1339),
.A2(n_1054),
.B(n_1047),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1372),
.A2(n_1125),
.B1(n_1042),
.B2(n_1133),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1272),
.A2(n_1125),
.B1(n_1042),
.B2(n_1133),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1342),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1330),
.A2(n_1125),
.B(n_1062),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1227),
.A2(n_384),
.B(n_321),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1256),
.B(n_1062),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1233),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1287),
.A2(n_646),
.B(n_624),
.Y(n_1508)
);

AOI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1257),
.A2(n_646),
.B(n_624),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1227),
.A2(n_646),
.B(n_624),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1251),
.A2(n_646),
.B(n_624),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1251),
.A2(n_646),
.B(n_624),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1344),
.A2(n_428),
.B(n_426),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1257),
.A2(n_646),
.B(n_593),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1261),
.A2(n_289),
.B(n_297),
.Y(n_1515)
);

INVx5_ASAP7_75t_L g1516 ( 
.A(n_1341),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1240),
.B(n_1259),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1328),
.A2(n_646),
.B(n_593),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1318),
.B(n_137),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1245),
.B(n_23),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1261),
.A2(n_593),
.B(n_447),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1240),
.B(n_335),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1250),
.A2(n_447),
.B(n_311),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1337),
.A2(n_370),
.B1(n_415),
.B2(n_411),
.Y(n_1524)
);

NAND4xp25_ASAP7_75t_L g1525 ( 
.A(n_1329),
.B(n_1291),
.C(n_1343),
.D(n_1314),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1262),
.A2(n_447),
.B(n_234),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1254),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1285),
.B(n_447),
.C(n_399),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1259),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1244),
.A2(n_447),
.B1(n_397),
.B2(n_396),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1268),
.B(n_26),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1234),
.B(n_139),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1253),
.A2(n_231),
.B(n_226),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1335),
.B(n_27),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1263),
.A2(n_380),
.B(n_344),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1286),
.B(n_140),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1309),
.A2(n_338),
.B(n_336),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1304),
.A2(n_212),
.B(n_204),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1332),
.B(n_141),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1354),
.A2(n_194),
.B(n_193),
.Y(n_1540)
);

AOI211xp5_ASAP7_75t_L g1541 ( 
.A1(n_1386),
.A2(n_333),
.B(n_332),
.C(n_325),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1281),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1285),
.A2(n_319),
.B(n_28),
.C(n_29),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1352),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1322),
.Y(n_1545)
);

OAI222xp33_ASAP7_75t_L g1546 ( 
.A1(n_1270),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C1(n_30),
.C2(n_31),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1373),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1354),
.A2(n_183),
.B(n_175),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1327),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1357),
.B(n_37),
.Y(n_1550)
);

NOR2xp67_ASAP7_75t_SL g1551 ( 
.A(n_1311),
.B(n_1388),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1331),
.A2(n_171),
.B(n_162),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1385),
.A2(n_159),
.B(n_155),
.Y(n_1553)
);

AO31x2_ASAP7_75t_L g1554 ( 
.A1(n_1301),
.A2(n_38),
.A3(n_39),
.B(n_41),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1281),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1263),
.A2(n_154),
.B(n_149),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1385),
.A2(n_1323),
.B(n_1336),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1289),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1332),
.B(n_148),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1307),
.A2(n_1310),
.B(n_1355),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1281),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1295),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1387),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1356),
.B(n_49),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1296),
.B(n_49),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1295),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_SL g1567 ( 
.A1(n_1284),
.A2(n_50),
.B(n_54),
.C(n_55),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1366),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1273),
.A2(n_56),
.B(n_58),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1295),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1246),
.B(n_58),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1545),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1411),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1493),
.A2(n_1321),
.B(n_1359),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1495),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1568),
.A2(n_1313),
.B1(n_1362),
.B2(n_1374),
.C(n_1363),
.Y(n_1576)
);

AND2x2_ASAP7_75t_SL g1577 ( 
.A(n_1407),
.B(n_1326),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1393),
.A2(n_1358),
.B1(n_1321),
.B2(n_1326),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1441),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1517),
.B(n_1296),
.Y(n_1580)
);

OAI222xp33_ASAP7_75t_L g1581 ( 
.A1(n_1393),
.A2(n_1296),
.B1(n_1284),
.B2(n_1279),
.C1(n_1243),
.C2(n_1293),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1495),
.Y(n_1582)
);

INVxp67_ASAP7_75t_SL g1583 ( 
.A(n_1455),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1522),
.A2(n_1360),
.B1(n_1375),
.B2(n_1324),
.C(n_1293),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1543),
.B(n_1317),
.C(n_1223),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1465),
.A2(n_1393),
.B(n_1440),
.Y(n_1586)
);

AO31x2_ASAP7_75t_L g1587 ( 
.A1(n_1480),
.A2(n_1290),
.A3(n_1288),
.B(n_1295),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1393),
.A2(n_1358),
.B1(n_1361),
.B2(n_1322),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1393),
.A2(n_1361),
.B1(n_1388),
.B2(n_1341),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1565),
.A2(n_1377),
.B1(n_1296),
.B2(n_1275),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1545),
.A2(n_1388),
.B1(n_1341),
.B2(n_1302),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1529),
.A2(n_1388),
.B1(n_1341),
.B2(n_1292),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1447),
.A2(n_1223),
.B1(n_1340),
.B2(n_1280),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1478),
.A2(n_1452),
.B1(n_1446),
.B2(n_1402),
.Y(n_1594)
);

OR2x6_ASAP7_75t_L g1595 ( 
.A(n_1473),
.B(n_1280),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1558),
.A2(n_1377),
.B1(n_61),
.B2(n_63),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_SL g1597 ( 
.A(n_1405),
.B(n_59),
.C(n_61),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1399),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1425),
.A2(n_1463),
.B1(n_1525),
.B2(n_1565),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1473),
.B(n_1275),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1423),
.B(n_63),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1475),
.A2(n_1260),
.B(n_1349),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1564),
.A2(n_1260),
.B1(n_66),
.B2(n_67),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_R g1604 ( 
.A(n_1499),
.B(n_65),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1425),
.A2(n_1260),
.B1(n_68),
.B2(n_70),
.Y(n_1605)
);

AOI222xp33_ASAP7_75t_L g1606 ( 
.A1(n_1546),
.A2(n_1260),
.B1(n_70),
.B2(n_73),
.C1(n_74),
.C2(n_76),
.Y(n_1606)
);

CKINVDCx11_ASAP7_75t_R g1607 ( 
.A(n_1431),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1507),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1525),
.A2(n_66),
.B1(n_73),
.B2(n_74),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1411),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1423),
.B(n_77),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1424),
.B(n_1349),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1417),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1520),
.B(n_81),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1541),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1396),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1443),
.B(n_88),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1527),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1475),
.A2(n_1450),
.B(n_1449),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1527),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1394),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1541),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1520),
.B(n_95),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1469),
.A2(n_1349),
.B(n_96),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1424),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1455),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1464),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1421),
.B(n_100),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1531),
.B(n_107),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1468),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1394),
.A2(n_108),
.B1(n_109),
.B2(n_113),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1469),
.A2(n_113),
.B(n_115),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1531),
.B(n_116),
.Y(n_1633)
);

NOR3xp33_ASAP7_75t_SL g1634 ( 
.A(n_1468),
.B(n_1549),
.C(n_1571),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1400),
.A2(n_1401),
.B1(n_1544),
.B2(n_1486),
.Y(n_1635)
);

INVx6_ASAP7_75t_L g1636 ( 
.A(n_1489),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1547),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1443),
.B(n_1458),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1405),
.A2(n_1513),
.B1(n_1430),
.B2(n_1438),
.C(n_1560),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1491),
.B(n_1550),
.Y(n_1640)
);

BUFx8_ASAP7_75t_L g1641 ( 
.A(n_1462),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1547),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1534),
.B(n_1550),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1392),
.Y(n_1644)
);

INVx4_ASAP7_75t_L g1645 ( 
.A(n_1516),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1524),
.A2(n_1502),
.B1(n_1402),
.B2(n_1501),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1473),
.A2(n_1490),
.B1(n_1489),
.B2(n_1563),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1427),
.Y(n_1648)
);

NAND2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1427),
.B(n_1399),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1400),
.A2(n_1401),
.B1(n_1534),
.B2(n_1481),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1503),
.B(n_1516),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1436),
.A2(n_1481),
.B1(n_1490),
.B2(n_1489),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1481),
.A2(n_1473),
.B1(n_1552),
.B2(n_1535),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1436),
.A2(n_1481),
.B1(n_1490),
.B2(n_1489),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_R g1655 ( 
.A(n_1481),
.B(n_1487),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1445),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_L g1657 ( 
.A(n_1551),
.B(n_1481),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1456),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1481),
.A2(n_1552),
.B1(n_1535),
.B2(n_1528),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1530),
.A2(n_1497),
.B1(n_1460),
.B2(n_1466),
.Y(n_1660)
);

BUFx2_ASAP7_75t_SL g1661 ( 
.A(n_1392),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1421),
.B(n_1490),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1460),
.A2(n_1466),
.B1(n_1552),
.B2(n_1490),
.Y(n_1663)
);

AOI222xp33_ASAP7_75t_L g1664 ( 
.A1(n_1456),
.A2(n_1528),
.B1(n_1426),
.B2(n_1457),
.C1(n_1428),
.C2(n_1412),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1535),
.A2(n_1488),
.B1(n_1485),
.B2(n_1477),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1427),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1412),
.B(n_1428),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1551),
.B(n_1429),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1453),
.B(n_1454),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1392),
.B(n_1479),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1453),
.B(n_1454),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1483),
.A2(n_1496),
.B1(n_1479),
.B2(n_1506),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1457),
.B(n_1467),
.Y(n_1673)
);

NAND2x1_ASAP7_75t_L g1674 ( 
.A(n_1498),
.B(n_1506),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1498),
.B(n_1422),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1399),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1498),
.B(n_1422),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1445),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1422),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1448),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1479),
.A2(n_1506),
.B1(n_1442),
.B2(n_1498),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1516),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1448),
.Y(n_1683)
);

NAND2xp33_ASAP7_75t_R g1684 ( 
.A(n_1556),
.B(n_1506),
.Y(n_1684)
);

INVx4_ASAP7_75t_SL g1685 ( 
.A(n_1476),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1516),
.B(n_1442),
.Y(n_1686)
);

AO31x2_ASAP7_75t_L g1687 ( 
.A1(n_1480),
.A2(n_1566),
.A3(n_1561),
.B(n_1542),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1516),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1390),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1532),
.B(n_1536),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1449),
.A2(n_1450),
.B(n_1451),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1532),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1451),
.A2(n_1439),
.B(n_1461),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1391),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1391),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1535),
.A2(n_1477),
.B1(n_1485),
.B2(n_1488),
.Y(n_1696)
);

NAND4xp25_ASAP7_75t_L g1697 ( 
.A(n_1567),
.B(n_1537),
.C(n_1532),
.D(n_1536),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1439),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1532),
.B(n_1536),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1397),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1404),
.Y(n_1701)
);

INVx4_ASAP7_75t_L g1702 ( 
.A(n_1539),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1413),
.A2(n_1410),
.B1(n_1569),
.B2(n_1505),
.Y(n_1703)
);

NAND2xp33_ASAP7_75t_SL g1704 ( 
.A(n_1418),
.B(n_1519),
.Y(n_1704)
);

NAND3x1_ASAP7_75t_L g1705 ( 
.A(n_1555),
.B(n_1570),
.C(n_1562),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1404),
.A2(n_1505),
.B1(n_1539),
.B2(n_1559),
.Y(n_1706)
);

CKINVDCx16_ASAP7_75t_R g1707 ( 
.A(n_1519),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1390),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1539),
.B(n_1559),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1395),
.A2(n_1521),
.B(n_1523),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1555),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1397),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1437),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1559),
.B(n_1476),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1559),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1519),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1570),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1538),
.A2(n_1540),
.B(n_1548),
.C(n_1553),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1439),
.B(n_1414),
.Y(n_1719)
);

NAND2x1p5_ASAP7_75t_L g1720 ( 
.A(n_1500),
.B(n_1519),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1414),
.B(n_1476),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1413),
.A2(n_1410),
.B1(n_1569),
.B2(n_1505),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1413),
.A2(n_1410),
.B1(n_1569),
.B2(n_1505),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1500),
.B(n_1435),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1403),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1437),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1403),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1476),
.Y(n_1729)
);

AOI21x1_ASAP7_75t_SL g1730 ( 
.A1(n_1515),
.A2(n_1554),
.B(n_1533),
.Y(n_1730)
);

AO22x1_ASAP7_75t_SL g1731 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1566),
.B2(n_1561),
.Y(n_1731)
);

OR2x6_ASAP7_75t_L g1732 ( 
.A(n_1435),
.B(n_1504),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1389),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1542),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1437),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1395),
.A2(n_1521),
.B(n_1523),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1437),
.Y(n_1737)
);

AO31x2_ASAP7_75t_L g1738 ( 
.A1(n_1419),
.A2(n_1515),
.A3(n_1554),
.B(n_1569),
.Y(n_1738)
);

BUFx4f_ASAP7_75t_SL g1739 ( 
.A(n_1471),
.Y(n_1739)
);

OR2x6_ASAP7_75t_L g1740 ( 
.A(n_1504),
.B(n_1461),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1444),
.B(n_1398),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1403),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1515),
.B(n_1414),
.C(n_1556),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1432),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1444),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1414),
.A2(n_1556),
.B1(n_1432),
.B2(n_1515),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1554),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1398),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1471),
.B(n_1554),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1556),
.A2(n_1514),
.B1(n_1509),
.B2(n_1434),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1432),
.A2(n_1538),
.B1(n_1420),
.B2(n_1548),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1471),
.B(n_1554),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1406),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1492),
.B(n_1484),
.Y(n_1754)
);

INVx6_ASAP7_75t_L g1755 ( 
.A(n_1492),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1406),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_SL g1757 ( 
.A(n_1526),
.B(n_1514),
.C(n_1509),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1470),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1420),
.B(n_1408),
.Y(n_1759)
);

AOI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1609),
.A2(n_1416),
.B1(n_1512),
.B2(n_1511),
.C(n_1494),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1607),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1594),
.B(n_1470),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1609),
.A2(n_1434),
.B1(n_1557),
.B2(n_1415),
.Y(n_1763)
);

OAI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1634),
.A2(n_1639),
.B1(n_1616),
.B2(n_1596),
.C(n_1606),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1613),
.A2(n_1434),
.B1(n_1557),
.B2(n_1415),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1643),
.B(n_1494),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1615),
.A2(n_1434),
.B1(n_1416),
.B2(n_1484),
.Y(n_1767)
);

OAI211xp5_ASAP7_75t_L g1768 ( 
.A1(n_1621),
.A2(n_1512),
.B(n_1511),
.C(n_1408),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1607),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1613),
.A2(n_1409),
.B1(n_1474),
.B2(n_1482),
.Y(n_1770)
);

OAI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1622),
.A2(n_1409),
.B1(n_1474),
.B2(n_1482),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1638),
.B(n_1580),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1575),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1640),
.B(n_1459),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1582),
.B(n_1510),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1680),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1605),
.A2(n_1518),
.B1(n_1510),
.B2(n_1433),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1605),
.A2(n_1518),
.B1(n_1472),
.B2(n_1508),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1572),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1625),
.A2(n_1472),
.B1(n_1508),
.B2(n_1597),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1608),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1625),
.A2(n_1597),
.B1(n_1616),
.B2(n_1599),
.Y(n_1782)
);

BUFx4f_ASAP7_75t_L g1783 ( 
.A(n_1577),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1699),
.A2(n_1702),
.B(n_1692),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1641),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1599),
.A2(n_1621),
.B1(n_1590),
.B2(n_1603),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1692),
.A2(n_1702),
.B(n_1709),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1627),
.A2(n_1631),
.B1(n_1574),
.B2(n_1634),
.C(n_1713),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1601),
.B(n_1611),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1631),
.A2(n_1627),
.B1(n_1585),
.B2(n_1576),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1614),
.A2(n_1623),
.B1(n_1629),
.B2(n_1633),
.C(n_1617),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1618),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1590),
.A2(n_1664),
.B1(n_1577),
.B2(n_1632),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1632),
.A2(n_1635),
.B1(n_1647),
.B2(n_1646),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1620),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_L g1796 ( 
.A1(n_1703),
.A2(n_1723),
.B(n_1722),
.C(n_1653),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1650),
.A2(n_1578),
.B1(n_1709),
.B2(n_1707),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1657),
.A2(n_1704),
.B(n_1706),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_R g1799 ( 
.A1(n_1588),
.A2(n_1628),
.B(n_1591),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1637),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1659),
.B(n_1722),
.C(n_1703),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1650),
.A2(n_1715),
.B1(n_1628),
.B2(n_1635),
.Y(n_1802)
);

BUFx4f_ASAP7_75t_L g1803 ( 
.A(n_1598),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_L g1804 ( 
.A(n_1659),
.B(n_1723),
.C(n_1653),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1647),
.A2(n_1663),
.B1(n_1660),
.B2(n_1697),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1663),
.A2(n_1698),
.B1(n_1714),
.B2(n_1593),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1743),
.B(n_1746),
.C(n_1668),
.Y(n_1807)
);

BUFx4f_ASAP7_75t_SL g1808 ( 
.A(n_1630),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_SL g1809 ( 
.A1(n_1739),
.A2(n_1714),
.B1(n_1655),
.B2(n_1715),
.Y(n_1809)
);

OAI211xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1610),
.A2(n_1747),
.B(n_1695),
.C(n_1694),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1644),
.A2(n_1573),
.B1(n_1658),
.B2(n_1652),
.Y(n_1811)
);

BUFx10_ASAP7_75t_L g1812 ( 
.A(n_1579),
.Y(n_1812)
);

AOI21xp33_ASAP7_75t_L g1813 ( 
.A1(n_1684),
.A2(n_1746),
.B(n_1752),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1573),
.Y(n_1814)
);

OAI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1654),
.A2(n_1586),
.B1(n_1716),
.B2(n_1672),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1726),
.A2(n_1735),
.B1(n_1737),
.B2(n_1581),
.C(n_1612),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1642),
.A2(n_1739),
.B1(n_1704),
.B2(n_1626),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1711),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1679),
.B(n_1690),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1626),
.B(n_1667),
.Y(n_1820)
);

AOI33xp33_ASAP7_75t_L g1821 ( 
.A1(n_1604),
.A2(n_1665),
.A3(n_1696),
.B1(n_1670),
.B2(n_1712),
.B3(n_1700),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1716),
.A2(n_1584),
.B1(n_1688),
.B2(n_1661),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1676),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1684),
.A2(n_1595),
.B1(n_1636),
.B2(n_1675),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1636),
.A2(n_1734),
.B1(n_1749),
.B2(n_1729),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1677),
.A2(n_1718),
.B1(n_1651),
.B2(n_1592),
.Y(n_1826)
);

OAI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1759),
.A2(n_1718),
.B(n_1719),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1598),
.B(n_1581),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1602),
.A2(n_1751),
.B(n_1589),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1669),
.Y(n_1830)
);

OAI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1595),
.A2(n_1674),
.B1(n_1662),
.B2(n_1681),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_L g1832 ( 
.A(n_1665),
.B(n_1696),
.C(n_1641),
.Y(n_1832)
);

AO221x2_ASAP7_75t_L g1833 ( 
.A1(n_1750),
.A2(n_1730),
.B1(n_1721),
.B2(n_1753),
.C(n_1756),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1598),
.B(n_1666),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1727),
.A2(n_1624),
.B1(n_1583),
.B2(n_1744),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1648),
.B(n_1666),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1727),
.A2(n_1624),
.B1(n_1583),
.B2(n_1744),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1649),
.A2(n_1720),
.B1(n_1645),
.B2(n_1682),
.Y(n_1838)
);

AOI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1711),
.A2(n_1717),
.B1(n_1742),
.B2(n_1728),
.C(n_1725),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1671),
.B(n_1673),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1655),
.Y(n_1841)
);

OAI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1600),
.A2(n_1701),
.B1(n_1682),
.B2(n_1645),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1731),
.B(n_1656),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1701),
.A2(n_1745),
.B1(n_1755),
.B2(n_1686),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1757),
.A2(n_1748),
.B1(n_1693),
.B2(n_1741),
.C(n_1755),
.Y(n_1845)
);

OAI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1757),
.A2(n_1741),
.B1(n_1755),
.B2(n_1724),
.C(n_1708),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1685),
.A2(n_1678),
.B1(n_1683),
.B2(n_1733),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1733),
.B(n_1754),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1724),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1689),
.A2(n_1758),
.B1(n_1754),
.B2(n_1619),
.C(n_1691),
.Y(n_1850)
);

OAI211xp5_ASAP7_75t_L g1851 ( 
.A1(n_1730),
.A2(n_1758),
.B(n_1710),
.C(n_1736),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1705),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1685),
.A2(n_1732),
.B1(n_1740),
.B2(n_1738),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1738),
.A2(n_1587),
.B1(n_1687),
.B2(n_1732),
.C(n_1740),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1738),
.A2(n_1609),
.B1(n_1393),
.B2(n_1517),
.Y(n_1855)
);

AOI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1609),
.A2(n_985),
.B1(n_910),
.B2(n_1625),
.C(n_689),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1575),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1598),
.Y(n_1858)
);

AOI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1603),
.A2(n_1505),
.B(n_1515),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1609),
.A2(n_1393),
.B1(n_1517),
.B2(n_1613),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1596),
.A2(n_910),
.B1(n_1089),
.B2(n_1090),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_SL g1862 ( 
.A1(n_1596),
.A2(n_1393),
.B1(n_1218),
.B2(n_837),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1575),
.Y(n_1863)
);

AOI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1603),
.A2(n_1505),
.B(n_1515),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1575),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1643),
.B(n_1638),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1572),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1609),
.B(n_1613),
.C(n_1639),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1643),
.B(n_1638),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1871)
);

OAI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1615),
.A2(n_1393),
.B1(n_1218),
.B2(n_1282),
.Y(n_1872)
);

OR2x6_ASAP7_75t_L g1873 ( 
.A(n_1595),
.B(n_1393),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1575),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1875)
);

OAI21xp33_ASAP7_75t_L g1876 ( 
.A1(n_1609),
.A2(n_1597),
.B(n_1613),
.Y(n_1876)
);

AO21x2_ASAP7_75t_L g1877 ( 
.A1(n_1743),
.A2(n_1757),
.B(n_1718),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1692),
.Y(n_1878)
);

OAI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1609),
.A2(n_1060),
.B1(n_910),
.B2(n_856),
.C(n_853),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1609),
.A2(n_1393),
.B1(n_1517),
.B2(n_1613),
.Y(n_1880)
);

AO31x2_ASAP7_75t_L g1881 ( 
.A1(n_1718),
.A2(n_1747),
.A3(n_1728),
.B(n_1742),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1609),
.A2(n_985),
.B1(n_910),
.B2(n_1625),
.C(n_689),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1609),
.A2(n_1393),
.B1(n_1517),
.B2(n_1613),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1638),
.B(n_1643),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1638),
.Y(n_1888)
);

BUFx4f_ASAP7_75t_L g1889 ( 
.A(n_1577),
.Y(n_1889)
);

OAI211xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1639),
.A2(n_1059),
.B(n_1034),
.C(n_793),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1643),
.B(n_1638),
.Y(n_1891)
);

AO21x2_ASAP7_75t_L g1892 ( 
.A1(n_1743),
.A2(n_1757),
.B(n_1718),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1643),
.B(n_1638),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1730),
.A2(n_1736),
.B(n_1710),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1643),
.B(n_1638),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1609),
.A2(n_689),
.B(n_1493),
.Y(n_1897)
);

OA21x2_ASAP7_75t_L g1898 ( 
.A1(n_1743),
.A2(n_1722),
.B(n_1703),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1572),
.Y(n_1899)
);

OAI21xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1609),
.A2(n_1546),
.B(n_1613),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1609),
.A2(n_1393),
.B1(n_1517),
.B2(n_1613),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1714),
.B(n_1715),
.Y(n_1902)
);

INVx4_ASAP7_75t_L g1903 ( 
.A(n_1692),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1641),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1643),
.B(n_1638),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1754),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1638),
.B(n_1643),
.Y(n_1907)
);

AOI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1603),
.A2(n_1505),
.B(n_1515),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1909)
);

OAI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1615),
.A2(n_1393),
.B1(n_1218),
.B2(n_1282),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1575),
.Y(n_1911)
);

AO21x2_ASAP7_75t_L g1912 ( 
.A1(n_1743),
.A2(n_1757),
.B(n_1718),
.Y(n_1912)
);

OAI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1609),
.A2(n_1060),
.B(n_910),
.C(n_1621),
.Y(n_1913)
);

AOI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1609),
.A2(n_985),
.B1(n_910),
.B2(n_1625),
.C(n_689),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1609),
.A2(n_1393),
.B1(n_1517),
.B2(n_1613),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1917)
);

NAND4xp25_ASAP7_75t_L g1918 ( 
.A(n_1609),
.B(n_722),
.C(n_793),
.D(n_1034),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1606),
.A2(n_1609),
.B1(n_1596),
.B2(n_1218),
.Y(n_1919)
);

BUFx4f_ASAP7_75t_SL g1920 ( 
.A(n_1630),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_SL g1921 ( 
.A1(n_1596),
.A2(n_1393),
.B1(n_1218),
.B2(n_837),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1906),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1906),
.B(n_1766),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1906),
.B(n_1833),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1867),
.B(n_1870),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1772),
.B(n_1820),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1891),
.B(n_1894),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1841),
.Y(n_1928)
);

INVxp33_ASAP7_75t_L g1929 ( 
.A(n_1789),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1818),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1795),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1896),
.B(n_1905),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1773),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1833),
.B(n_1827),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1781),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1808),
.B(n_1920),
.Y(n_1936)
);

NOR4xp25_ASAP7_75t_SL g1937 ( 
.A(n_1900),
.B(n_1764),
.C(n_1876),
.D(n_1788),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1792),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1833),
.B(n_1877),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1902),
.B(n_1873),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1800),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1774),
.B(n_1888),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1877),
.B(n_1892),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1840),
.B(n_1830),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1849),
.Y(n_1945)
);

OAI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1879),
.A2(n_1914),
.B1(n_1883),
.B2(n_1856),
.C(n_1866),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1892),
.B(n_1912),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1857),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1912),
.B(n_1898),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1898),
.B(n_1881),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1898),
.B(n_1881),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1882),
.B(n_1909),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1902),
.B(n_1863),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1761),
.B(n_1769),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1776),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1865),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1874),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1902),
.B(n_1911),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1823),
.Y(n_1959)
);

INVx1_ASAP7_75t_SL g1960 ( 
.A(n_1868),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1869),
.A2(n_1875),
.B1(n_1866),
.B2(n_1919),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1886),
.B(n_1907),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1881),
.B(n_1848),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1779),
.B(n_1899),
.Y(n_1964)
);

OR2x6_ASAP7_75t_L g1965 ( 
.A(n_1873),
.B(n_1798),
.Y(n_1965)
);

AND2x2_ASAP7_75t_SL g1966 ( 
.A(n_1783),
.B(n_1889),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1807),
.Y(n_1967)
);

OAI221xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1782),
.A2(n_1918),
.B1(n_1871),
.B2(n_1919),
.C(n_1887),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1816),
.B(n_1762),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_L g1970 ( 
.A1(n_1871),
.A2(n_1887),
.B1(n_1893),
.B2(n_1917),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1843),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1829),
.B(n_1850),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1775),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1852),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1895),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1845),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1762),
.B(n_1821),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1826),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1853),
.B(n_1765),
.Y(n_1979)
);

INVxp67_ASAP7_75t_L g1980 ( 
.A(n_1846),
.Y(n_1980)
);

INVx3_ASAP7_75t_SL g1981 ( 
.A(n_1814),
.Y(n_1981)
);

INVx4_ASAP7_75t_L g1982 ( 
.A(n_1783),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_L g1983 ( 
.A(n_1913),
.B(n_1890),
.C(n_1897),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1841),
.Y(n_1984)
);

AOI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1859),
.A2(n_1864),
.B(n_1908),
.Y(n_1985)
);

AO21x2_ASAP7_75t_L g1986 ( 
.A1(n_1801),
.A2(n_1804),
.B(n_1796),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1858),
.Y(n_1987)
);

INVxp67_ASAP7_75t_SL g1988 ( 
.A(n_1854),
.Y(n_1988)
);

BUFx3_ASAP7_75t_L g1989 ( 
.A(n_1889),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1763),
.B(n_1813),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1770),
.B(n_1777),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1836),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1810),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1821),
.B(n_1828),
.Y(n_1994)
);

INVxp67_ASAP7_75t_L g1995 ( 
.A(n_1828),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1851),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1805),
.B(n_1806),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1805),
.B(n_1806),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1803),
.B(n_1811),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1831),
.Y(n_2000)
);

AO21x2_ASAP7_75t_L g2001 ( 
.A1(n_1767),
.A2(n_1771),
.B(n_1768),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1777),
.B(n_1837),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1815),
.B(n_1855),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1835),
.B(n_1837),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1923),
.B(n_1835),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_R g2006 ( 
.A(n_1937),
.B(n_1769),
.Y(n_2006)
);

OAI211xp5_ASAP7_75t_SL g2007 ( 
.A1(n_1983),
.A2(n_1960),
.B(n_1946),
.C(n_1961),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1928),
.Y(n_2008)
);

OAI211xp5_ASAP7_75t_L g2009 ( 
.A1(n_1934),
.A2(n_1861),
.B(n_1782),
.C(n_1786),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1986),
.A2(n_1786),
.B1(n_1793),
.B2(n_1875),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1942),
.B(n_1832),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1931),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1955),
.Y(n_2013)
);

NAND2xp33_ASAP7_75t_SL g2014 ( 
.A(n_1981),
.B(n_1878),
.Y(n_2014)
);

O2A1O1Ixp33_ASAP7_75t_L g2015 ( 
.A1(n_1946),
.A2(n_1968),
.B(n_1983),
.C(n_1967),
.Y(n_2015)
);

OR2x6_ASAP7_75t_L g2016 ( 
.A(n_1965),
.B(n_1802),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1931),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1933),
.Y(n_2018)
);

OR2x6_ASAP7_75t_L g2019 ( 
.A(n_1965),
.B(n_1797),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1933),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1942),
.B(n_1794),
.Y(n_2021)
);

AOI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_1968),
.A2(n_1790),
.B1(n_1893),
.B2(n_1885),
.C(n_1917),
.Y(n_2022)
);

OAI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1969),
.A2(n_1884),
.B1(n_1916),
.B2(n_1901),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1923),
.B(n_1817),
.Y(n_2024)
);

AOI221xp5_ASAP7_75t_L g2025 ( 
.A1(n_1969),
.A2(n_1915),
.B1(n_1885),
.B2(n_1880),
.C(n_1860),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1935),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_R g2027 ( 
.A(n_1936),
.B(n_1814),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1923),
.B(n_1844),
.Y(n_2028)
);

INVx1_ASAP7_75t_SL g2029 ( 
.A(n_1981),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1924),
.B(n_1819),
.Y(n_2030)
);

OAI31xp33_ASAP7_75t_L g2031 ( 
.A1(n_1967),
.A2(n_1793),
.A3(n_1915),
.B(n_1910),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1924),
.B(n_1834),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1924),
.B(n_1794),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1992),
.B(n_1784),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_1977),
.A2(n_1872),
.B1(n_1791),
.B2(n_1862),
.C(n_1921),
.Y(n_2035)
);

INVx4_ASAP7_75t_L g2036 ( 
.A(n_1981),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1986),
.A2(n_1824),
.B1(n_1825),
.B2(n_1847),
.Y(n_2037)
);

BUFx6f_ASAP7_75t_L g2038 ( 
.A(n_1966),
.Y(n_2038)
);

NAND3xp33_ASAP7_75t_L g2039 ( 
.A(n_1943),
.B(n_1780),
.C(n_1839),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_1986),
.A2(n_1847),
.B1(n_1780),
.B2(n_1809),
.Y(n_2040)
);

OAI33xp33_ASAP7_75t_L g2041 ( 
.A1(n_1994),
.A2(n_1822),
.A3(n_1842),
.B1(n_1838),
.B2(n_1799),
.B3(n_1812),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1940),
.B(n_1904),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1960),
.B(n_1812),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1935),
.Y(n_2044)
);

OAI31xp33_ASAP7_75t_L g2045 ( 
.A1(n_1970),
.A2(n_1904),
.A3(n_1778),
.B(n_1785),
.Y(n_2045)
);

OAI31xp33_ASAP7_75t_L g2046 ( 
.A1(n_1997),
.A2(n_1998),
.A3(n_1977),
.B(n_1972),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1964),
.Y(n_2047)
);

OAI211xp5_ASAP7_75t_SL g2048 ( 
.A1(n_1930),
.A2(n_1760),
.B(n_1787),
.C(n_1778),
.Y(n_2048)
);

AOI33xp33_ASAP7_75t_L g2049 ( 
.A1(n_1937),
.A2(n_1812),
.A3(n_1878),
.B1(n_1903),
.B2(n_1934),
.B3(n_1939),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1938),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1941),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1941),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_SL g2053 ( 
.A1(n_1986),
.A2(n_1878),
.B1(n_1903),
.B2(n_1997),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1954),
.B(n_1903),
.Y(n_2054)
);

AOI211xp5_ASAP7_75t_L g2055 ( 
.A1(n_1934),
.A2(n_1939),
.B(n_1947),
.C(n_1943),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1930),
.Y(n_2056)
);

AOI221xp5_ASAP7_75t_L g2057 ( 
.A1(n_1994),
.A2(n_1988),
.B1(n_1990),
.B2(n_1993),
.C(n_1949),
.Y(n_2057)
);

AOI211xp5_ASAP7_75t_L g2058 ( 
.A1(n_1939),
.A2(n_1943),
.B(n_1947),
.C(n_1990),
.Y(n_2058)
);

AO21x2_ASAP7_75t_L g2059 ( 
.A1(n_1985),
.A2(n_1949),
.B(n_1947),
.Y(n_2059)
);

OAI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_2003),
.A2(n_1998),
.B1(n_1976),
.B2(n_1972),
.Y(n_2060)
);

INVx4_ASAP7_75t_L g2061 ( 
.A(n_1982),
.Y(n_2061)
);

OAI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_1972),
.A2(n_2003),
.B(n_1993),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1973),
.Y(n_2063)
);

INVx2_ASAP7_75t_SL g2064 ( 
.A(n_1953),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1953),
.B(n_1958),
.Y(n_2065)
);

NAND2xp33_ASAP7_75t_SL g2066 ( 
.A(n_1996),
.B(n_1945),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_SL g2067 ( 
.A1(n_1966),
.A2(n_1978),
.B1(n_1929),
.B2(n_1928),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1978),
.A2(n_1999),
.B1(n_1990),
.B2(n_1966),
.Y(n_2068)
);

NAND3xp33_ASAP7_75t_L g2069 ( 
.A(n_1949),
.B(n_1976),
.C(n_1988),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1948),
.Y(n_2070)
);

NAND3xp33_ASAP7_75t_L g2071 ( 
.A(n_1996),
.B(n_1974),
.C(n_1980),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1958),
.B(n_1979),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1979),
.B(n_1925),
.Y(n_2073)
);

OAI211xp5_ASAP7_75t_SL g2074 ( 
.A1(n_1974),
.A2(n_1959),
.B(n_1992),
.C(n_1980),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1959),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1948),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_1952),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1979),
.B(n_1925),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1927),
.B(n_1932),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1922),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1927),
.B(n_1932),
.Y(n_2081)
);

NOR2x1_ASAP7_75t_SL g2082 ( 
.A(n_1965),
.B(n_1989),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1940),
.B(n_1965),
.Y(n_2083)
);

NOR2x1_ASAP7_75t_L g2084 ( 
.A(n_1928),
.B(n_1984),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2073),
.B(n_1991),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2063),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2018),
.Y(n_2087)
);

NAND2x1p5_ASAP7_75t_L g2088 ( 
.A(n_2038),
.B(n_1982),
.Y(n_2088)
);

NOR2x1_ASAP7_75t_L g2089 ( 
.A(n_2084),
.B(n_1984),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2073),
.B(n_1926),
.Y(n_2090)
);

INVx2_ASAP7_75t_SL g2091 ( 
.A(n_2080),
.Y(n_2091)
);

NOR4xp25_ASAP7_75t_SL g2092 ( 
.A(n_2066),
.B(n_1945),
.C(n_2000),
.D(n_1987),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2078),
.B(n_2012),
.Y(n_2093)
);

NOR3xp33_ASAP7_75t_L g2094 ( 
.A(n_2015),
.B(n_1985),
.C(n_1991),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2059),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2078),
.B(n_1926),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2072),
.B(n_1991),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2017),
.B(n_1963),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2020),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2072),
.B(n_2079),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2059),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2026),
.Y(n_2102)
);

AND2x4_ASAP7_75t_SL g2103 ( 
.A(n_2038),
.B(n_1982),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2044),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2079),
.B(n_2001),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2059),
.B(n_1973),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2077),
.B(n_1962),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2058),
.B(n_1963),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2013),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2057),
.B(n_1963),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2056),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2081),
.B(n_2001),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2050),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2081),
.B(n_2001),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2065),
.B(n_2001),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2065),
.B(n_2002),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2005),
.B(n_2002),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2005),
.B(n_2002),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2034),
.B(n_1956),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2055),
.B(n_1956),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2047),
.B(n_1962),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_2080),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2024),
.B(n_1951),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2024),
.B(n_2028),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2051),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2052),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2070),
.B(n_1957),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2076),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2028),
.B(n_1951),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2064),
.B(n_2032),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2064),
.B(n_1951),
.Y(n_2131)
);

NOR2x1_ASAP7_75t_SL g2132 ( 
.A(n_2038),
.B(n_1965),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2032),
.B(n_1950),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2033),
.B(n_1957),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2030),
.B(n_1950),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2030),
.B(n_1950),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2082),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_2066),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2033),
.B(n_1922),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2021),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_2071),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2047),
.B(n_1952),
.Y(n_2142)
);

NAND2xp33_ASAP7_75t_R g2143 ( 
.A(n_2027),
.B(n_2004),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2087),
.Y(n_2144)
);

AND2x4_ASAP7_75t_SL g2145 ( 
.A(n_2139),
.B(n_2042),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_2090),
.B(n_2096),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2087),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2094),
.B(n_2062),
.Y(n_2148)
);

NAND2x1_ASAP7_75t_L g2149 ( 
.A(n_2138),
.B(n_2089),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2131),
.Y(n_2150)
);

AOI21xp5_ASAP7_75t_L g2151 ( 
.A1(n_2110),
.A2(n_2039),
.B(n_2069),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2113),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2113),
.Y(n_2153)
);

BUFx3_ASAP7_75t_L g2154 ( 
.A(n_2111),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_2142),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2094),
.B(n_2060),
.Y(n_2156)
);

INVx2_ASAP7_75t_SL g2157 ( 
.A(n_2142),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_2090),
.B(n_2021),
.Y(n_2158)
);

OAI32xp33_ASAP7_75t_L g2159 ( 
.A1(n_2110),
.A2(n_2141),
.A3(n_2108),
.B1(n_2143),
.B2(n_2007),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2085),
.B(n_2008),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2125),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2125),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2126),
.Y(n_2163)
);

NAND2xp33_ASAP7_75t_L g2164 ( 
.A(n_2089),
.B(n_2014),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2131),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2126),
.Y(n_2166)
);

NOR2x1_ASAP7_75t_L g2167 ( 
.A(n_2138),
.B(n_2008),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2141),
.B(n_2046),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_2100),
.B(n_2082),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2090),
.B(n_2011),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_2100),
.B(n_2042),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2096),
.B(n_2011),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2128),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2131),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2128),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2099),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2099),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2099),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2102),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2085),
.B(n_2042),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2102),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2124),
.B(n_2068),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2085),
.B(n_2029),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2124),
.B(n_2049),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2109),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2097),
.B(n_2075),
.Y(n_2186)
);

AND2x4_ASAP7_75t_L g2187 ( 
.A(n_2100),
.B(n_2083),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2107),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2097),
.B(n_2075),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2121),
.B(n_2043),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_2138),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2108),
.A2(n_2023),
.B(n_2009),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2096),
.B(n_1944),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2097),
.B(n_1944),
.Y(n_2194)
);

OAI21xp33_ASAP7_75t_L g2195 ( 
.A1(n_2105),
.A2(n_2049),
.B(n_2022),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2109),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2109),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_SL g2198 ( 
.A(n_2124),
.Y(n_2198)
);

AOI22x1_ASAP7_75t_SL g2199 ( 
.A1(n_2137),
.A2(n_2036),
.B1(n_2006),
.B2(n_2061),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2143),
.A2(n_2010),
.B1(n_2025),
.B2(n_2035),
.Y(n_2200)
);

NOR2x1p5_ASAP7_75t_SL g2201 ( 
.A(n_2101),
.B(n_1975),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2102),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2104),
.Y(n_2203)
);

OAI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_2151),
.A2(n_2120),
.B(n_2112),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2144),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2147),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2146),
.Y(n_2207)
);

OAI211xp5_ASAP7_75t_L g2208 ( 
.A1(n_2159),
.A2(n_2092),
.B(n_2031),
.C(n_2095),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2170),
.B(n_2142),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2152),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2192),
.B(n_2105),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2153),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2170),
.B(n_2121),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2171),
.B(n_2187),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2172),
.B(n_2121),
.Y(n_2215)
);

NAND2xp33_ASAP7_75t_R g2216 ( 
.A(n_2199),
.B(n_2092),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2172),
.B(n_2134),
.Y(n_2217)
);

CKINVDCx16_ASAP7_75t_R g2218 ( 
.A(n_2198),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_2186),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2146),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2169),
.B(n_2116),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2171),
.B(n_2105),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2148),
.B(n_2112),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2161),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2162),
.Y(n_2225)
);

INVx2_ASAP7_75t_SL g2226 ( 
.A(n_2186),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2158),
.B(n_2134),
.Y(n_2227)
);

NOR3xp33_ASAP7_75t_L g2228 ( 
.A(n_2159),
.B(n_2041),
.C(n_2095),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2169),
.B(n_2116),
.Y(n_2229)
);

NOR4xp25_ASAP7_75t_SL g2230 ( 
.A(n_2191),
.B(n_2140),
.C(n_2074),
.D(n_2014),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2163),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_2176),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2150),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2171),
.B(n_2112),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2177),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2195),
.B(n_2114),
.Y(n_2236)
);

OAI33xp33_ASAP7_75t_L g2237 ( 
.A1(n_2156),
.A2(n_2120),
.A3(n_2106),
.B1(n_2119),
.B2(n_2140),
.B3(n_2086),
.Y(n_2237)
);

NOR3xp33_ASAP7_75t_SL g2238 ( 
.A(n_2184),
.B(n_2048),
.C(n_2067),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2187),
.B(n_2114),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2187),
.B(n_2169),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2158),
.B(n_2098),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_R g2242 ( 
.A(n_2164),
.B(n_2036),
.Y(n_2242)
);

INVxp67_ASAP7_75t_L g2243 ( 
.A(n_2189),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2168),
.B(n_2119),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2167),
.B(n_2116),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2182),
.A2(n_2053),
.B1(n_2114),
.B2(n_2115),
.Y(n_2246)
);

NAND5xp2_ASAP7_75t_SL g2247 ( 
.A(n_2189),
.B(n_2115),
.C(n_2045),
.D(n_2139),
.E(n_2130),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_2149),
.Y(n_2248)
);

AND2x4_ASAP7_75t_L g2249 ( 
.A(n_2180),
.B(n_2154),
.Y(n_2249)
);

NAND2xp33_ASAP7_75t_SL g2250 ( 
.A(n_2149),
.B(n_2036),
.Y(n_2250)
);

INVx1_ASAP7_75t_SL g2251 ( 
.A(n_2188),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2166),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2155),
.B(n_2111),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2173),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_2160),
.Y(n_2255)
);

INVx5_ASAP7_75t_L g2256 ( 
.A(n_2191),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2155),
.B(n_2115),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_2194),
.B(n_2098),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2175),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2213),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2218),
.B(n_2200),
.Y(n_2261)
);

OAI21xp33_ASAP7_75t_L g2262 ( 
.A1(n_2204),
.A2(n_2157),
.B(n_2154),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2244),
.B(n_2251),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2232),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2232),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2244),
.B(n_2157),
.Y(n_2266)
);

OAI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_2208),
.A2(n_2164),
.B(n_2106),
.Y(n_2267)
);

AOI211xp5_ASAP7_75t_L g2268 ( 
.A1(n_2228),
.A2(n_2106),
.B(n_2101),
.C(n_2199),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2235),
.Y(n_2269)
);

OAI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_2211),
.A2(n_2019),
.B1(n_2016),
.B2(n_2117),
.Y(n_2270)
);

NAND2x1_ASAP7_75t_L g2271 ( 
.A(n_2245),
.B(n_2160),
.Y(n_2271)
);

OAI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2238),
.A2(n_2194),
.B1(n_2180),
.B2(n_2145),
.Y(n_2272)
);

NAND2x1p5_ASAP7_75t_L g2273 ( 
.A(n_2256),
.B(n_2038),
.Y(n_2273)
);

OAI222xp33_ASAP7_75t_L g2274 ( 
.A1(n_2236),
.A2(n_2118),
.B1(n_2117),
.B2(n_1995),
.C1(n_2140),
.C2(n_2037),
.Y(n_2274)
);

INVxp67_ASAP7_75t_L g2275 ( 
.A(n_2219),
.Y(n_2275)
);

NAND3xp33_ASAP7_75t_L g2276 ( 
.A(n_2216),
.B(n_2256),
.C(n_2230),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_L g2277 ( 
.A1(n_2247),
.A2(n_2004),
.B1(n_2118),
.B2(n_2117),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2237),
.A2(n_2118),
.B1(n_2004),
.B2(n_2129),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2235),
.Y(n_2279)
);

INVx1_ASAP7_75t_SL g2280 ( 
.A(n_2242),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_2243),
.B(n_2190),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2205),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2214),
.B(n_2245),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2215),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2246),
.A2(n_2129),
.B1(n_2040),
.B2(n_1995),
.Y(n_2285)
);

INVx1_ASAP7_75t_SL g2286 ( 
.A(n_2242),
.Y(n_2286)
);

NAND3xp33_ASAP7_75t_L g2287 ( 
.A(n_2216),
.B(n_2101),
.C(n_2202),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2214),
.B(n_2183),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2206),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2245),
.B(n_2183),
.Y(n_2290)
);

A2O1A1Ixp33_ASAP7_75t_SL g2291 ( 
.A1(n_2248),
.A2(n_2101),
.B(n_2203),
.C(n_2178),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2210),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2221),
.B(n_2145),
.Y(n_2293)
);

OAI21xp33_ASAP7_75t_L g2294 ( 
.A1(n_2223),
.A2(n_2150),
.B(n_2174),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2212),
.Y(n_2295)
);

OAI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2256),
.A2(n_2129),
.B(n_2123),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2224),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2225),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2226),
.B(n_2193),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_2209),
.B(n_2207),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2226),
.B(n_2135),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2261),
.Y(n_2302)
);

INVx2_ASAP7_75t_SL g2303 ( 
.A(n_2283),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2276),
.A2(n_2256),
.B(n_2253),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2261),
.B(n_2255),
.Y(n_2305)
);

NAND3xp33_ASAP7_75t_L g2306 ( 
.A(n_2268),
.B(n_2250),
.C(n_2220),
.Y(n_2306)
);

OAI21xp33_ASAP7_75t_L g2307 ( 
.A1(n_2267),
.A2(n_2207),
.B(n_2220),
.Y(n_2307)
);

AOI31xp33_ASAP7_75t_L g2308 ( 
.A1(n_2280),
.A2(n_2250),
.A3(n_2249),
.B(n_2240),
.Y(n_2308)
);

OAI21xp33_ASAP7_75t_SL g2309 ( 
.A1(n_2277),
.A2(n_2248),
.B(n_2240),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2264),
.Y(n_2310)
);

OAI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2277),
.A2(n_2249),
.B1(n_2229),
.B2(n_2221),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2300),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2275),
.B(n_2299),
.Y(n_2313)
);

INVxp67_ASAP7_75t_SL g2314 ( 
.A(n_2263),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2299),
.B(n_2231),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2260),
.Y(n_2316)
);

OAI32xp33_ASAP7_75t_L g2317 ( 
.A1(n_2262),
.A2(n_2248),
.A3(n_2257),
.B1(n_2241),
.B2(n_2217),
.Y(n_2317)
);

NOR2x1p5_ASAP7_75t_L g2318 ( 
.A(n_2271),
.B(n_2249),
.Y(n_2318)
);

OAI21xp5_ASAP7_75t_L g2319 ( 
.A1(n_2285),
.A2(n_2234),
.B(n_2222),
.Y(n_2319)
);

NOR4xp25_ASAP7_75t_SL g2320 ( 
.A(n_2265),
.B(n_2259),
.C(n_2254),
.D(n_2252),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2281),
.B(n_2227),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2288),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2288),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2269),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2279),
.Y(n_2325)
);

OAI21xp33_ASAP7_75t_L g2326 ( 
.A1(n_2266),
.A2(n_2222),
.B(n_2234),
.Y(n_2326)
);

CKINVDCx16_ASAP7_75t_R g2327 ( 
.A(n_2281),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2282),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2286),
.B(n_2193),
.Y(n_2329)
);

HB1xp67_ASAP7_75t_L g2330 ( 
.A(n_2260),
.Y(n_2330)
);

AOI21xp33_ASAP7_75t_L g2331 ( 
.A1(n_2291),
.A2(n_2287),
.B(n_2298),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2289),
.Y(n_2332)
);

INVxp33_ASAP7_75t_L g2333 ( 
.A(n_2305),
.Y(n_2333)
);

INVxp67_ASAP7_75t_SL g2334 ( 
.A(n_2316),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2330),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2312),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2327),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2327),
.B(n_2283),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_2322),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_SL g2340 ( 
.A(n_2320),
.B(n_2290),
.Y(n_2340)
);

AND4x1_ASAP7_75t_L g2341 ( 
.A(n_2304),
.B(n_2278),
.C(n_2296),
.D(n_2290),
.Y(n_2341)
);

INVxp67_ASAP7_75t_SL g2342 ( 
.A(n_2314),
.Y(n_2342)
);

CKINVDCx16_ASAP7_75t_R g2343 ( 
.A(n_2303),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2322),
.B(n_2284),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2312),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2323),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2323),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2328),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2303),
.B(n_2318),
.Y(n_2349)
);

XOR2x2_ASAP7_75t_L g2350 ( 
.A(n_2306),
.B(n_2273),
.Y(n_2350)
);

OAI221xp5_ASAP7_75t_L g2351 ( 
.A1(n_2309),
.A2(n_2291),
.B1(n_2284),
.B2(n_2273),
.C(n_2272),
.Y(n_2351)
);

XNOR2xp5_ASAP7_75t_L g2352 ( 
.A(n_2302),
.B(n_2270),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2328),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2308),
.B(n_2221),
.Y(n_2354)
);

XOR2xp5_ASAP7_75t_L g2355 ( 
.A(n_2313),
.B(n_2292),
.Y(n_2355)
);

OR2x2_ASAP7_75t_L g2356 ( 
.A(n_2321),
.B(n_2295),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2333),
.B(n_2307),
.Y(n_2357)
);

NOR3x1_ASAP7_75t_L g2358 ( 
.A(n_2334),
.B(n_2311),
.C(n_2315),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2339),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2339),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2340),
.B(n_2331),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2339),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2351),
.A2(n_2318),
.B1(n_2329),
.B2(n_2301),
.Y(n_2363)
);

INVxp67_ASAP7_75t_L g2364 ( 
.A(n_2338),
.Y(n_2364)
);

AOI211xp5_ASAP7_75t_L g2365 ( 
.A1(n_2338),
.A2(n_2317),
.B(n_2309),
.C(n_2319),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2335),
.Y(n_2366)
);

INVx2_ASAP7_75t_SL g2367 ( 
.A(n_2349),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2337),
.B(n_2293),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2337),
.B(n_2332),
.Y(n_2369)
);

OA211x2_ASAP7_75t_L g2370 ( 
.A1(n_2354),
.A2(n_2326),
.B(n_2294),
.C(n_2317),
.Y(n_2370)
);

NOR2xp67_ASAP7_75t_L g2371 ( 
.A(n_2335),
.B(n_2344),
.Y(n_2371)
);

NAND3xp33_ASAP7_75t_L g2372 ( 
.A(n_2361),
.B(n_2342),
.C(n_2336),
.Y(n_2372)
);

AOI32xp33_ASAP7_75t_L g2373 ( 
.A1(n_2365),
.A2(n_2363),
.A3(n_2361),
.B1(n_2357),
.B2(n_2362),
.Y(n_2373)
);

AOI221xp5_ASAP7_75t_SL g2374 ( 
.A1(n_2357),
.A2(n_2355),
.B1(n_2349),
.B2(n_2347),
.C(n_2346),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2359),
.Y(n_2375)
);

AOI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_2369),
.A2(n_2336),
.B1(n_2345),
.B2(n_2355),
.C(n_2353),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2364),
.B(n_2343),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2367),
.B(n_2343),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2371),
.A2(n_2350),
.B(n_2352),
.Y(n_2379)
);

AOI211xp5_ASAP7_75t_L g2380 ( 
.A1(n_2368),
.A2(n_2356),
.B(n_2346),
.C(n_2347),
.Y(n_2380)
);

OAI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2370),
.A2(n_2356),
.B1(n_2229),
.B2(n_2293),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2367),
.A2(n_2350),
.B(n_2352),
.Y(n_2382)
);

OAI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2360),
.A2(n_2229),
.B1(n_2348),
.B2(n_2353),
.Y(n_2383)
);

AOI322xp5_ASAP7_75t_L g2384 ( 
.A1(n_2366),
.A2(n_2345),
.A3(n_2348),
.B1(n_2341),
.B2(n_2332),
.C1(n_2325),
.C2(n_2324),
.Y(n_2384)
);

AOI211xp5_ASAP7_75t_SL g2385 ( 
.A1(n_2378),
.A2(n_2325),
.B(n_2324),
.C(n_2310),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2377),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2372),
.Y(n_2387)
);

AOI222xp33_ASAP7_75t_L g2388 ( 
.A1(n_2376),
.A2(n_2310),
.B1(n_2274),
.B2(n_2358),
.C1(n_2297),
.C2(n_2201),
.Y(n_2388)
);

XOR2xp5_ASAP7_75t_L g2389 ( 
.A(n_2379),
.B(n_2132),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2380),
.B(n_2374),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_2375),
.Y(n_2391)
);

OA22x2_ASAP7_75t_L g2392 ( 
.A1(n_2381),
.A2(n_2233),
.B1(n_2239),
.B2(n_2086),
.Y(n_2392)
);

AOI222xp33_ASAP7_75t_L g2393 ( 
.A1(n_2390),
.A2(n_2387),
.B1(n_2384),
.B2(n_2383),
.C1(n_2386),
.C2(n_2391),
.Y(n_2393)
);

NOR2x1_ASAP7_75t_L g2394 ( 
.A(n_2391),
.B(n_2382),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2385),
.B(n_2373),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2392),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_2389),
.B(n_2233),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2388),
.Y(n_2398)
);

AOI222xp33_ASAP7_75t_L g2399 ( 
.A1(n_2390),
.A2(n_2201),
.B1(n_2123),
.B2(n_1971),
.C1(n_2197),
.C2(n_2196),
.Y(n_2399)
);

INVxp33_ASAP7_75t_L g2400 ( 
.A(n_2391),
.Y(n_2400)
);

AOI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2388),
.A2(n_2239),
.B1(n_2135),
.B2(n_2136),
.Y(n_2401)
);

OA22x2_ASAP7_75t_L g2402 ( 
.A1(n_2396),
.A2(n_2122),
.B1(n_2091),
.B2(n_2179),
.Y(n_2402)
);

AO22x2_ASAP7_75t_L g2403 ( 
.A1(n_2395),
.A2(n_2197),
.B1(n_2196),
.B2(n_2185),
.Y(n_2403)
);

NAND5xp2_ASAP7_75t_L g2404 ( 
.A(n_2393),
.B(n_2088),
.C(n_2054),
.D(n_2136),
.E(n_2135),
.Y(n_2404)
);

NAND3xp33_ASAP7_75t_L g2405 ( 
.A(n_2394),
.B(n_2181),
.C(n_2185),
.Y(n_2405)
);

AOI221xp5_ASAP7_75t_L g2406 ( 
.A1(n_2398),
.A2(n_2123),
.B1(n_2136),
.B2(n_2165),
.C(n_2174),
.Y(n_2406)
);

OAI211xp5_ASAP7_75t_SL g2407 ( 
.A1(n_2399),
.A2(n_2258),
.B(n_2165),
.C(n_2093),
.Y(n_2407)
);

XOR2xp5_ASAP7_75t_L g2408 ( 
.A(n_2403),
.B(n_2400),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2405),
.Y(n_2409)
);

OR4x2_ASAP7_75t_L g2410 ( 
.A(n_2404),
.B(n_2401),
.C(n_2397),
.D(n_1984),
.Y(n_2410)
);

AOI22xp5_ASAP7_75t_L g2411 ( 
.A1(n_2407),
.A2(n_2133),
.B1(n_1971),
.B2(n_2139),
.Y(n_2411)
);

AO22x2_ASAP7_75t_L g2412 ( 
.A1(n_2408),
.A2(n_2402),
.B1(n_2406),
.B2(n_2107),
.Y(n_2412)
);

OAI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2412),
.A2(n_2409),
.B(n_2411),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2413),
.B(n_2410),
.Y(n_2414)
);

CKINVDCx20_ASAP7_75t_R g2415 ( 
.A(n_2413),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2414),
.B(n_2130),
.Y(n_2416)
);

OAI222xp33_ASAP7_75t_L g2417 ( 
.A1(n_2415),
.A2(n_2137),
.B1(n_2088),
.B2(n_2133),
.C1(n_2019),
.C2(n_2107),
.Y(n_2417)
);

CKINVDCx20_ASAP7_75t_R g2418 ( 
.A(n_2416),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2417),
.A2(n_2093),
.B(n_2127),
.Y(n_2419)
);

AOI22xp33_ASAP7_75t_SL g2420 ( 
.A1(n_2418),
.A2(n_2038),
.B1(n_2103),
.B2(n_2137),
.Y(n_2420)
);

OAI221xp5_ASAP7_75t_R g2421 ( 
.A1(n_2420),
.A2(n_2419),
.B1(n_2091),
.B2(n_2122),
.C(n_2130),
.Y(n_2421)
);

OAI31xp33_ASAP7_75t_L g2422 ( 
.A1(n_2421),
.A2(n_2088),
.A3(n_2103),
.B(n_2137),
.Y(n_2422)
);


endmodule