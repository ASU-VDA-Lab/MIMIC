module fake_jpeg_14794_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_63),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_36),
.B1(n_42),
.B2(n_34),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_65),
.B(n_41),
.C(n_40),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_2),
.B(n_3),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_35),
.B1(n_37),
.B2(n_4),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_44),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_80),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_64),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_86),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_47),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_49),
.B1(n_45),
.B2(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_107),
.B1(n_77),
.B2(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_90),
.B1(n_85),
.B2(n_89),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_99),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_103),
.C(n_104),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_94),
.B1(n_82),
.B2(n_11),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_118),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_123),
.C(n_125),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_105),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_13),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_8),
.C(n_9),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_122),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_129),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_126),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_131),
.B(n_15),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_137),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_21),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_140),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_22),
.Y(n_142)
);


endmodule