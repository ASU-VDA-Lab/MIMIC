module real_jpeg_33527_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_0),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_1),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_1),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_1),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_1),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_1),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_1),
.B(n_506),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_2),
.A2(n_19),
.B(n_545),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_2),
.B(n_546),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_3),
.Y(n_144)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_5),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_5),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_39),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_5),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_5),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_5),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_5),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_5),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_6),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_6),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_6),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_7),
.Y(n_236)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_7),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_7),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_8),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_9),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_9),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_9),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_9),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_9),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_9),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_9),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

NAND2x1_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_10),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_10),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_10),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_10),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_10),
.B(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_11),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_12),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_12),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_12),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_12),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g344 ( 
.A(n_12),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_12),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_12),
.B(n_430),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_12),
.B(n_464),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_13),
.Y(n_198)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_14),
.Y(n_248)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_14),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_15),
.Y(n_280)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_15),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_16),
.B(n_238),
.Y(n_237)
);

BUFx24_ASAP7_75t_L g289 ( 
.A(n_16),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_16),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_16),
.B(n_397),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g482 ( 
.A(n_16),
.B(n_57),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_17),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_17),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_17),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_17),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_17),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_17),
.B(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_17),
.B(n_510),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_159),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_157),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_129),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_22),
.B(n_129),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_73),
.C(n_93),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_24),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_50),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_25),
.B(n_51),
.C(n_63),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_36),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_27),
.B(n_120),
.C(n_126),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_27),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_27),
.A2(n_28),
.B1(n_126),
.B2(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_27),
.B(n_190),
.C(n_199),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_27),
.A2(n_28),
.B1(n_200),
.B2(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_31),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_31),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_32),
.Y(n_134)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_35),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_36),
.A2(n_37),
.B(n_133),
.C(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_42),
.C(n_45),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_38),
.B(n_45),
.Y(n_118)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_42),
.B(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_44),
.Y(n_175)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_44),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_46),
.B(n_191),
.C(n_195),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_46),
.B(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XOR2x1_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_63),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.C(n_59),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_75),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_54),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_76),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_78),
.C(n_79),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_76),
.B1(n_78),
.B2(n_99),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_55),
.B(n_342),
.C(n_344),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_55),
.A2(n_76),
.B1(n_342),
.B2(n_382),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_58),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_59),
.B(n_66),
.C(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_59),
.B(n_111),
.C(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_59),
.B(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

XOR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_65),
.A2(n_66),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_65),
.B(n_103),
.C(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_65),
.B(n_222),
.Y(n_351)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_68),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_68),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_68),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_69),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_72),
.Y(n_299)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_73),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.C(n_83),
.Y(n_73)
);

XNOR2x2_ASAP7_75t_SL g202 ( 
.A(n_74),
.B(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_77),
.B(n_83),
.Y(n_203)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_80),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_79),
.A2(n_80),
.B1(n_121),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_121),
.C(n_123),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_80),
.B(n_240),
.Y(n_424)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_82),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.C(n_90),
.Y(n_83)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_84),
.A2(n_150),
.B1(n_151),
.B2(n_155),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_87),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_94),
.B(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_116),
.C(n_119),
.Y(n_94)
);

XNOR2x2_ASAP7_75t_L g204 ( 
.A(n_95),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_114),
.B2(n_115),
.Y(n_95)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_101),
.B(n_104),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_103),
.B(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_104),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.C(n_111),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2x1_ASAP7_75t_SL g171 ( 
.A(n_106),
.B(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_112),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_111),
.A2(n_112),
.B1(n_298),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_117),
.B(n_119),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_122),
.B(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_123),
.B(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_123),
.A2(n_124),
.B1(n_429),
.B2(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_177),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_124),
.B(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_125),
.Y(n_339)
);

INVx8_ASAP7_75t_L g507 ( 
.A(n_125),
.Y(n_507)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_156),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_151),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_151),
.B(n_232),
.C(n_244),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_152),
.A2(n_153),
.B1(n_244),
.B2(n_245),
.Y(n_310)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_154),
.Y(n_398)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21x1_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_256),
.B(n_540),
.Y(n_159)
);

NAND2x1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_209),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_162),
.A2(n_542),
.B(n_543),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_206),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_164),
.B(n_544),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_202),
.C(n_204),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_166),
.B(n_202),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_183),
.C(n_188),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_180),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_169),
.B(n_172),
.Y(n_314)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_176),
.B(n_179),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_177),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_177),
.B(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_177),
.A2(n_230),
.B1(n_336),
.B2(n_337),
.Y(n_379)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_179),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_179),
.A2(n_403),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_180),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_180),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_194),
.Y(n_487)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_206),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_254),
.Y(n_209)
);

NAND2xp67_ASAP7_75t_SL g542 ( 
.A(n_210),
.B(n_254),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_218),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_212),
.B(n_215),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_218),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_231),
.C(n_249),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_220),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.C(n_228),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_221),
.B(n_228),
.Y(n_357)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_226),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_250),
.B1(n_251),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_232),
.A2(n_233),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_237),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_242),
.Y(n_464)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_361),
.B(n_531),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_321),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_318),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_259),
.A2(n_318),
.B1(n_322),
.B2(n_359),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_317),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_260),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_267),
.B(n_312),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_267),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_262),
.A2(n_263),
.B1(n_312),
.B2(n_313),
.Y(n_360)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_269),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_294),
.C(n_308),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_270),
.B(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.C(n_281),
.Y(n_270)
);

XOR2x2_ASAP7_75t_L g410 ( 
.A(n_271),
.B(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_274),
.A2(n_275),
.B(n_277),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_274),
.B(n_282),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_288),
.C(n_290),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_284),
.B(n_332),
.Y(n_331)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_286),
.B(n_343),
.Y(n_342)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_288),
.A2(n_290),
.B1(n_291),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_289),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_289),
.B(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_293),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_295),
.B(n_309),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.C(n_304),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_304),
.Y(n_328)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_303),
.Y(n_427)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_317),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_L g537 ( 
.A(n_318),
.B(n_538),
.C(n_539),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_359),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_322),
.B(n_359),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_352),
.C(n_355),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_324),
.B(n_415),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.C(n_349),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_326),
.B(n_350),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_329),
.B(n_406),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_334),
.B(n_348),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_330),
.A2(n_331),
.B1(n_385),
.B2(n_387),
.Y(n_384)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_340),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_340),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_335),
.A2(n_340),
.B1(n_341),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_343),
.B(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_344),
.B(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_347),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_353),
.B(n_356),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_412),
.C(n_417),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_404),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_363),
.B(n_404),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_383),
.C(n_388),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_364),
.B(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_379),
.C(n_380),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_365),
.B(n_379),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.C(n_373),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g472 ( 
.A(n_367),
.B(n_374),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_369),
.B(n_472),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_R g525 ( 
.A(n_369),
.B(n_472),
.Y(n_525)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_422),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_L g437 ( 
.A(n_384),
.B(n_388),
.Y(n_437)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_385),
.Y(n_387)
);

XOR2x2_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_394),
.C(n_409),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.C(n_403),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_396),
.B1(n_399),
.B2(n_400),
.Y(n_434)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_408),
.C(n_410),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AOI21x1_ASAP7_75t_L g533 ( 
.A1(n_413),
.A2(n_534),
.B(n_535),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_414),
.B(n_416),
.Y(n_534)
);

OAI21x1_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_438),
.B(n_529),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_436),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_420),
.B(n_530),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_423),
.C(n_433),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_421),
.B(n_527),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_423),
.B(n_433),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.C(n_428),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_424),
.A2(n_425),
.B1(n_426),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_429),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_434),
.Y(n_435)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_436),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_522),
.B(n_528),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_478),
.B(n_521),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_468),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_441),
.B(n_468),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_460),
.C(n_465),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_442),
.A2(n_443),
.B1(n_489),
.B2(n_491),
.Y(n_488)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_454),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_449),
.B2(n_453),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_453),
.C(n_454),
.Y(n_470)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_449),
.Y(n_453)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_460),
.A2(n_465),
.B1(n_466),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_460),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_463),
.Y(n_481)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_475),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_473),
.B2(n_474),
.Y(n_469)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_470),
.Y(n_474)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_471),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_474),
.B(n_524),
.C(n_525),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_475),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_492),
.B(n_520),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_488),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_480),
.B(n_488),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.C(n_483),
.Y(n_480)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_517),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_489),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_513),
.B(n_519),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_508),
.B(n_512),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_499),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_499),
.Y(n_512)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_505),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_500),
.B(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_505),
.Y(n_514)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_515),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_518),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_526),
.Y(n_528)
);

O2A1O1Ixp33_ASAP7_75t_SL g531 ( 
.A1(n_532),
.A2(n_533),
.B(n_536),
.C(n_537),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_541),
.Y(n_540)
);


endmodule