module real_jpeg_8936_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_18),
.B(n_50),
.C(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_18),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_8),
.B(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_7),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_23),
.B1(n_37),
.B2(n_38),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_17),
.B(n_25),
.C(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_18),
.B1(n_20),
.B2(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_15),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_80),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_79),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_56),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_13),
.B(n_56),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_31),
.C(n_46),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_14),
.A2(n_46),
.B1(n_88),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_14),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_22),
.B(n_26),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_15),
.A2(n_22),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_17),
.B(n_25),
.C(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_25),
.Y(n_30)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_SL g34 ( 
.A1(n_18),
.A2(n_21),
.B(n_28),
.Y(n_34)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_20),
.A2(n_28),
.B(n_51),
.C(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_28),
.B(n_50),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_31),
.A2(n_32),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_35),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_36),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_37),
.B(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_69),
.B(n_71),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_46),
.B(n_86),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_52),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_74),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_73),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_72),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_84),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_77),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_95),
.C(n_103),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_107),
.B(n_113),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_98),
.B(n_106),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_89),
.B(n_97),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_96),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_100),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_109),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);


endmodule