module fake_aes_7979_n_1150 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1150);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1150;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_1122;
wire n_779;
wire n_993;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1097;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1024;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1063;
wire n_767;
wire n_828;
wire n_1014;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_649;
wire n_526;
wire n_276;
wire n_527;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_666;
wire n_423;
wire n_342;
wire n_621;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_1110;
wire n_327;
wire n_944;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_137), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_19), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_250), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_52), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_48), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_223), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_176), .Y(n_263) );
BUFx8_ASAP7_75t_SL g264 ( .A(n_147), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_114), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_217), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_136), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_20), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_138), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_149), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_12), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_226), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_75), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_125), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_14), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_4), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_102), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_162), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_133), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_120), .Y(n_281) );
BUFx5_ASAP7_75t_L g282 ( .A(n_80), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_98), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_233), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_39), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_55), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_104), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_212), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_154), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_49), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_8), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_109), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_9), .Y(n_293) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_75), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_179), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_178), .Y(n_296) );
INVxp33_ASAP7_75t_L g297 ( .A(n_96), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_62), .Y(n_298) );
BUFx2_ASAP7_75t_SL g299 ( .A(n_34), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_209), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_132), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_187), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_216), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_82), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_157), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_170), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_166), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_215), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_57), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_56), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_202), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_12), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_164), .Y(n_313) );
INVxp33_ASAP7_75t_SL g314 ( .A(n_139), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_229), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_214), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_150), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_69), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_144), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_50), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_25), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g322 ( .A(n_45), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_8), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_210), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_140), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_224), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_85), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_172), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_183), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_106), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_84), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_97), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_186), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_198), .Y(n_335) );
NOR2xp67_ASAP7_75t_L g336 ( .A(n_91), .B(n_41), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_232), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_143), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_19), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_71), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_189), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_35), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_118), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_116), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_167), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_95), .B(n_255), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_201), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_159), .Y(n_348) );
CKINVDCx16_ASAP7_75t_R g349 ( .A(n_55), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_244), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_168), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_128), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_193), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_207), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_88), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_245), .Y(n_356) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_153), .B(n_213), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_190), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_174), .Y(n_359) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_2), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_161), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_219), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_5), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_93), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_42), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_156), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_35), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_243), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_74), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_152), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_185), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_196), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_155), .Y(n_373) );
XOR2xp5_ASAP7_75t_L g374 ( .A(n_27), .B(n_130), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_54), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_1), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_175), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_119), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_158), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_237), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_25), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_103), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_211), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_145), .Y(n_384) );
CKINVDCx14_ASAP7_75t_R g385 ( .A(n_141), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_38), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_282), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_282), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_282), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_326), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_282), .Y(n_391) );
AND2x6_ASAP7_75t_L g392 ( .A(n_346), .B(n_87), .Y(n_392) );
BUFx12f_ASAP7_75t_L g393 ( .A(n_265), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_369), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_326), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_322), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_326), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_282), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_326), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_258), .Y(n_400) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_258), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_282), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_273), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_282), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_309), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_298), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_308), .B(n_0), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_298), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_312), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_308), .B(n_0), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_273), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_349), .B(n_1), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_376), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_376), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_386), .B(n_2), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_269), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_309), .B(n_310), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_257), .B(n_3), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_283), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_283), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_351), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_310), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_342), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_393), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_422), .B(n_337), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_387), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_388), .B(n_269), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
BUFx10_ASAP7_75t_L g431 ( .A(n_392), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_392), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
AOI22xp5_ASAP7_75t_SL g434 ( .A1(n_396), .A2(n_261), .B1(n_323), .B2(n_318), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_422), .B(n_385), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_411), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_389), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_411), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_389), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_417), .B(n_342), .Y(n_445) );
INVx4_ASAP7_75t_L g446 ( .A(n_392), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_392), .A2(n_268), .B1(n_271), .B2(n_260), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_391), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_391), .Y(n_449) );
NOR2x1p5_ASAP7_75t_L g450 ( .A(n_393), .B(n_274), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_392), .A2(n_286), .B1(n_290), .B2(n_277), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_398), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_398), .B(n_338), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_402), .B(n_338), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_392), .Y(n_455) );
NAND2xp33_ASAP7_75t_L g456 ( .A(n_392), .B(n_296), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_394), .B(n_297), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_402), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_394), .B(n_340), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_393), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_412), .B(n_360), .C(n_304), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_395), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_411), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_404), .B(n_358), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_404), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_409), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_417), .B(n_358), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_416), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_417), .B(n_380), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_416), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_415), .B(n_363), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_395), .Y(n_473) );
NOR2x1p5_ASAP7_75t_L g474 ( .A(n_415), .B(n_274), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_457), .B(n_417), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_425), .A2(n_263), .B1(n_270), .B2(n_256), .Y(n_476) );
INVx2_ASAP7_75t_SL g477 ( .A(n_466), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_466), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_445), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_456), .A2(n_410), .B(n_407), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_425), .A2(n_263), .B1(n_270), .B2(n_256), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_460), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_431), .Y(n_483) );
NOR2xp67_ASAP7_75t_SL g484 ( .A(n_432), .B(n_265), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_457), .B(n_410), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_445), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_430), .B(n_259), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_472), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_468), .A2(n_423), .B(n_405), .C(n_416), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_439), .B(n_423), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_430), .B(n_262), .Y(n_493) );
AND2x4_ASAP7_75t_SL g494 ( .A(n_439), .B(n_315), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_468), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_471), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_425), .B(n_266), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_447), .A2(n_418), .B1(n_408), .B2(n_413), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_430), .B(n_278), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_467), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_467), .A2(n_470), .B(n_447), .C(n_451), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_459), .B(n_278), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_430), .B(n_287), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_437), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_430), .B(n_267), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_474), .B(n_287), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_451), .A2(n_418), .B1(n_408), .B2(n_413), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_424), .Y(n_510) );
OR2x6_ASAP7_75t_SL g511 ( .A(n_434), .B(n_276), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_437), .B(n_289), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_437), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_424), .B(n_289), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_438), .B(n_272), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_431), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_428), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_441), .B(n_306), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_461), .B(n_276), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_428), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_441), .A2(n_382), .B(n_380), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_443), .B(n_463), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_461), .B(n_285), .Y(n_523) );
NAND2xp33_ASAP7_75t_L g524 ( .A(n_443), .B(n_307), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_463), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_426), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_426), .B(n_427), .Y(n_527) );
NAND2xp33_ASAP7_75t_L g528 ( .A(n_427), .B(n_331), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_436), .B(n_442), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_438), .B(n_331), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_436), .B(n_347), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_442), .B(n_347), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_450), .A2(n_348), .B1(n_356), .B2(n_315), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_438), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_444), .B(n_355), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_431), .Y(n_536) );
CKINVDCx11_ASAP7_75t_R g537 ( .A(n_434), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_438), .B(n_275), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_453), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_432), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_448), .B(n_314), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_438), .B(n_446), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_446), .A2(n_261), .B1(n_323), .B2(n_318), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_446), .B(n_279), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_449), .B(n_314), .Y(n_545) );
INVx5_ASAP7_75t_L g546 ( .A(n_446), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_452), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_450), .B(n_291), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_454), .A2(n_464), .B1(n_356), .B2(n_361), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_452), .B(n_359), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_464), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_458), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_465), .B(n_359), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_465), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_455), .A2(n_414), .B1(n_406), .B2(n_320), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_431), .B(n_362), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_431), .B(n_366), .Y(n_558) );
AND3x1_ASAP7_75t_SL g559 ( .A(n_511), .B(n_367), .C(n_374), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_553), .A2(n_293), .B(n_328), .C(n_321), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_479), .Y(n_561) );
CKINVDCx8_ASAP7_75t_R g562 ( .A(n_482), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_501), .A2(n_294), .B(n_339), .C(n_332), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_478), .B(n_497), .Y(n_564) );
O2A1O1Ixp5_ASAP7_75t_L g565 ( .A1(n_475), .A2(n_280), .B(n_284), .C(n_281), .Y(n_565) );
BUFx2_ASAP7_75t_L g566 ( .A(n_510), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_502), .A2(n_299), .B1(n_367), .B2(n_365), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_547), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_542), .A2(n_433), .B(n_429), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_537), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_504), .B(n_381), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_487), .B(n_366), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_485), .Y(n_573) );
A2O1A1Ixp33_ASAP7_75t_L g574 ( .A1(n_552), .A2(n_375), .B(n_336), .C(n_406), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_494), .B(n_264), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_514), .B(n_295), .Y(n_576) );
AO21x1_ASAP7_75t_L g577 ( .A1(n_521), .A2(n_292), .B(n_288), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g578 ( .A(n_528), .B(n_370), .C(n_368), .Y(n_578) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_546), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_486), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_555), .Y(n_581) );
OA22x2_ASAP7_75t_L g582 ( .A1(n_476), .A2(n_414), .B1(n_384), .B2(n_371), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_489), .A2(n_462), .B(n_440), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_488), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_508), .B(n_302), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_541), .A2(n_305), .B(n_311), .C(n_303), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_519), .A2(n_384), .B1(n_316), .B2(n_317), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_481), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_493), .A2(n_473), .B(n_319), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_495), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_523), .B(n_313), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_513), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_513), .Y(n_593) );
AOI21x1_ASAP7_75t_L g594 ( .A1(n_493), .A2(n_473), .B(n_357), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_545), .B(n_300), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_499), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_546), .B(n_301), .Y(n_598) );
BUFx2_ASAP7_75t_L g599 ( .A(n_549), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_503), .A2(n_325), .B1(n_327), .B2(n_324), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_545), .A2(n_330), .B(n_333), .C(n_329), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_526), .B(n_334), .Y(n_602) );
BUFx4f_ASAP7_75t_L g603 ( .A(n_548), .Y(n_603) );
BUFx8_ASAP7_75t_L g604 ( .A(n_543), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_506), .Y(n_605) );
O2A1O1Ixp5_ASAP7_75t_L g606 ( .A1(n_507), .A2(n_341), .B(n_343), .C(n_335), .Y(n_606) );
O2A1O1Ixp5_ASAP7_75t_L g607 ( .A1(n_507), .A2(n_345), .B(n_350), .C(n_344), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_534), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_492), .A2(n_400), .B1(n_403), .B2(n_401), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_531), .B(n_377), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_532), .B(n_378), .Y(n_611) );
NOR2xp33_ASAP7_75t_SL g612 ( .A(n_546), .B(n_383), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_491), .A2(n_354), .B(n_364), .C(n_353), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_533), .B(n_4), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_SL g615 ( .A1(n_515), .A2(n_373), .B(n_379), .C(n_372), .Y(n_615) );
AOI22x1_ASAP7_75t_L g616 ( .A1(n_480), .A2(n_403), .B1(n_419), .B2(n_401), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_546), .B(n_400), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_498), .A2(n_400), .B1(n_403), .B2(n_401), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_535), .A2(n_352), .B(n_351), .C(n_390), .Y(n_619) );
CKINVDCx6p67_ASAP7_75t_R g620 ( .A(n_512), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_540), .B(n_400), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_540), .B(n_352), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_515), .A2(n_473), .B(n_403), .Y(n_623) );
BUFx12f_ASAP7_75t_L g624 ( .A(n_551), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_498), .A2(n_401), .B1(n_419), .B2(n_403), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_525), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_550), .B(n_5), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_554), .A2(n_390), .B(n_9), .C(n_6), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_509), .B(n_7), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_522), .Y(n_630) );
NOR2xp33_ASAP7_75t_R g631 ( .A(n_524), .B(n_10), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_556), .B(n_401), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_517), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_539), .B(n_10), .Y(n_634) );
NAND2xp33_ASAP7_75t_L g635 ( .A(n_483), .B(n_401), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_483), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_500), .B(n_11), .Y(n_637) );
INVx5_ASAP7_75t_L g638 ( .A(n_534), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_538), .A2(n_390), .B(n_14), .C(n_11), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_483), .B(n_401), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_520), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_556), .B(n_403), .Y(n_642) );
NAND2x1_ASAP7_75t_SL g643 ( .A(n_509), .B(n_13), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_518), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_538), .B(n_419), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_544), .A2(n_420), .B(n_419), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_544), .A2(n_17), .B(n_15), .C(n_16), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_SL g648 ( .A1(n_484), .A2(n_421), .B(n_420), .C(n_419), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_505), .B(n_17), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_483), .B(n_420), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_530), .A2(n_18), .B(n_20), .C(n_21), .Y(n_651) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_516), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_557), .B(n_420), .Y(n_653) );
INVx5_ASAP7_75t_L g654 ( .A(n_516), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_558), .A2(n_420), .B1(n_421), .B2(n_397), .Y(n_655) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_516), .A2(n_469), .B(n_435), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_516), .B(n_18), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_536), .A2(n_421), .B1(n_420), .B2(n_399), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_536), .B(n_21), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_536), .A2(n_421), .B1(n_397), .B2(n_399), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_490), .B(n_22), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_490), .B(n_22), .Y(n_662) );
NAND2xp33_ASAP7_75t_L g663 ( .A(n_483), .B(n_397), .Y(n_663) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_546), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_502), .A2(n_397), .B1(n_399), .B2(n_24), .Y(n_665) );
O2A1O1Ixp5_ASAP7_75t_L g666 ( .A1(n_475), .A2(n_469), .B(n_435), .C(n_131), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_477), .B(n_397), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_553), .A2(n_399), .B(n_397), .C(n_469), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_490), .B(n_23), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_542), .A2(n_469), .B(n_435), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_479), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_502), .A2(n_399), .B1(n_26), .B2(n_27), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_490), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_501), .A2(n_28), .B(n_29), .C(n_30), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_477), .B(n_435), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_478), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_478), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_479), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_477), .B(n_435), .Y(n_679) );
AO31x2_ASAP7_75t_L g680 ( .A1(n_625), .A2(n_618), .A3(n_600), .B(n_577), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_588), .A2(n_469), .B1(n_31), .B2(n_32), .Y(n_681) );
AOI22x1_ASAP7_75t_SL g682 ( .A1(n_570), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_682) );
AO31x2_ASAP7_75t_L g683 ( .A1(n_625), .A2(n_33), .A3(n_34), .B(n_36), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_676), .B(n_33), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_565), .A2(n_90), .B(n_89), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_590), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_677), .B(n_37), .Y(n_687) );
AO21x1_ASAP7_75t_L g688 ( .A1(n_600), .A2(n_94), .B(n_92), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_673), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_568), .Y(n_690) );
INVx4_ASAP7_75t_L g691 ( .A(n_654), .Y(n_691) );
INVx2_ASAP7_75t_SL g692 ( .A(n_603), .Y(n_692) );
INVx3_ASAP7_75t_SL g693 ( .A(n_620), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_627), .A2(n_40), .B(n_43), .C(n_44), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_595), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_597), .Y(n_696) );
NOR2xp67_ASAP7_75t_L g697 ( .A(n_654), .B(n_99), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_574), .A2(n_44), .B(n_45), .C(n_46), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_613), .A2(n_46), .B(n_47), .C(n_49), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_562), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_632), .A2(n_101), .B(n_100), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_654), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_662), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_L g705 ( .A1(n_586), .A2(n_51), .B(n_52), .C(n_53), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_637), .A2(n_53), .B(n_54), .C(n_57), .Y(n_706) );
O2A1O1Ixp5_ASAP7_75t_SL g707 ( .A1(n_672), .A2(n_173), .B(n_253), .C(n_252), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_581), .Y(n_708) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_566), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_599), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_710) );
OAI21x1_ASAP7_75t_L g711 ( .A1(n_616), .A2(n_171), .B(n_251), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_561), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_654), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_649), .A2(n_59), .B(n_61), .C(n_62), .Y(n_714) );
BUFx4_ASAP7_75t_R g715 ( .A(n_559), .Y(n_715) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_636), .Y(n_716) );
BUFx8_ASAP7_75t_L g717 ( .A(n_624), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_61), .B1(n_63), .B2(n_64), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_603), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_572), .B(n_63), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g721 ( .A1(n_628), .A2(n_64), .B(n_65), .C(n_66), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_602), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_722) );
BUFx3_ASAP7_75t_L g723 ( .A(n_604), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_569), .A2(n_180), .B(n_249), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_602), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g726 ( .A1(n_642), .A2(n_181), .B(n_248), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_630), .A2(n_68), .B1(n_70), .B2(n_72), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_575), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_573), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_666), .A2(n_177), .B(n_247), .Y(n_730) );
BUFx2_ASAP7_75t_L g731 ( .A(n_631), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_675), .A2(n_169), .B(n_246), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_567), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_661), .A2(n_73), .B(n_74), .C(n_76), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_633), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_679), .A2(n_182), .B(n_241), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_640), .A2(n_165), .B(n_240), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_580), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g739 ( .A1(n_669), .A2(n_73), .B(n_76), .C(n_77), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_612), .B(n_78), .Y(n_740) );
AO32x2_ASAP7_75t_L g741 ( .A1(n_665), .A2(n_78), .A3(n_79), .B1(n_80), .B2(n_81), .Y(n_741) );
AO31x2_ASAP7_75t_L g742 ( .A1(n_655), .A2(n_79), .A3(n_81), .B(n_82), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_591), .B(n_83), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g744 ( .A(n_579), .B(n_83), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g745 ( .A1(n_639), .A2(n_84), .B(n_85), .C(n_86), .Y(n_745) );
OA21x2_ASAP7_75t_L g746 ( .A1(n_668), .A2(n_105), .B(n_107), .Y(n_746) );
NOR2x1_ASAP7_75t_R g747 ( .A(n_629), .B(n_108), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_584), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_650), .A2(n_110), .B(n_111), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_582), .A2(n_112), .B1(n_113), .B2(n_115), .Y(n_750) );
BUFx2_ASAP7_75t_L g751 ( .A(n_622), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_579), .Y(n_752) );
AO32x2_ASAP7_75t_L g753 ( .A1(n_672), .A2(n_117), .A3(n_121), .B1(n_122), .B2(n_123), .Y(n_753) );
AO31x2_ASAP7_75t_L g754 ( .A1(n_655), .A2(n_124), .A3(n_126), .B(n_127), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_560), .B(n_129), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_601), .A2(n_134), .B(n_135), .Y(n_756) );
OR2x6_ASAP7_75t_L g757 ( .A(n_582), .B(n_142), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_644), .A2(n_146), .B1(n_148), .B2(n_151), .Y(n_758) );
BUFx3_ASAP7_75t_L g759 ( .A(n_664), .Y(n_759) );
OR2x6_ASAP7_75t_L g760 ( .A(n_664), .B(n_160), .Y(n_760) );
AO21x2_ASAP7_75t_L g761 ( .A1(n_594), .A2(n_163), .B(n_184), .Y(n_761) );
BUFx12f_ASAP7_75t_L g762 ( .A(n_638), .Y(n_762) );
BUFx3_ASAP7_75t_L g763 ( .A(n_605), .Y(n_763) );
BUFx12f_ASAP7_75t_L g764 ( .A(n_638), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_621), .A2(n_191), .B(n_192), .Y(n_765) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_636), .Y(n_766) );
OA21x2_ASAP7_75t_L g767 ( .A1(n_643), .A2(n_194), .B(n_195), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_L g768 ( .A1(n_651), .A2(n_197), .B(n_199), .C(n_200), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g769 ( .A1(n_587), .A2(n_203), .B(n_205), .C(n_206), .Y(n_769) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_636), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g771 ( .A(n_652), .B(n_208), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_638), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_678), .Y(n_773) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_652), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_671), .Y(n_775) );
BUFx12f_ASAP7_75t_L g776 ( .A(n_652), .Y(n_776) );
NAND2x1_ASAP7_75t_L g777 ( .A(n_608), .B(n_218), .Y(n_777) );
AO21x2_ASAP7_75t_L g778 ( .A1(n_648), .A2(n_220), .B(n_221), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_571), .A2(n_222), .B1(n_225), .B2(n_227), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g780 ( .A1(n_674), .A2(n_228), .B(n_230), .C(n_231), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_653), .A2(n_234), .B(n_235), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_L g782 ( .A1(n_563), .A2(n_236), .B(n_238), .C(n_239), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_610), .A2(n_254), .B(n_611), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_583), .A2(n_623), .B(n_635), .Y(n_784) );
OAI21x1_ASAP7_75t_L g785 ( .A1(n_646), .A2(n_660), .B(n_645), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_L g786 ( .A1(n_647), .A2(n_596), .B(n_615), .C(n_576), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_645), .A2(n_667), .B(n_626), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_634), .A2(n_585), .B1(n_608), .B2(n_578), .Y(n_788) );
A2O1A1Ixp33_ASAP7_75t_L g789 ( .A1(n_606), .A2(n_607), .B(n_657), .C(n_659), .Y(n_789) );
O2A1O1Ixp33_ASAP7_75t_L g790 ( .A1(n_619), .A2(n_598), .B(n_617), .C(n_593), .Y(n_790) );
A2O1A1Ixp33_ASAP7_75t_L g791 ( .A1(n_589), .A2(n_592), .B(n_609), .C(n_658), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_660), .Y(n_792) );
OAI21x1_ASAP7_75t_L g793 ( .A1(n_663), .A2(n_656), .B(n_616), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_676), .Y(n_794) );
NAND2x1p5_ASAP7_75t_L g795 ( .A(n_603), .B(n_676), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_588), .B(n_476), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_676), .B(n_490), .Y(n_797) );
INVx4_ASAP7_75t_L g798 ( .A(n_654), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g799 ( .A1(n_627), .A2(n_565), .B(n_564), .C(n_613), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_670), .A2(n_529), .B(n_527), .Y(n_800) );
NOR2x1_ASAP7_75t_SL g801 ( .A(n_654), .B(n_579), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_695), .B(n_696), .Y(n_802) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_800), .A2(n_799), .B(n_792), .Y(n_803) );
OR2x6_ASAP7_75t_L g804 ( .A(n_760), .B(n_795), .Y(n_804) );
AO221x2_ASAP7_75t_L g805 ( .A1(n_718), .A2(n_725), .B1(n_722), .B2(n_727), .C(n_756), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_707), .A2(n_785), .B(n_685), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_738), .B(n_748), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_686), .Y(n_808) );
NAND2x1p5_ASAP7_75t_L g809 ( .A(n_691), .B(n_798), .Y(n_809) );
BUFx6f_ASAP7_75t_L g810 ( .A(n_776), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_702), .Y(n_811) );
INVx3_ASAP7_75t_L g812 ( .A(n_691), .Y(n_812) );
OR2x6_ASAP7_75t_L g813 ( .A(n_760), .B(n_692), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_789), .A2(n_787), .B(n_791), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_712), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_729), .Y(n_816) );
INVx5_ASAP7_75t_L g817 ( .A(n_760), .Y(n_817) );
OA21x2_ASAP7_75t_L g818 ( .A1(n_701), .A2(n_726), .B(n_756), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_709), .B(n_693), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_751), .B(n_794), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_735), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_773), .B(n_775), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_684), .B(n_689), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_790), .A2(n_720), .B(n_704), .Y(n_824) );
OA21x2_ASAP7_75t_L g825 ( .A1(n_688), .A2(n_768), .B(n_780), .Y(n_825) );
O2A1O1Ixp33_ASAP7_75t_L g826 ( .A1(n_734), .A2(n_739), .B(n_694), .C(n_699), .Y(n_826) );
OAI21x1_ASAP7_75t_L g827 ( .A1(n_771), .A2(n_777), .B(n_724), .Y(n_827) );
BUFx3_ASAP7_75t_L g828 ( .A(n_717), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_689), .B(n_763), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_690), .Y(n_830) );
BUFx2_ASAP7_75t_L g831 ( .A(n_762), .Y(n_831) );
INVx3_ASAP7_75t_L g832 ( .A(n_798), .Y(n_832) );
INVx4_ASAP7_75t_L g833 ( .A(n_764), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_708), .Y(n_834) );
A2O1A1Ixp33_ASAP7_75t_L g835 ( .A1(n_782), .A2(n_705), .B(n_721), .C(n_745), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_723), .A2(n_687), .B1(n_755), .B2(n_788), .Y(n_836) );
NOR2xp67_ASAP7_75t_L g837 ( .A(n_700), .B(n_728), .Y(n_837) );
BUFx2_ASAP7_75t_L g838 ( .A(n_759), .Y(n_838) );
AOI22xp33_ASAP7_75t_SL g839 ( .A1(n_682), .A2(n_744), .B1(n_698), .B2(n_747), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_683), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_683), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_680), .B(n_747), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_779), .A2(n_681), .B1(n_750), .B2(n_703), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_680), .B(n_772), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_761), .A2(n_767), .B(n_766), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_680), .B(n_772), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_713), .B(n_801), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_752), .Y(n_848) );
BUFx4_ASAP7_75t_SL g849 ( .A(n_717), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_740), .A2(n_752), .B1(n_758), .B2(n_779), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_742), .Y(n_851) );
OR2x4_ASAP7_75t_L g852 ( .A(n_715), .B(n_716), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_706), .B(n_714), .Y(n_853) );
AND2x4_ASAP7_75t_L g854 ( .A(n_697), .B(n_716), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_774), .B(n_770), .Y(n_855) );
OA21x2_ASAP7_75t_L g856 ( .A1(n_781), .A2(n_769), .B(n_732), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_770), .B(n_742), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_770), .B(n_736), .Y(n_858) );
OA21x2_ASAP7_75t_L g859 ( .A1(n_765), .A2(n_749), .B(n_737), .Y(n_859) );
INVx2_ASAP7_75t_SL g860 ( .A(n_754), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_754), .B(n_746), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_741), .A2(n_710), .B1(n_760), .B2(n_757), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_753), .B(n_778), .Y(n_863) );
AO21x2_ASAP7_75t_L g864 ( .A1(n_778), .A2(n_685), .B(n_792), .Y(n_864) );
OA21x2_ASAP7_75t_L g865 ( .A1(n_793), .A2(n_730), .B(n_711), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_695), .B(n_696), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g867 ( .A1(n_800), .A2(n_600), .B(n_799), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_731), .A2(n_604), .B1(n_434), .B2(n_494), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g869 ( .A1(n_786), .A2(n_799), .B(n_743), .C(n_627), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_695), .B(n_696), .Y(n_870) );
OR2x2_ASAP7_75t_L g871 ( .A(n_797), .B(n_490), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_712), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_695), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_712), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_695), .B(n_696), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_712), .Y(n_876) );
OR2x2_ASAP7_75t_L g877 ( .A(n_797), .B(n_490), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_797), .B(n_490), .Y(n_878) );
OAI221xp5_ASAP7_75t_SL g879 ( .A1(n_710), .A2(n_481), .B1(n_476), .B2(n_567), .C(n_533), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_717), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_796), .A2(n_604), .B1(n_733), .B2(n_599), .Y(n_881) );
NAND2x1p5_ASAP7_75t_L g882 ( .A(n_691), .B(n_798), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_695), .B(n_696), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_695), .B(n_696), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_695), .B(n_696), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_800), .A2(n_600), .B(n_799), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_695), .B(n_696), .Y(n_887) );
BUFx8_ASAP7_75t_L g888 ( .A(n_700), .Y(n_888) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_800), .A2(n_784), .B(n_783), .Y(n_889) );
OA21x2_ASAP7_75t_L g890 ( .A1(n_793), .A2(n_730), .B(n_711), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_712), .Y(n_891) );
OAI21xp5_ASAP7_75t_L g892 ( .A1(n_800), .A2(n_600), .B(n_799), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_712), .Y(n_893) );
AND2x4_ASAP7_75t_L g894 ( .A(n_692), .B(n_719), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_695), .B(n_696), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_695), .B(n_696), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_712), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_844), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_844), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_846), .Y(n_900) );
NOR2x1_ASAP7_75t_SL g901 ( .A(n_813), .B(n_804), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_846), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_813), .A2(n_804), .B1(n_862), .B2(n_817), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_808), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_802), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_851), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_805), .A2(n_839), .B1(n_868), .B2(n_881), .Y(n_907) );
BUFx2_ASAP7_75t_L g908 ( .A(n_817), .Y(n_908) );
AOI22xp5_ASAP7_75t_SL g909 ( .A1(n_828), .A2(n_880), .B1(n_849), .B2(n_833), .Y(n_909) );
BUFx2_ASAP7_75t_L g910 ( .A(n_817), .Y(n_910) );
INVx2_ASAP7_75t_SL g911 ( .A(n_810), .Y(n_911) );
AND2x4_ASAP7_75t_L g912 ( .A(n_813), .B(n_817), .Y(n_912) );
NOR2x1_ASAP7_75t_R g913 ( .A(n_833), .B(n_831), .Y(n_913) );
NAND3xp33_ASAP7_75t_L g914 ( .A(n_869), .B(n_840), .C(n_841), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_815), .B(n_816), .Y(n_915) );
OAI21xp5_ASAP7_75t_L g916 ( .A1(n_835), .A2(n_824), .B(n_826), .Y(n_916) );
INVx4_ASAP7_75t_L g917 ( .A(n_810), .Y(n_917) );
OR2x2_ASAP7_75t_L g918 ( .A(n_822), .B(n_842), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_872), .B(n_874), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_878), .B(n_871), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_822), .B(n_842), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_877), .B(n_811), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_807), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_879), .B(n_819), .Y(n_924) );
OR2x6_ASAP7_75t_L g925 ( .A(n_809), .B(n_882), .Y(n_925) );
OA21x2_ASAP7_75t_L g926 ( .A1(n_861), .A2(n_803), .B(n_814), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_873), .B(n_866), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_847), .B(n_812), .Y(n_928) );
INVxp67_ASAP7_75t_SL g929 ( .A(n_866), .Y(n_929) );
AO21x2_ASAP7_75t_L g930 ( .A1(n_806), .A2(n_803), .B(n_889), .Y(n_930) );
OR2x6_ASAP7_75t_L g931 ( .A(n_809), .B(n_882), .Y(n_931) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_829), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_870), .B(n_887), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_876), .B(n_891), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_870), .B(n_885), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g936 ( .A(n_836), .B(n_886), .C(n_867), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_857), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_823), .A2(n_853), .B1(n_843), .B2(n_820), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_857), .Y(n_939) );
OA21x2_ASAP7_75t_L g940 ( .A1(n_845), .A2(n_892), .B(n_867), .Y(n_940) );
NAND2x1_ASAP7_75t_L g941 ( .A(n_854), .B(n_860), .Y(n_941) );
OR2x2_ASAP7_75t_L g942 ( .A(n_875), .B(n_884), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_875), .Y(n_943) );
INVx3_ASAP7_75t_L g944 ( .A(n_812), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_853), .A2(n_884), .B1(n_896), .B2(n_895), .C(n_887), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_883), .B(n_885), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_893), .B(n_897), .Y(n_947) );
INVx3_ASAP7_75t_L g948 ( .A(n_832), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_830), .B(n_834), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_821), .B(n_896), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_883), .B(n_895), .Y(n_951) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_838), .Y(n_952) );
BUFx3_ASAP7_75t_L g953 ( .A(n_832), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_848), .B(n_892), .Y(n_954) );
AO21x2_ASAP7_75t_L g955 ( .A1(n_886), .A2(n_863), .B(n_864), .Y(n_955) );
INVx3_ASAP7_75t_L g956 ( .A(n_827), .Y(n_956) );
CKINVDCx11_ASAP7_75t_R g957 ( .A(n_894), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_865), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_855), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_855), .B(n_850), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_858), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_837), .B(n_852), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_858), .Y(n_963) );
INVx5_ASAP7_75t_L g964 ( .A(n_888), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_825), .B(n_843), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_825), .B(n_818), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_890), .Y(n_967) );
INVx3_ASAP7_75t_L g968 ( .A(n_859), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_906), .Y(n_969) );
INVx2_ASAP7_75t_L g970 ( .A(n_958), .Y(n_970) );
AND2x4_ASAP7_75t_L g971 ( .A(n_961), .B(n_859), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_951), .B(n_856), .Y(n_972) );
AND2x4_ASAP7_75t_L g973 ( .A(n_961), .B(n_856), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_951), .B(n_965), .Y(n_974) );
BUFx2_ASAP7_75t_L g975 ( .A(n_908), .Y(n_975) );
BUFx3_ASAP7_75t_L g976 ( .A(n_925), .Y(n_976) );
BUFx2_ASAP7_75t_L g977 ( .A(n_908), .Y(n_977) );
OAI31xp33_ASAP7_75t_L g978 ( .A1(n_907), .A2(n_924), .A3(n_903), .B(n_942), .Y(n_978) );
INVx3_ASAP7_75t_L g979 ( .A(n_941), .Y(n_979) );
NOR2x1_ASAP7_75t_L g980 ( .A(n_925), .B(n_931), .Y(n_980) );
AND2x2_ASAP7_75t_SL g981 ( .A(n_912), .B(n_910), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_918), .B(n_921), .Y(n_982) );
NOR2x1_ASAP7_75t_L g983 ( .A(n_925), .B(n_931), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_929), .A2(n_942), .B1(n_938), .B2(n_945), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_918), .B(n_921), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_937), .B(n_939), .Y(n_986) );
AO21x2_ASAP7_75t_L g987 ( .A1(n_916), .A2(n_967), .B(n_936), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_939), .B(n_959), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_950), .B(n_898), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_950), .B(n_899), .Y(n_990) );
AND2x4_ASAP7_75t_L g991 ( .A(n_963), .B(n_899), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_933), .A2(n_946), .B1(n_935), .B2(n_943), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_905), .B(n_923), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_900), .Y(n_994) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_920), .B(n_957), .Y(n_995) );
INVx4_ASAP7_75t_L g996 ( .A(n_925), .Y(n_996) );
NOR2x1_ASAP7_75t_SL g997 ( .A(n_931), .B(n_953), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_900), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_902), .B(n_960), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_932), .B(n_954), .Y(n_1000) );
NOR2x1_ASAP7_75t_SL g1001 ( .A(n_931), .B(n_953), .Y(n_1001) );
OR2x2_ASAP7_75t_L g1002 ( .A(n_954), .B(n_960), .Y(n_1002) );
BUFx3_ASAP7_75t_L g1003 ( .A(n_928), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_949), .B(n_947), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_949), .B(n_919), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_927), .B(n_904), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_915), .B(n_934), .Y(n_1007) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_910), .Y(n_1008) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_912), .Y(n_1009) );
INVx2_ASAP7_75t_L g1010 ( .A(n_968), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_912), .A2(n_952), .B1(n_922), .B2(n_962), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_1002), .B(n_914), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_969), .Y(n_1013) );
AND2x4_ASAP7_75t_SL g1014 ( .A(n_996), .B(n_928), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_1004), .B(n_947), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_974), .B(n_966), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_974), .B(n_966), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_969), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_970), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_1000), .B(n_926), .Y(n_1020) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_972), .B(n_956), .Y(n_1021) );
INVx3_ASAP7_75t_L g1022 ( .A(n_979), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_982), .B(n_926), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_975), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_982), .B(n_985), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_999), .B(n_926), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_999), .B(n_940), .Y(n_1027) );
INVx1_ASAP7_75t_SL g1028 ( .A(n_1005), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_972), .B(n_940), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_985), .B(n_955), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_989), .B(n_940), .Y(n_1031) );
INVx1_ASAP7_75t_SL g1032 ( .A(n_1005), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_989), .B(n_940), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_990), .B(n_955), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_990), .B(n_955), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_1007), .B(n_928), .Y(n_1036) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_977), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1007), .B(n_917), .Y(n_1038) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_995), .B(n_913), .Y(n_1039) );
INVx2_ASAP7_75t_SL g1040 ( .A(n_980), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_991), .B(n_930), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_992), .B(n_917), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_992), .B(n_917), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_991), .B(n_930), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1034), .B(n_988), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1013), .Y(n_1046) );
NOR2xp67_ASAP7_75t_L g1047 ( .A(n_1022), .B(n_996), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1013), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1016), .B(n_987), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1019), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_1028), .B(n_987), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1018), .Y(n_1052) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_1032), .B(n_987), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_1030), .B(n_987), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1016), .B(n_971), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1034), .B(n_988), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1018), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1017), .B(n_971), .Y(n_1058) );
NAND4xp75_ASAP7_75t_L g1059 ( .A(n_1039), .B(n_980), .C(n_983), .D(n_978), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1060 ( .A(n_1030), .B(n_986), .Y(n_1060) );
BUFx2_ASAP7_75t_L g1061 ( .A(n_1037), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1017), .B(n_971), .Y(n_1062) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_1025), .B(n_986), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1027), .B(n_971), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1027), .B(n_973), .Y(n_1065) );
INVx2_ASAP7_75t_SL g1066 ( .A(n_1037), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1035), .B(n_994), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1031), .B(n_973), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1031), .B(n_973), .Y(n_1069) );
INVx3_ASAP7_75t_L g1070 ( .A(n_1022), .Y(n_1070) );
INVx2_ASAP7_75t_SL g1071 ( .A(n_1037), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1023), .B(n_998), .Y(n_1072) );
NOR2x1_ASAP7_75t_L g1073 ( .A(n_1042), .B(n_983), .Y(n_1073) );
INVx3_ASAP7_75t_L g1074 ( .A(n_1022), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1064), .B(n_1033), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1049), .B(n_1033), .Y(n_1076) );
AND2x4_ASAP7_75t_L g1077 ( .A(n_1065), .B(n_1021), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1046), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1064), .B(n_1029), .Y(n_1079) );
INVx1_ASAP7_75t_SL g1080 ( .A(n_1063), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1065), .B(n_1029), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1068), .B(n_1041), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1049), .B(n_1012), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1046), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_1063), .B(n_909), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1048), .Y(n_1086) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_1061), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1048), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1050), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1068), .B(n_1041), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1069), .B(n_1044), .Y(n_1091) );
NOR2x1p5_ASAP7_75t_SL g1092 ( .A(n_1059), .B(n_1010), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1060), .B(n_1023), .Y(n_1093) );
O2A1O1Ixp33_ASAP7_75t_SL g1094 ( .A1(n_1066), .A2(n_1011), .B(n_1040), .C(n_1043), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1052), .Y(n_1095) );
INVx3_ASAP7_75t_L g1096 ( .A(n_1070), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_1060), .B(n_1020), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1067), .B(n_1012), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1052), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1057), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1067), .B(n_1026), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1057), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1080), .B(n_1045), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1089), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1079), .B(n_1069), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1097), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1098), .B(n_1045), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1083), .B(n_1056), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1076), .B(n_1051), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1093), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1079), .B(n_1055), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g1112 ( .A(n_1094), .B(n_1073), .C(n_1054), .Y(n_1112) );
OAI21xp33_ASAP7_75t_L g1113 ( .A1(n_1092), .A2(n_1058), .B(n_1062), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1101), .B(n_1056), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1078), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1078), .Y(n_1116) );
AOI31xp33_ASAP7_75t_SL g1117 ( .A1(n_1085), .A2(n_1038), .A3(n_1053), .B(n_1051), .Y(n_1117) );
AOI322xp5_ASAP7_75t_L g1118 ( .A1(n_1113), .A2(n_1075), .A3(n_1081), .B1(n_1082), .B2(n_1090), .C1(n_1091), .C2(n_1077), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_1106), .A2(n_1087), .B1(n_1077), .B2(n_1062), .Y(n_1119) );
OAI32xp33_ASAP7_75t_L g1120 ( .A1(n_1112), .A2(n_1087), .A3(n_1096), .B1(n_1072), .B2(n_1024), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_1107), .B(n_1077), .Y(n_1121) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_1117), .A2(n_1096), .B1(n_1061), .B2(n_1071), .C(n_1066), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1106), .B(n_1084), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1104), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_1110), .A2(n_1003), .B1(n_1021), .B2(n_1026), .Y(n_1125) );
OAI31xp33_ASAP7_75t_L g1126 ( .A1(n_1105), .A2(n_984), .A3(n_1096), .B(n_1014), .Y(n_1126) );
NAND3xp33_ASAP7_75t_L g1127 ( .A(n_1126), .B(n_964), .C(n_1116), .Y(n_1127) );
NAND2xp5_ASAP7_75t_SL g1128 ( .A(n_1118), .B(n_1047), .Y(n_1128) );
O2A1O1Ixp33_ASAP7_75t_L g1129 ( .A1(n_1120), .A2(n_1103), .B(n_1109), .C(n_911), .Y(n_1129) );
AOI222xp33_ASAP7_75t_L g1130 ( .A1(n_1122), .A2(n_1092), .B1(n_1116), .B2(n_1115), .C1(n_1108), .C2(n_1114), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_1128), .A2(n_1123), .B1(n_1121), .B2(n_1125), .C(n_1124), .Y(n_1131) );
OAI211xp5_ASAP7_75t_SL g1132 ( .A1(n_1130), .A2(n_1119), .B(n_1123), .C(n_1006), .Y(n_1132) );
OA211x2_ASAP7_75t_L g1133 ( .A1(n_1127), .A2(n_1036), .B(n_901), .C(n_993), .Y(n_1133) );
NAND5xp2_ASAP7_75t_L g1134 ( .A(n_1129), .B(n_1009), .C(n_1008), .D(n_1111), .E(n_993), .Y(n_1134) );
AOI22xp5_ASAP7_75t_L g1135 ( .A1(n_1132), .A2(n_981), .B1(n_1070), .B2(n_1074), .Y(n_1135) );
OAI211xp5_ASAP7_75t_L g1136 ( .A1(n_1131), .A2(n_976), .B(n_1074), .C(n_1070), .Y(n_1136) );
AND3x2_ASAP7_75t_L g1137 ( .A(n_1133), .B(n_997), .C(n_1001), .Y(n_1137) );
XNOR2xp5_ASAP7_75t_L g1138 ( .A(n_1137), .B(n_1134), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1135), .Y(n_1139) );
CKINVDCx20_ASAP7_75t_R g1140 ( .A(n_1136), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_1140), .A2(n_976), .B1(n_981), .B2(n_1014), .Y(n_1141) );
AND4x1_ASAP7_75t_L g1142 ( .A(n_1139), .B(n_1015), .C(n_1100), .D(n_1099), .Y(n_1142) );
XNOR2xp5_ASAP7_75t_L g1143 ( .A(n_1141), .B(n_1138), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1142), .Y(n_1144) );
OAI22xp5_ASAP7_75t_SL g1145 ( .A1(n_1143), .A2(n_976), .B1(n_1074), .B2(n_979), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_1144), .A2(n_948), .B1(n_944), .B2(n_1095), .C(n_1084), .Y(n_1146) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1145), .Y(n_1147) );
AOI222xp33_ASAP7_75t_L g1148 ( .A1(n_1146), .A2(n_1102), .B1(n_1100), .B2(n_1095), .C1(n_1086), .C2(n_1088), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1147), .B(n_1086), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_1149), .A2(n_1148), .B1(n_1022), .B2(n_1021), .Y(n_1150) );
endmodule