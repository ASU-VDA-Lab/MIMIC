module fake_jpeg_2878_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_28),
.B1(n_24),
.B2(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_59),
.B1(n_55),
.B2(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_28),
.B1(n_24),
.B2(n_29),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_31),
.B1(n_22),
.B2(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_23),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_31),
.B1(n_26),
.B2(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_31),
.B1(n_26),
.B2(n_17),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_20),
.B(n_33),
.C(n_34),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_27),
.B(n_19),
.C(n_21),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_81),
.B(n_64),
.C(n_96),
.Y(n_100)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_85),
.Y(n_104)
);

AO22x2_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_47),
.B1(n_40),
.B2(n_37),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_71),
.B(n_69),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_65),
.B(n_66),
.Y(n_106)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_27),
.B1(n_51),
.B2(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_89),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_27),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_95),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_93),
.B1(n_55),
.B2(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_53),
.B(n_19),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_98),
.B1(n_7),
.B2(n_8),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_51),
.B1(n_66),
.B2(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_7),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_79),
.B(n_72),
.C(n_85),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_64),
.A3(n_34),
.B1(n_33),
.B2(n_21),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_65),
.C(n_61),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_14),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2x1_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_27),
.Y(n_109)
);

NOR2x1_ASAP7_75t_R g130 ( 
.A(n_109),
.B(n_103),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_117),
.B1(n_90),
.B2(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_0),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_6),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_73),
.B1(n_3),
.B2(n_6),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_122),
.B1(n_128),
.B2(n_116),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_109),
.B(n_114),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_134),
.B1(n_115),
.B2(n_104),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_79),
.B1(n_94),
.B2(n_76),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_76),
.B1(n_75),
.B2(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_1),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_132),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_104),
.B(n_102),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_6),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_7),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_146),
.B1(n_118),
.B2(n_127),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_148),
.B1(n_121),
.B2(n_125),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_145),
.B(n_152),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_98),
.B1(n_101),
.B2(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_108),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_105),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_153),
.C(n_133),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_105),
.C(n_108),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_164),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_123),
.B(n_135),
.C(n_119),
.D(n_121),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_156),
.A2(n_159),
.B(n_163),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_158),
.B1(n_165),
.B2(n_166),
.Y(n_170)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_141),
.B(n_144),
.C(n_148),
.D(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_131),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_121),
.B1(n_134),
.B2(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_149),
.C(n_140),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.C(n_172),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_151),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_146),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_174),
.C(n_172),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_155),
.B1(n_143),
.B2(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_159),
.B1(n_156),
.B2(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_169),
.A2(n_152),
.B1(n_111),
.B2(n_11),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_111),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_173),
.B(n_168),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_181),
.B(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_190),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_184),
.B(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_177),
.C(n_111),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_191),
.B(n_10),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_193),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_189),
.B(n_10),
.C(n_11),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_192),
.B(n_10),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_197),
.B(n_196),
.Y(n_198)
);


endmodule