module fake_netlist_1_9047_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_10), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_4), .B(n_1), .Y(n_15) );
NOR2xp67_ASAP7_75t_L g16 ( .A(n_8), .B(n_4), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AO21x2_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_16), .B(n_15), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_13), .Y(n_21) );
O2A1O1Ixp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_20), .B(n_16), .C(n_18), .Y(n_22) );
O2A1O1Ixp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_2), .B(n_3), .C(n_14), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
OAI22xp5_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_25) );
AOI22xp33_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_7), .B1(n_9), .B2(n_12), .Y(n_26) );
endmodule