module real_aes_16158_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g555 ( .A(n_0), .Y(n_555) );
INVx1_ASAP7_75t_L g678 ( .A(n_1), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g1434 ( .A1(n_1), .A2(n_245), .B1(n_1407), .B2(n_1411), .Y(n_1434) );
INVx1_ASAP7_75t_L g1054 ( .A(n_2), .Y(n_1054) );
INVx1_ASAP7_75t_L g1166 ( .A(n_3), .Y(n_1166) );
AOI221x1_ASAP7_75t_SL g1182 ( .A1(n_3), .A2(n_4), .B1(n_753), .B2(n_838), .C(n_1183), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_4), .A2(n_28), .B1(n_1171), .B2(n_1172), .Y(n_1177) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_5), .A2(n_505), .B(n_646), .C(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g670 ( .A(n_5), .Y(n_670) );
AOI221x1_ASAP7_75t_SL g691 ( .A1(n_6), .A2(n_286), .B1(n_692), .B2(n_694), .C(n_696), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g771 ( .A1(n_6), .A2(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g332 ( .A(n_7), .Y(n_332) );
OAI211xp5_ASAP7_75t_L g440 ( .A1(n_7), .A2(n_441), .B(n_446), .C(n_459), .Y(n_440) );
INVx1_ASAP7_75t_L g1055 ( .A(n_8), .Y(n_1055) );
INVx1_ASAP7_75t_L g1090 ( .A(n_9), .Y(n_1090) );
XNOR2xp5_ASAP7_75t_L g1307 ( .A(n_10), .B(n_1308), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1443 ( .A1(n_10), .A2(n_67), .B1(n_1407), .B2(n_1411), .Y(n_1443) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_11), .Y(n_1275) );
INVx1_ASAP7_75t_L g918 ( .A(n_12), .Y(n_918) );
INVx1_ASAP7_75t_L g1202 ( .A(n_13), .Y(n_1202) );
OAI211xp5_ASAP7_75t_L g1240 ( .A1(n_13), .A2(n_375), .B(n_931), .C(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g797 ( .A(n_14), .Y(n_797) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_14), .A2(n_148), .B1(n_853), .B2(n_858), .Y(n_852) );
INVx1_ASAP7_75t_L g1644 ( .A(n_15), .Y(n_1644) );
AOI22xp33_ASAP7_75t_L g1660 ( .A1(n_15), .A2(n_128), .B1(n_775), .B2(n_1661), .Y(n_1660) );
AOI21xp33_ASAP7_75t_L g1175 ( .A1(n_16), .A2(n_454), .B(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1190 ( .A(n_16), .Y(n_1190) );
INVx1_ASAP7_75t_L g311 ( .A(n_17), .Y(n_311) );
AND2x2_ASAP7_75t_L g429 ( .A(n_17), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g472 ( .A(n_17), .B(n_261), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_17), .B(n_321), .Y(n_550) );
OAI211xp5_ASAP7_75t_SL g1070 ( .A1(n_18), .A2(n_886), .B(n_980), .C(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1082 ( .A(n_18), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g800 ( .A1(n_19), .A2(n_287), .B1(n_801), .B2(n_804), .C(n_805), .Y(n_800) );
INVx1_ASAP7_75t_L g845 ( .A(n_19), .Y(n_845) );
OAI211xp5_ASAP7_75t_L g878 ( .A1(n_20), .A2(n_879), .B(n_880), .C(n_886), .Y(n_878) );
INVx1_ASAP7_75t_L g894 ( .A(n_20), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_21), .A2(n_214), .B1(n_835), .B2(n_1268), .Y(n_1267) );
AOI221xp5_ASAP7_75t_L g1300 ( .A1(n_21), .A2(n_108), .B1(n_457), .B2(n_1301), .C(n_1302), .Y(n_1300) );
INVx1_ASAP7_75t_L g1341 ( .A(n_22), .Y(n_1341) );
INVx1_ASAP7_75t_L g1316 ( .A(n_23), .Y(n_1316) );
INVx1_ASAP7_75t_L g1257 ( .A(n_24), .Y(n_1257) );
INVx2_ASAP7_75t_L g1410 ( .A(n_25), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_25), .B(n_123), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_25), .B(n_1416), .Y(n_1418) );
INVx1_ASAP7_75t_L g1091 ( .A(n_26), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_27), .A2(n_193), .B1(n_870), .B2(n_872), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_27), .A2(n_193), .B1(n_896), .B2(n_897), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_28), .A2(n_211), .B1(n_753), .B2(n_1186), .C(n_1188), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1428 ( .A1(n_29), .A2(n_44), .B1(n_1414), .B2(n_1417), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_30), .A2(n_170), .B1(n_716), .B2(n_719), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_30), .A2(n_265), .B1(n_729), .B2(n_735), .C(n_739), .Y(n_728) );
INVx1_ASAP7_75t_L g975 ( .A(n_31), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g1386 ( .A1(n_32), .A2(n_281), .B1(n_510), .B2(n_960), .Y(n_1386) );
OAI22xp33_ASAP7_75t_L g1394 ( .A1(n_32), .A2(n_281), .B1(n_672), .B2(n_1207), .Y(n_1394) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_33), .A2(n_65), .B1(n_510), .B2(n_511), .Y(n_509) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_33), .A2(n_65), .B1(n_528), .B2(n_531), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_34), .A2(n_48), .B1(n_313), .B2(n_877), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g888 ( .A1(n_34), .A2(n_48), .B1(n_889), .B2(n_890), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g1433 ( .A1(n_35), .A2(n_146), .B1(n_1414), .B2(n_1417), .Y(n_1433) );
OAI211xp5_ASAP7_75t_L g1339 ( .A1(n_36), .A2(n_375), .B(n_636), .C(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1351 ( .A(n_36), .Y(n_1351) );
INVx1_ASAP7_75t_L g1359 ( .A(n_37), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_38), .A2(n_243), .B1(n_398), .B2(n_401), .Y(n_1255) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_38), .A2(n_77), .B1(n_1157), .B2(n_1283), .C(n_1285), .Y(n_1282) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_39), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_40), .A2(n_153), .B1(n_1337), .B2(n_1381), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g1388 ( .A1(n_40), .A2(n_153), .B1(n_877), .B2(n_1389), .Y(n_1388) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_41), .A2(n_215), .B1(n_369), .B2(n_498), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_41), .A2(n_215), .B1(n_313), .B2(n_537), .Y(n_659) );
INVx1_ASAP7_75t_L g1615 ( .A(n_42), .Y(n_1615) );
INVx1_ASAP7_75t_L g1223 ( .A(n_43), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_45), .A2(n_266), .B1(n_413), .B2(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g447 ( .A(n_45), .Y(n_447) );
INVx1_ASAP7_75t_L g917 ( .A(n_46), .Y(n_917) );
INVx1_ASAP7_75t_L g626 ( .A(n_47), .Y(n_626) );
INVx1_ASAP7_75t_L g1201 ( .A(n_49), .Y(n_1201) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_50), .A2(n_112), .B1(n_1407), .B2(n_1421), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_51), .A2(n_117), .B1(n_1407), .B2(n_1493), .Y(n_1492) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_52), .A2(n_194), .B1(n_877), .B2(n_1204), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1239 ( .A1(n_52), .A2(n_194), .B1(n_496), .B2(n_1079), .Y(n_1239) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_53), .A2(n_164), .B1(n_792), .B2(n_793), .C(n_794), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_53), .A2(n_91), .B1(n_398), .B2(n_843), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g1110 ( .A1(n_54), .A2(n_76), .B1(n_956), .B2(n_957), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g1119 ( .A1(n_54), .A2(n_76), .B1(n_496), .B2(n_966), .Y(n_1119) );
AOI22xp33_ASAP7_75t_SL g396 ( .A1(n_55), .A2(n_137), .B1(n_397), .B2(n_401), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_55), .A2(n_266), .B1(n_457), .B2(n_458), .Y(n_464) );
INVx1_ASAP7_75t_L g507 ( .A(n_56), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_57), .A2(n_202), .B1(n_436), .B2(n_709), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_57), .A2(n_120), .B1(n_838), .B2(n_839), .Y(n_837) );
OAI22xp5_ASAP7_75t_SL g1152 ( .A1(n_58), .A2(n_213), .B1(n_816), .B2(n_822), .Y(n_1152) );
INVx1_ASAP7_75t_L g1156 ( .A(n_58), .Y(n_1156) );
INVx1_ASAP7_75t_L g913 ( .A(n_59), .Y(n_913) );
INVx1_ASAP7_75t_L g340 ( .A(n_60), .Y(n_340) );
INVx1_ASAP7_75t_L g348 ( .A(n_60), .Y(n_348) );
INVx1_ASAP7_75t_L g411 ( .A(n_61), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_61), .A2(n_275), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g614 ( .A(n_62), .Y(n_614) );
INVx1_ASAP7_75t_L g1115 ( .A(n_63), .Y(n_1115) );
OAI211xp5_ASAP7_75t_L g1122 ( .A1(n_63), .A2(n_505), .B(n_1123), .C(n_1124), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g1439 ( .A1(n_64), .A2(n_159), .B1(n_1407), .B2(n_1421), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1612 ( .A1(n_64), .A2(n_1613), .B1(n_1662), .B2(n_1663), .Y(n_1612) );
INVxp67_ASAP7_75t_L g1663 ( .A(n_64), .Y(n_1663) );
AOI22xp33_ASAP7_75t_L g1668 ( .A1(n_64), .A2(n_1669), .B1(n_1671), .B2(n_1674), .Y(n_1668) );
INVx1_ASAP7_75t_L g1342 ( .A(n_66), .Y(n_1342) );
OAI211xp5_ASAP7_75t_L g1347 ( .A1(n_66), .A2(n_517), .B(n_1348), .C(n_1350), .Y(n_1347) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_68), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_69), .A2(n_258), .B1(n_1414), .B2(n_1417), .Y(n_1494) );
CKINVDCx5p33_ASAP7_75t_R g1625 ( .A(n_70), .Y(n_1625) );
INVx1_ASAP7_75t_L g1094 ( .A(n_71), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_72), .A2(n_328), .B1(n_329), .B2(n_489), .Y(n_327) );
INVxp67_ASAP7_75t_L g489 ( .A(n_72), .Y(n_489) );
INVx1_ASAP7_75t_L g304 ( .A(n_73), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_74), .Y(n_1008) );
INVx2_ASAP7_75t_L g336 ( .A(n_75), .Y(n_336) );
AOI22xp33_ASAP7_75t_SL g1270 ( .A1(n_77), .A2(n_218), .B1(n_833), .B2(n_1271), .Y(n_1270) );
XOR2x2_ASAP7_75t_L g492 ( .A(n_78), .B(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_79), .A2(n_255), .B1(n_821), .B2(n_823), .Y(n_820) );
INVx1_ASAP7_75t_L g924 ( .A(n_80), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g1646 ( .A1(n_81), .A2(n_295), .B1(n_1171), .B2(n_1301), .Y(n_1646) );
INVx1_ASAP7_75t_L g1652 ( .A(n_81), .Y(n_1652) );
INVx1_ASAP7_75t_L g819 ( .A(n_82), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_83), .Y(n_1030) );
INVx1_ASAP7_75t_L g1057 ( .A(n_84), .Y(n_1057) );
OAI211xp5_ASAP7_75t_L g949 ( .A1(n_85), .A2(n_886), .B(n_950), .C(n_951), .Y(n_949) );
INVx1_ASAP7_75t_L g964 ( .A(n_85), .Y(n_964) );
OAI211xp5_ASAP7_75t_L g1197 ( .A1(n_86), .A2(n_1198), .B(n_1199), .C(n_1200), .Y(n_1197) );
INVx1_ASAP7_75t_L g1242 ( .A(n_86), .Y(n_1242) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_87), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_87), .A2(n_250), .B1(n_471), .B2(n_473), .C(n_478), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_88), .A2(n_128), .B1(n_1172), .B2(n_1633), .Y(n_1632) );
AOI22xp33_ASAP7_75t_L g1653 ( .A1(n_88), .A2(n_230), .B1(n_756), .B2(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g885 ( .A(n_89), .Y(n_885) );
OAI211xp5_ASAP7_75t_L g891 ( .A1(n_89), .A2(n_375), .B(n_646), .C(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g574 ( .A(n_90), .Y(n_574) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_91), .Y(n_808) );
INVx1_ASAP7_75t_L g1265 ( .A(n_92), .Y(n_1265) );
XOR2x2_ASAP7_75t_L g865 ( .A(n_93), .B(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g653 ( .A(n_94), .Y(n_653) );
OAI211xp5_ASAP7_75t_L g660 ( .A1(n_94), .A2(n_661), .B(n_663), .C(n_667), .Y(n_660) );
XOR2x2_ASAP7_75t_L g996 ( .A(n_95), .B(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_95), .A2(n_125), .B1(n_1407), .B2(n_1411), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_96), .Y(n_1004) );
INVx1_ASAP7_75t_L g1063 ( .A(n_97), .Y(n_1063) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_98), .A2(n_221), .B1(n_313), .B2(n_957), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g1034 ( .A1(n_98), .A2(n_221), .B1(n_498), .B2(n_889), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_99), .A2(n_151), .B1(n_1414), .B2(n_1417), .Y(n_1459) );
OAI221xp5_ASAP7_75t_SL g1621 ( .A1(n_100), .A2(n_109), .B1(n_1622), .B2(n_1623), .C(n_1624), .Y(n_1621) );
INVx1_ASAP7_75t_L g1639 ( .A(n_100), .Y(n_1639) );
INVx1_ASAP7_75t_L g631 ( .A(n_101), .Y(n_631) );
INVx1_ASAP7_75t_L g1174 ( .A(n_102), .Y(n_1174) );
INVx1_ASAP7_75t_L g630 ( .A(n_103), .Y(n_630) );
INVx1_ASAP7_75t_L g1059 ( .A(n_104), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_105), .Y(n_362) );
INVx1_ASAP7_75t_L g1061 ( .A(n_106), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_107), .A2(n_127), .B1(n_672), .B2(n_874), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_107), .A2(n_127), .B1(n_655), .B2(n_1121), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_108), .A2(n_152), .B1(n_838), .B2(n_839), .Y(n_1254) );
INVx1_ASAP7_75t_L g1648 ( .A(n_109), .Y(n_1648) );
INVx1_ASAP7_75t_L g1100 ( .A(n_110), .Y(n_1100) );
XNOR2xp5_ASAP7_75t_L g1672 ( .A(n_111), .B(n_1673), .Y(n_1672) );
OA222x2_ASAP7_75t_L g680 ( .A1(n_113), .A2(n_244), .B1(n_265), .B2(n_681), .C1(n_685), .C2(n_689), .Y(n_680) );
INVx1_ASAP7_75t_L g752 ( .A(n_113), .Y(n_752) );
INVx1_ASAP7_75t_L g1366 ( .A(n_114), .Y(n_1366) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_115), .A2(n_1194), .B1(n_1195), .B2(n_1245), .Y(n_1193) );
INVxp67_ASAP7_75t_SL g1245 ( .A(n_115), .Y(n_1245) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_116), .Y(n_306) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_116), .B(n_304), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_118), .A2(n_144), .B1(n_529), .B2(n_874), .Y(n_1075) );
OAI22xp33_ASAP7_75t_L g1083 ( .A1(n_118), .A2(n_144), .B1(n_960), .B2(n_1041), .Y(n_1083) );
INVx1_ASAP7_75t_L g1362 ( .A(n_119), .Y(n_1362) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_120), .A2(n_190), .B1(n_461), .B2(n_462), .C(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g977 ( .A(n_121), .Y(n_977) );
INVx1_ASAP7_75t_L g986 ( .A(n_122), .Y(n_986) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_123), .B(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1416 ( .A(n_123), .Y(n_1416) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_124), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_126), .A2(n_201), .B1(n_1414), .B2(n_1417), .Y(n_1438) );
INVx1_ASAP7_75t_L g569 ( .A(n_129), .Y(n_569) );
INVx1_ASAP7_75t_L g1114 ( .A(n_130), .Y(n_1114) );
INVx1_ASAP7_75t_L g1074 ( .A(n_131), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g1080 ( .A1(n_131), .A2(n_505), .B(n_962), .C(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1363 ( .A(n_132), .Y(n_1363) );
INVx1_ASAP7_75t_L g1050 ( .A(n_133), .Y(n_1050) );
INVx1_ASAP7_75t_L g1085 ( .A(n_134), .Y(n_1085) );
INVx1_ASAP7_75t_L g1360 ( .A(n_135), .Y(n_1360) );
INVx1_ASAP7_75t_L g1619 ( .A(n_136), .Y(n_1619) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_137), .A2(n_452), .B(n_454), .Y(n_451) );
OAI211xp5_ASAP7_75t_L g1382 ( .A1(n_138), .A2(n_501), .B(n_505), .C(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1393 ( .A(n_138), .Y(n_1393) );
INVx2_ASAP7_75t_L g380 ( .A(n_139), .Y(n_380) );
INVx1_ASAP7_75t_L g422 ( .A(n_139), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_139), .B(n_336), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_140), .A2(n_272), .B1(n_510), .B2(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_140), .A2(n_272), .B1(n_672), .B2(n_673), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_141), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_142), .A2(n_290), .B1(n_496), .B2(n_498), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g536 ( .A1(n_142), .A2(n_290), .B1(n_313), .B2(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g1211 ( .A(n_143), .Y(n_1211) );
INVx1_ASAP7_75t_L g1317 ( .A(n_145), .Y(n_1317) );
INVx1_ASAP7_75t_L g1385 ( .A(n_147), .Y(n_1385) );
OAI211xp5_ASAP7_75t_L g1391 ( .A1(n_147), .A2(n_663), .B(n_914), .C(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g798 ( .A(n_148), .Y(n_798) );
INVx1_ASAP7_75t_L g971 ( .A(n_149), .Y(n_971) );
INVx1_ASAP7_75t_L g1101 ( .A(n_150), .Y(n_1101) );
INVx1_ASAP7_75t_L g1287 ( .A(n_152), .Y(n_1287) );
INVxp67_ASAP7_75t_SL g1263 ( .A(n_154), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_154), .A2(n_270), .B1(n_554), .B2(n_1295), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_155), .A2(n_285), .B1(n_436), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_155), .A2(n_268), .B1(n_754), .B2(n_775), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_156), .A2(n_183), .B1(n_528), .B2(n_531), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g1040 ( .A1(n_156), .A2(n_183), .B1(n_511), .B2(n_1041), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_157), .A2(n_276), .B1(n_1414), .B2(n_1417), .Y(n_1413) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_158), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g1458 ( .A1(n_160), .A2(n_161), .B1(n_1407), .B2(n_1411), .Y(n_1458) );
INVx1_ASAP7_75t_L g1312 ( .A(n_162), .Y(n_1312) );
INVx1_ASAP7_75t_L g372 ( .A(n_163), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_163), .A2(n_203), .B1(n_426), .B2(n_434), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_164), .A2(n_208), .B1(n_831), .B2(n_833), .Y(n_830) );
INVx1_ASAP7_75t_L g1219 ( .A(n_165), .Y(n_1219) );
INVx1_ASAP7_75t_L g1134 ( .A(n_166), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_167), .A2(n_242), .B1(n_672), .B2(n_673), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_167), .A2(n_242), .B1(n_896), .B2(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g1031 ( .A(n_168), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g1035 ( .A1(n_168), .A2(n_505), .B(n_1036), .C(n_1038), .Y(n_1035) );
INVx1_ASAP7_75t_L g1322 ( .A(n_169), .Y(n_1322) );
INVx1_ASAP7_75t_L g755 ( .A(n_170), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_171), .A2(n_199), .B1(n_655), .B2(n_1344), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_171), .A2(n_199), .B1(n_531), .B2(n_672), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_172), .A2(n_181), .B1(n_1414), .B2(n_1417), .Y(n_1442) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_173), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_174), .Y(n_707) );
INVx1_ASAP7_75t_L g617 ( .A(n_175), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_176), .Y(n_619) );
INVx1_ASAP7_75t_L g391 ( .A(n_177), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g460 ( .A1(n_177), .A2(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g923 ( .A(n_178), .Y(n_923) );
INVx1_ASAP7_75t_L g1095 ( .A(n_179), .Y(n_1095) );
INVx1_ASAP7_75t_L g1277 ( .A(n_180), .Y(n_1277) );
OAI211xp5_ASAP7_75t_L g1026 ( .A1(n_182), .A2(n_886), .B(n_1027), .C(n_1029), .Y(n_1026) );
INVx1_ASAP7_75t_L g1039 ( .A(n_182), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_184), .A2(n_293), .B1(n_956), .B2(n_957), .Y(n_955) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_184), .A2(n_293), .B1(n_369), .B2(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g1365 ( .A(n_185), .Y(n_1365) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_186), .A2(n_232), .B1(n_537), .B2(n_956), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1078 ( .A1(n_186), .A2(n_232), .B1(n_369), .B2(n_1079), .Y(n_1078) );
BUFx3_ASAP7_75t_L g342 ( .A(n_187), .Y(n_342) );
INVx1_ASAP7_75t_L g1222 ( .A(n_188), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1422 ( .A1(n_189), .A2(n_191), .B1(n_1414), .B2(n_1417), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_190), .A2(n_202), .B1(n_644), .B2(n_835), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g1429 ( .A1(n_192), .A2(n_262), .B1(n_1407), .B2(n_1411), .Y(n_1429) );
CKINVDCx5p33_ASAP7_75t_R g1260 ( .A(n_195), .Y(n_1260) );
INVx1_ASAP7_75t_L g1098 ( .A(n_196), .Y(n_1098) );
INVx1_ASAP7_75t_L g1305 ( .A(n_197), .Y(n_1305) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_198), .Y(n_318) );
INVx1_ASAP7_75t_L g1618 ( .A(n_200), .Y(n_1618) );
INVx1_ASAP7_75t_L g367 ( .A(n_203), .Y(n_367) );
INVx1_ASAP7_75t_L g1324 ( .A(n_204), .Y(n_1324) );
INVx1_ASAP7_75t_L g1371 ( .A(n_205), .Y(n_1371) );
INVx1_ASAP7_75t_L g1319 ( .A(n_206), .Y(n_1319) );
INVx1_ASAP7_75t_L g508 ( .A(n_207), .Y(n_508) );
OAI211xp5_ASAP7_75t_L g514 ( .A1(n_207), .A2(n_515), .B(n_517), .C(n_520), .Y(n_514) );
INVxp67_ASAP7_75t_SL g806 ( .A(n_208), .Y(n_806) );
INVx1_ASAP7_75t_L g981 ( .A(n_209), .Y(n_981) );
INVx1_ASAP7_75t_L g903 ( .A(n_210), .Y(n_903) );
AOI21xp33_ASAP7_75t_L g1167 ( .A1(n_211), .A2(n_1168), .B(n_1169), .Y(n_1167) );
INVx1_ASAP7_75t_L g1097 ( .A(n_212), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g1161 ( .A(n_213), .Y(n_1161) );
INVx1_ASAP7_75t_L g1286 ( .A(n_214), .Y(n_1286) );
XOR2x2_ASAP7_75t_L g784 ( .A(n_216), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g883 ( .A(n_217), .Y(n_883) );
INVx1_ASAP7_75t_L g1303 ( .A(n_218), .Y(n_1303) );
INVx1_ASAP7_75t_L g973 ( .A(n_219), .Y(n_973) );
INVx1_ASAP7_75t_L g611 ( .A(n_220), .Y(n_611) );
INVx1_ASAP7_75t_L g552 ( .A(n_222), .Y(n_552) );
INVx1_ASAP7_75t_L g564 ( .A(n_223), .Y(n_564) );
OAI222xp33_ASAP7_75t_L g1136 ( .A1(n_224), .A2(n_263), .B1(n_279), .B2(n_823), .C1(n_1137), .C2(n_1141), .Y(n_1136) );
XOR2x2_ASAP7_75t_L g604 ( .A(n_225), .B(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_226), .A2(n_296), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g1189 ( .A(n_226), .Y(n_1189) );
OAI211xp5_ASAP7_75t_L g499 ( .A1(n_227), .A2(n_500), .B(n_505), .C(n_506), .Y(n_499) );
INVx1_ASAP7_75t_L g526 ( .A(n_227), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_228), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_229), .Y(n_1001) );
AOI21xp33_ASAP7_75t_L g1645 ( .A1(n_230), .A2(n_454), .B(n_1176), .Y(n_1645) );
INVx1_ASAP7_75t_L g652 ( .A(n_231), .Y(n_652) );
INVx1_ASAP7_75t_L g906 ( .A(n_233), .Y(n_906) );
INVx1_ASAP7_75t_L g1217 ( .A(n_234), .Y(n_1217) );
INVx1_ASAP7_75t_L g1320 ( .A(n_235), .Y(n_1320) );
INVx1_ASAP7_75t_L g559 ( .A(n_236), .Y(n_559) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_237), .Y(n_317) );
INVx1_ASAP7_75t_L g1213 ( .A(n_238), .Y(n_1213) );
INVx1_ASAP7_75t_L g1228 ( .A(n_239), .Y(n_1228) );
OAI22xp33_ASAP7_75t_L g1336 ( .A1(n_240), .A2(n_256), .B1(n_498), .B2(n_1337), .Y(n_1336) );
OAI22xp33_ASAP7_75t_L g1346 ( .A1(n_240), .A2(n_256), .B1(n_313), .B2(n_957), .Y(n_1346) );
OAI211xp5_ASAP7_75t_L g1111 ( .A1(n_241), .A2(n_914), .B(n_1112), .C(n_1113), .Y(n_1111) );
INVx1_ASAP7_75t_L g1125 ( .A(n_241), .Y(n_1125) );
INVx1_ASAP7_75t_L g1304 ( .A(n_243), .Y(n_1304) );
INVx1_ASAP7_75t_L g740 ( .A(n_244), .Y(n_740) );
INVx1_ASAP7_75t_L g357 ( .A(n_246), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_247), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g1629 ( .A1(n_248), .A2(n_257), .B1(n_695), .B2(n_1169), .C(n_1630), .Y(n_1629) );
INVx1_ASAP7_75t_L g1651 ( .A(n_248), .Y(n_1651) );
OAI22xp33_ASAP7_75t_L g1205 ( .A1(n_249), .A2(n_264), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
OAI22xp33_ASAP7_75t_L g1243 ( .A1(n_249), .A2(n_264), .B1(n_897), .B2(n_1121), .Y(n_1243) );
INVx1_ASAP7_75t_L g350 ( .A(n_250), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g1150 ( .A(n_251), .Y(n_1150) );
INVx1_ASAP7_75t_L g1314 ( .A(n_252), .Y(n_1314) );
INVx1_ASAP7_75t_L g571 ( .A(n_253), .Y(n_571) );
INVx1_ASAP7_75t_L g623 ( .A(n_254), .Y(n_623) );
OAI211xp5_ASAP7_75t_L g787 ( .A1(n_255), .A2(n_788), .B(n_790), .C(n_796), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1658 ( .A1(n_257), .A2(n_295), .B1(n_389), .B2(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g985 ( .A(n_259), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g1626 ( .A(n_260), .Y(n_1626) );
BUFx3_ASAP7_75t_L g321 ( .A(n_261), .Y(n_321) );
INVx1_ASAP7_75t_L g430 ( .A(n_261), .Y(n_430) );
XOR2x2_ASAP7_75t_L g1354 ( .A(n_262), .B(n_1355), .Y(n_1354) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_267), .Y(n_706) );
INVx1_ASAP7_75t_L g697 ( .A(n_268), .Y(n_697) );
INVx1_ASAP7_75t_L g915 ( .A(n_269), .Y(n_915) );
INVxp67_ASAP7_75t_SL g1279 ( .A(n_270), .Y(n_1279) );
INVx1_ASAP7_75t_L g1227 ( .A(n_271), .Y(n_1227) );
INVx1_ASAP7_75t_L g1384 ( .A(n_273), .Y(n_1384) );
XOR2x2_ASAP7_75t_L g946 ( .A(n_274), .B(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g395 ( .A(n_275), .Y(n_395) );
INVx1_ASAP7_75t_L g385 ( .A(n_277), .Y(n_385) );
INVx1_ASAP7_75t_L g421 ( .A(n_277), .Y(n_421) );
INVx2_ASAP7_75t_L g488 ( .A(n_277), .Y(n_488) );
INVx1_ASAP7_75t_L g577 ( .A(n_278), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_279), .A2(n_284), .B1(n_434), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1368 ( .A(n_280), .Y(n_1368) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_282), .Y(n_724) );
XNOR2xp5_ASAP7_75t_L g1043 ( .A(n_283), .B(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1151 ( .A(n_284), .Y(n_1151) );
INVx1_ASAP7_75t_L g769 ( .A(n_285), .Y(n_769) );
INVx1_ASAP7_75t_L g768 ( .A(n_286), .Y(n_768) );
INVx1_ASAP7_75t_L g848 ( .A(n_287), .Y(n_848) );
INVx1_ASAP7_75t_L g979 ( .A(n_288), .Y(n_979) );
INVx1_ASAP7_75t_L g1048 ( .A(n_289), .Y(n_1048) );
INVx1_ASAP7_75t_L g1072 ( .A(n_291), .Y(n_1072) );
INVx1_ASAP7_75t_L g953 ( .A(n_292), .Y(n_953) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_292), .A2(n_505), .B(n_962), .C(n_963), .Y(n_961) );
INVx1_ASAP7_75t_L g952 ( .A(n_294), .Y(n_952) );
INVx1_ASAP7_75t_L g1184 ( .A(n_296), .Y(n_1184) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_322), .B(n_1400), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_307), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g1667 ( .A(n_301), .B(n_310), .Y(n_1667) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g1670 ( .A(n_303), .B(n_306), .Y(n_1670) );
INVx1_ASAP7_75t_L g1675 ( .A(n_303), .Y(n_1675) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g1677 ( .A(n_306), .B(n_1675), .Y(n_1677) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g540 ( .A(n_310), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g455 ( .A(n_311), .B(n_321), .Y(n_455) );
AND2x4_ASAP7_75t_L g463 ( .A(n_311), .B(n_320), .Y(n_463) );
INVx1_ASAP7_75t_L g1204 ( .A(n_312), .Y(n_1204) );
AND2x4_ASAP7_75t_SL g1666 ( .A(n_312), .B(n_1667), .Y(n_1666) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_314), .B(n_319), .Y(n_313) );
OR2x6_ASAP7_75t_L g529 ( .A(n_314), .B(n_530), .Y(n_529) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_314), .Y(n_573) );
INVxp67_ASAP7_75t_L g613 ( .A(n_314), .Y(n_613) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g554 ( .A(n_315), .Y(n_554) );
BUFx4f_ASAP7_75t_L g1234 ( .A(n_315), .Y(n_1234) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g432 ( .A(n_317), .Y(n_432) );
INVx2_ASAP7_75t_L g439 ( .A(n_317), .Y(n_439) );
AND2x2_ASAP7_75t_L g444 ( .A(n_317), .B(n_445), .Y(n_444) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_317), .B(n_318), .Y(n_450) );
AND2x2_ASAP7_75t_L g469 ( .A(n_317), .B(n_318), .Y(n_469) );
INVx1_ASAP7_75t_L g482 ( .A(n_317), .Y(n_482) );
INVx1_ASAP7_75t_L g433 ( .A(n_318), .Y(n_433) );
AND2x2_ASAP7_75t_L g438 ( .A(n_318), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g445 ( .A(n_318), .Y(n_445) );
BUFx2_ASAP7_75t_L g476 ( .A(n_318), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_318), .B(n_439), .Y(n_535) );
OR2x2_ASAP7_75t_L g563 ( .A(n_318), .B(n_432), .Y(n_563) );
OR2x6_ASAP7_75t_L g956 ( .A(n_319), .B(n_554), .Y(n_956) );
INVxp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g519 ( .A(n_320), .Y(n_519) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g522 ( .A(n_321), .Y(n_522) );
AND2x4_ASAP7_75t_L g525 ( .A(n_321), .B(n_481), .Y(n_525) );
XNOR2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_779), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
XNOR2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_490), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_377), .B(n_386), .C(n_423), .Y(n_329) );
NAND4xp25_ASAP7_75t_L g330 ( .A(n_331), .B(n_349), .C(n_366), .D(n_375), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_343), .B2(n_344), .Y(n_331) );
INVx2_ASAP7_75t_L g498 ( .A(n_333), .Y(n_498) );
INVx1_ASAP7_75t_L g890 ( .A(n_333), .Y(n_890) );
INVx1_ASAP7_75t_L g966 ( .A(n_333), .Y(n_966) );
INVx2_ASAP7_75t_L g1079 ( .A(n_333), .Y(n_1079) );
INVxp67_ASAP7_75t_L g1381 ( .A(n_333), .Y(n_1381) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
OR2x4_ASAP7_75t_L g374 ( .A(n_334), .B(n_370), .Y(n_374) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x6_ASAP7_75t_L g345 ( .A(n_335), .B(n_346), .Y(n_345) );
OR2x4_ASAP7_75t_L g369 ( .A(n_335), .B(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g376 ( .A(n_335), .B(n_364), .Y(n_376) );
NAND3x1_ASAP7_75t_L g419 ( .A(n_335), .B(n_420), .C(n_422), .Y(n_419) );
AND2x4_ASAP7_75t_L g733 ( .A(n_335), .B(n_734), .Y(n_733) );
NAND2x1p5_ASAP7_75t_L g766 ( .A(n_335), .B(n_422), .Y(n_766) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
NAND2xp33_ASAP7_75t_SL g406 ( .A(n_336), .B(n_380), .Y(n_406) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_337), .Y(n_592) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_337), .Y(n_644) );
INVx1_ASAP7_75t_L g1005 ( .A(n_337), .Y(n_1005) );
INVx2_ASAP7_75t_L g1378 ( .A(n_337), .Y(n_1378) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g390 ( .A(n_338), .Y(n_390) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_338), .Y(n_598) );
BUFx8_ASAP7_75t_L g772 ( .A(n_338), .Y(n_772) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
AND2x4_ASAP7_75t_L g399 ( .A(n_341), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_342), .B(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_342), .Y(n_356) );
AND2x4_ASAP7_75t_L g364 ( .A(n_342), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g960 ( .A(n_344), .Y(n_960) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g512 ( .A(n_345), .Y(n_512) );
INVx1_ASAP7_75t_L g656 ( .A(n_345), .Y(n_656) );
BUFx3_ASAP7_75t_L g897 ( .A(n_345), .Y(n_897) );
INVx1_ASAP7_75t_L g595 ( .A(n_346), .Y(n_595) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_346), .Y(n_1323) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
INVx1_ASAP7_75t_L g361 ( .A(n_348), .Y(n_361) );
INVx2_ASAP7_75t_L g365 ( .A(n_348), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_357), .B2(n_358), .C1(n_362), .C2(n_363), .Y(n_349) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_351), .A2(n_359), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_351), .A2(n_358), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g893 ( .A(n_352), .Y(n_893) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
AND2x4_ASAP7_75t_L g359 ( .A(n_353), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g651 ( .A(n_353), .B(n_355), .Y(n_651) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND3x4_ASAP7_75t_L g829 ( .A(n_354), .B(n_380), .C(n_487), .Y(n_829) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_356), .B(n_361), .Y(n_504) );
INVx2_ASAP7_75t_L g732 ( .A(n_356), .Y(n_732) );
AND2x4_ASAP7_75t_L g754 ( .A(n_356), .B(n_738), .Y(n_754) );
AOI211xp5_ASAP7_75t_SL g465 ( .A1(n_357), .A2(n_466), .B(n_470), .C(n_483), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_358), .A2(n_883), .B1(n_893), .B2(n_894), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_358), .A2(n_893), .B1(n_1201), .B2(n_1242), .Y(n_1241) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_359), .A2(n_651), .B1(n_652), .B2(n_653), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_359), .A2(n_651), .B1(n_952), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g1038 ( .A1(n_359), .A2(n_651), .B1(n_1030), .B2(n_1039), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_359), .A2(n_651), .B1(n_1072), .B2(n_1082), .Y(n_1081) );
AOI22xp33_ASAP7_75t_SL g1124 ( .A1(n_359), .A2(n_651), .B1(n_1114), .B2(n_1125), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_359), .A2(n_651), .B1(n_1384), .B2(n_1385), .Y(n_1383) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_362), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g416 ( .A(n_363), .Y(n_416) );
BUFx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
BUFx3_ASAP7_75t_L g743 ( .A(n_364), .Y(n_743) );
BUFx2_ASAP7_75t_L g756 ( .A(n_364), .Y(n_756) );
BUFx2_ASAP7_75t_L g833 ( .A(n_364), .Y(n_833) );
BUFx2_ASAP7_75t_L g864 ( .A(n_364), .Y(n_864) );
INVx1_ASAP7_75t_L g738 ( .A(n_365), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_372), .B2(n_373), .Y(n_366) );
INVx2_ASAP7_75t_L g889 ( .A(n_368), .Y(n_889) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g497 ( .A(n_369), .Y(n_497) );
INVx1_ASAP7_75t_L g1338 ( .A(n_369), .Y(n_1338) );
BUFx3_ASAP7_75t_L g587 ( .A(n_370), .Y(n_587) );
BUFx3_ASAP7_75t_L g764 ( .A(n_370), .Y(n_764) );
INVx2_ASAP7_75t_L g855 ( .A(n_370), .Y(n_855) );
BUFx4f_ASAP7_75t_L g930 ( .A(n_370), .Y(n_930) );
INVx1_ASAP7_75t_L g400 ( .A(n_371), .Y(n_400) );
INVx2_ASAP7_75t_L g1041 ( .A(n_373), .Y(n_1041) );
INVx1_ASAP7_75t_L g1121 ( .A(n_373), .Y(n_1121) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g510 ( .A(n_374), .Y(n_510) );
BUFx2_ASAP7_75t_L g896 ( .A(n_374), .Y(n_896) );
BUFx2_ASAP7_75t_L g1344 ( .A(n_374), .Y(n_1344) );
CKINVDCx8_ASAP7_75t_R g375 ( .A(n_376), .Y(n_375) );
CKINVDCx8_ASAP7_75t_R g505 ( .A(n_376), .Y(n_505) );
OAI31xp33_ASAP7_75t_L g494 ( .A1(n_377), .A2(n_495), .A3(n_499), .B(n_509), .Y(n_494) );
CKINVDCx14_ASAP7_75t_R g898 ( .A(n_377), .Y(n_898) );
OAI31xp33_ASAP7_75t_L g1033 ( .A1(n_377), .A2(n_1034), .A3(n_1035), .B(n_1040), .Y(n_1033) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .Y(n_377) );
AND2x2_ASAP7_75t_L g657 ( .A(n_378), .B(n_381), .Y(n_657) );
AND2x2_ASAP7_75t_L g967 ( .A(n_378), .B(n_381), .Y(n_967) );
AND2x2_ASAP7_75t_SL g1244 ( .A(n_378), .B(n_381), .Y(n_1244) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g734 ( .A(n_380), .Y(n_734) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g405 ( .A(n_383), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g581 ( .A(n_383), .Y(n_581) );
OR2x2_ASAP7_75t_L g818 ( .A(n_383), .B(n_760), .Y(n_818) );
AND2x2_ASAP7_75t_SL g983 ( .A(n_383), .B(n_455), .Y(n_983) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g542 ( .A(n_384), .Y(n_542) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_403), .B1(n_407), .B2(n_417), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_391), .B1(n_392), .B2(n_395), .C(n_396), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_388), .A2(n_913), .B1(n_923), .B2(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g408 ( .A(n_390), .Y(n_408) );
INVx3_ASAP7_75t_L g641 ( .A(n_390), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_392), .A2(n_617), .B1(n_630), .B2(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_392), .A2(n_591), .B1(n_768), .B2(n_769), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_392), .A2(n_1008), .B1(n_1009), .B2(n_1010), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1377 ( .A1(n_392), .A2(n_1363), .B1(n_1371), .B2(n_1378), .Y(n_1377) );
CKINVDCx8_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g410 ( .A(n_393), .Y(n_410) );
INVx3_ASAP7_75t_L g935 ( .A(n_393), .Y(n_935) );
INVx1_ASAP7_75t_L g992 ( .A(n_393), .Y(n_992) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g817 ( .A(n_394), .Y(n_817) );
BUFx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g414 ( .A(n_398), .Y(n_414) );
INVx2_ASAP7_75t_SL g832 ( .A(n_398), .Y(n_832) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx8_ASAP7_75t_L g742 ( .A(n_399), .Y(n_742) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_399), .Y(n_748) );
NAND2x1p5_ASAP7_75t_L g824 ( .A(n_399), .B(n_733), .Y(n_824) );
BUFx3_ASAP7_75t_L g1656 ( .A(n_399), .Y(n_1656) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g843 ( .A(n_402), .Y(n_843) );
INVx2_ASAP7_75t_L g1661 ( .A(n_402), .Y(n_1661) );
OAI33xp33_ASAP7_75t_L g1209 ( .A1(n_403), .A2(n_1210), .A3(n_1216), .B1(n_1220), .B2(n_1224), .B3(n_1226), .Y(n_1209) );
OAI33xp33_ASAP7_75t_L g1310 ( .A1(n_403), .A2(n_1011), .A3(n_1311), .B1(n_1315), .B2(n_1318), .B3(n_1321), .Y(n_1310) );
BUFx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx4f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx8_ASAP7_75t_L g583 ( .A(n_405), .Y(n_583) );
BUFx4f_ASAP7_75t_L g926 ( .A(n_405), .Y(n_926) );
BUFx2_ASAP7_75t_L g988 ( .A(n_405), .Y(n_988) );
BUFx2_ASAP7_75t_L g773 ( .A(n_406), .Y(n_773) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_410), .B2(n_411), .C(n_412), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_408), .A2(n_975), .B1(n_985), .B2(n_992), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_408), .A2(n_410), .B1(n_1054), .B2(n_1055), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_408), .A2(n_1057), .B1(n_1058), .B2(n_1059), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_408), .A2(n_992), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_409), .A2(n_448), .B(n_460), .C(n_464), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_410), .A2(n_915), .B1(n_924), .B2(n_937), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_410), .A2(n_977), .B1(n_986), .B2(n_994), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_410), .A2(n_994), .B1(n_1097), .B2(n_1098), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_410), .A2(n_1362), .B1(n_1368), .B2(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI33xp33_ASAP7_75t_L g925 ( .A1(n_417), .A2(n_926), .A3(n_927), .B1(n_934), .B2(n_936), .B3(n_939), .Y(n_925) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_418), .Y(n_1011) );
AOI221xp5_ASAP7_75t_L g1181 ( .A1(n_418), .A2(n_863), .B1(n_1182), .B2(n_1185), .C(n_1191), .Y(n_1181) );
NAND3xp33_ASAP7_75t_L g1657 ( .A(n_418), .B(n_1658), .C(n_1660), .Y(n_1657) );
INVx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g601 ( .A(n_419), .Y(n_601) );
OAI33xp33_ASAP7_75t_L g632 ( .A1(n_419), .A2(n_583), .A3(n_633), .B1(n_639), .B2(n_642), .B3(n_645), .Y(n_632) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g684 ( .A(n_421), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_421), .B(n_429), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_465), .B(n_484), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_440), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_427), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g722 ( .A(n_428), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
AND2x2_ASAP7_75t_L g435 ( .A(n_429), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g442 ( .A(n_429), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_SL g467 ( .A(n_429), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g726 ( .A(n_429), .B(n_443), .Y(n_726) );
AND2x4_ASAP7_75t_L g789 ( .A(n_429), .B(n_458), .Y(n_789) );
BUFx2_ASAP7_75t_L g1290 ( .A(n_429), .Y(n_1290) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_430), .Y(n_530) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_431), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_431), .B(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g710 ( .A(n_431), .Y(n_710) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_432), .Y(n_1163) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g1647 ( .A1(n_435), .A2(n_466), .B1(n_1615), .B2(n_1648), .Y(n_1647) );
AND2x4_ASAP7_75t_L g686 ( .A(n_436), .B(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_438), .Y(n_458) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_438), .Y(n_1172) );
BUFx3_ASAP7_75t_L g1301 ( .A(n_438), .Y(n_1301) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_442), .Y(n_799) );
BUFx6f_ASAP7_75t_L g1176 ( .A(n_443), .Y(n_1176) );
INVx2_ASAP7_75t_L g1293 ( .A(n_443), .Y(n_1293) );
INVx1_ASAP7_75t_L g1631 ( .A(n_443), .Y(n_1631) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g453 ( .A(n_444), .Y(n_453) );
AND2x4_ASAP7_75t_L g538 ( .A(n_444), .B(n_530), .Y(n_538) );
BUFx3_ASAP7_75t_L g1168 ( .A(n_444), .Y(n_1168) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_451), .C(n_456), .Y(n_446) );
INVx1_ASAP7_75t_L g1028 ( .A(n_448), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_448), .A2(n_976), .B1(n_1054), .B2(n_1057), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_448), .A2(n_976), .B1(n_1050), .B2(n_1063), .Y(n_1067) );
BUFx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g625 ( .A(n_449), .Y(n_625) );
OR2x2_ASAP7_75t_L g689 ( .A(n_449), .B(n_688), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_449), .B(n_1298), .Y(n_1297) );
BUFx2_ASAP7_75t_SL g1331 ( .A(n_449), .Y(n_1331) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_450), .Y(n_516) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g461 ( .A(n_453), .Y(n_461) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g579 ( .A(n_455), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g794 ( .A(n_455), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_455), .B(n_580), .Y(n_921) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_455), .A2(n_516), .B1(n_562), .B2(n_1303), .C(n_1304), .Y(n_1302) );
BUFx6f_ASAP7_75t_L g1157 ( .A(n_457), .Y(n_1157) );
A2O1A1Ixp33_ASAP7_75t_L g1296 ( .A1(n_457), .A2(n_1265), .B(n_1297), .C(n_1299), .Y(n_1296) );
INVx1_ASAP7_75t_L g1284 ( .A(n_458), .Y(n_1284) );
INVx2_ASAP7_75t_L g693 ( .A(n_461), .Y(n_693) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g1169 ( .A(n_463), .Y(n_1169) );
OAI221xp5_ASAP7_75t_L g1285 ( .A1(n_463), .A2(n_911), .B1(n_1022), .B2(n_1286), .C(n_1287), .Y(n_1285) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g803 ( .A(n_467), .Y(n_803) );
AND2x6_ASAP7_75t_L g483 ( .A(n_468), .B(n_472), .Y(n_483) );
AND2x2_ASAP7_75t_L g518 ( .A(n_468), .B(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_468), .Y(n_695) );
BUFx3_ASAP7_75t_L g792 ( .A(n_468), .Y(n_792) );
INVx1_ASAP7_75t_L g811 ( .A(n_468), .Y(n_811) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g666 ( .A(n_469), .Y(n_666) );
OR2x2_ASAP7_75t_L g683 ( .A(n_471), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g477 ( .A(n_472), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_472), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_472), .B(n_488), .Y(n_714) );
HB1xp67_ASAP7_75t_L g1164 ( .A(n_472), .Y(n_1164) );
BUFx2_ASAP7_75t_L g804 ( .A(n_473), .Y(n_804) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g1638 ( .A(n_475), .Y(n_1638) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g521 ( .A(n_476), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g718 ( .A(n_476), .Y(n_718) );
AND2x4_ASAP7_75t_L g882 ( .A(n_476), .B(n_522), .Y(n_882) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_476), .Y(n_1160) );
INVx1_ASAP7_75t_L g1299 ( .A(n_477), .Y(n_1299) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g719 ( .A(n_480), .B(n_542), .Y(n_719) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_SL g790 ( .A1(n_483), .A2(n_791), .B(n_795), .Y(n_790) );
INVx1_ASAP7_75t_L g812 ( .A(n_484), .Y(n_812) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_485), .Y(n_1180) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI31xp33_ASAP7_75t_L g1281 ( .A1(n_486), .A2(n_1282), .A3(n_1288), .B(n_1300), .Y(n_1281) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g549 ( .A(n_488), .Y(n_549) );
OAI22x1_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_675), .B1(n_676), .B2(n_778), .Y(n_490) );
INVx1_ASAP7_75t_L g778 ( .A(n_491), .Y(n_778) );
XNOR2x1_ASAP7_75t_L g491 ( .A(n_492), .B(n_604), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_513), .C(n_543), .Y(n_493) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI211xp5_ASAP7_75t_L g770 ( .A1(n_501), .A2(n_706), .B(n_771), .C(n_774), .Y(n_770) );
OAI22xp33_ASAP7_75t_L g989 ( .A1(n_501), .A2(n_971), .B1(n_979), .B2(n_990), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_501), .A2(n_930), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g589 ( .A(n_503), .Y(n_589) );
OR2x2_ASAP7_75t_L g822 ( .A(n_503), .B(n_818), .Y(n_822) );
BUFx6f_ASAP7_75t_L g1062 ( .A(n_503), .Y(n_1062) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g638 ( .A(n_504), .Y(n_638) );
BUFx3_ASAP7_75t_L g933 ( .A(n_504), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_507), .A2(n_521), .B1(n_523), .B2(n_526), .Y(n_520) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI31xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_527), .A3(n_536), .B(n_539), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_515), .A2(n_559), .B1(n_560), .B2(n_564), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_515), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_515), .A2(n_976), .B1(n_1094), .B2(n_1097), .Y(n_1104) );
INVx1_ASAP7_75t_L g1349 ( .A(n_515), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g1364 ( .A1(n_515), .A2(n_618), .B1(n_1365), .B2(n_1366), .Y(n_1364) );
BUFx4f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx4f_ASAP7_75t_L g570 ( .A(n_516), .Y(n_570) );
INVx4_ASAP7_75t_L g662 ( .A(n_516), .Y(n_662) );
OR2x6_ASAP7_75t_L g711 ( .A(n_516), .B(n_712), .Y(n_711) );
BUFx4f_ASAP7_75t_L g914 ( .A(n_516), .Y(n_914) );
BUFx6f_ASAP7_75t_L g950 ( .A(n_516), .Y(n_950) );
BUFx4f_ASAP7_75t_L g1198 ( .A(n_516), .Y(n_1198) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g886 ( .A(n_518), .Y(n_886) );
INVx1_ASAP7_75t_L g1199 ( .A(n_518), .Y(n_1199) );
AND2x2_ASAP7_75t_L g664 ( .A(n_519), .B(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_521), .A2(n_652), .B1(n_668), .B2(n_670), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_521), .A2(n_523), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_521), .A2(n_1072), .B1(n_1073), .B2(n_1074), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_521), .A2(n_1073), .B1(n_1114), .B2(n_1115), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_521), .A2(n_668), .B1(n_1341), .B2(n_1351), .Y(n_1350) );
OR2x2_ASAP7_75t_L g533 ( .A(n_522), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g1073 ( .A(n_524), .Y(n_1073) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g669 ( .A(n_525), .Y(n_669) );
BUFx3_ASAP7_75t_L g884 ( .A(n_525), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_525), .A2(n_882), .B1(n_952), .B2(n_953), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_525), .A2(n_882), .B1(n_1384), .B2(n_1393), .Y(n_1392) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_529), .Y(n_672) );
INVx1_ASAP7_75t_L g871 ( .A(n_529), .Y(n_871) );
HB1xp67_ASAP7_75t_L g1206 ( .A(n_529), .Y(n_1206) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g673 ( .A(n_532), .Y(n_673) );
INVx1_ASAP7_75t_L g1207 ( .A(n_532), .Y(n_1207) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g875 ( .A(n_533), .Y(n_875) );
INVx8_ASAP7_75t_L g557 ( .A(n_534), .Y(n_557) );
BUFx2_ASAP7_75t_L g807 ( .A(n_534), .Y(n_807) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx3_ASAP7_75t_SL g877 ( .A(n_538), .Y(n_877) );
CKINVDCx16_ASAP7_75t_R g957 ( .A(n_538), .Y(n_957) );
OAI31xp33_ASAP7_75t_L g948 ( .A1(n_539), .A2(n_949), .A3(n_954), .B(n_955), .Y(n_948) );
BUFx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
BUFx3_ASAP7_75t_L g674 ( .A(n_540), .Y(n_674) );
INVx1_ASAP7_75t_L g867 ( .A(n_540), .Y(n_867) );
OAI31xp33_ASAP7_75t_L g1069 ( .A1(n_540), .A2(n_1070), .A3(n_1075), .B(n_1076), .Y(n_1069) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_540), .Y(n_1117) );
OAI31xp33_ASAP7_75t_L g1196 ( .A1(n_540), .A2(n_1197), .A3(n_1203), .B(n_1205), .Y(n_1196) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g723 ( .A(n_542), .Y(n_723) );
INVxp67_ASAP7_75t_L g825 ( .A(n_542), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_582), .Y(n_543) );
OAI33xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_551), .A3(n_558), .B1(n_565), .B2(n_572), .B3(n_578), .Y(n_544) );
OAI33xp33_ASAP7_75t_L g1064 ( .A1(n_545), .A2(n_982), .A3(n_1065), .B1(n_1066), .B2(n_1067), .B3(n_1068), .Y(n_1064) );
OAI33xp33_ASAP7_75t_L g1357 ( .A1(n_545), .A2(n_578), .A3(n_1358), .B1(n_1361), .B2(n_1364), .B3(n_1367), .Y(n_1357) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g609 ( .A(n_548), .Y(n_609) );
INVx1_ASAP7_75t_L g703 ( .A(n_548), .Y(n_703) );
INVx2_ASAP7_75t_L g901 ( .A(n_548), .Y(n_901) );
INVx2_ASAP7_75t_L g1105 ( .A(n_548), .Y(n_1105) );
AND2x4_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g777 ( .A(n_549), .Y(n_777) );
OR2x6_ASAP7_75t_L g841 ( .A(n_549), .B(n_766), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B1(n_555), .B2(n_556), .Y(n_551) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_552), .A2(n_569), .B1(n_585), .B2(n_588), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_553), .A2(n_1314), .B1(n_1324), .B2(n_1333), .Y(n_1332) );
BUFx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_SL g629 ( .A(n_554), .Y(n_629) );
BUFx3_ASAP7_75t_L g698 ( .A(n_554), .Y(n_698) );
BUFx6f_ASAP7_75t_L g972 ( .A(n_554), .Y(n_972) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_555), .A2(n_571), .B1(n_585), .B2(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_556), .A2(n_628), .B1(n_1006), .B2(n_1010), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_556), .A2(n_1368), .B1(n_1369), .B2(n_1371), .Y(n_1367) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_557), .Y(n_576) );
INVx2_ASAP7_75t_SL g615 ( .A(n_557), .Y(n_615) );
INVx2_ASAP7_75t_L g700 ( .A(n_557), .Y(n_700) );
INVx4_ASAP7_75t_L g909 ( .A(n_557), .Y(n_909) );
INVx2_ASAP7_75t_L g1295 ( .A(n_557), .Y(n_1295) );
INVx1_ASAP7_75t_L g1327 ( .A(n_557), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_559), .A2(n_574), .B1(n_591), .B2(n_593), .Y(n_590) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g568 ( .A(n_563), .Y(n_568) );
INVx1_ASAP7_75t_L g622 ( .A(n_563), .Y(n_622) );
INVx2_ASAP7_75t_L g912 ( .A(n_563), .Y(n_912) );
BUFx2_ASAP7_75t_L g976 ( .A(n_563), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_564), .A2(n_577), .B1(n_593), .B2(n_597), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_566), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_566), .A2(n_980), .B1(n_1091), .B2(n_1101), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g1328 ( .A1(n_566), .A2(n_624), .B1(n_1312), .B2(n_1322), .Y(n_1328) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_566), .A2(n_624), .B1(n_1362), .B2(n_1363), .Y(n_1361) );
INVx4_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g618 ( .A(n_567), .Y(n_618) );
INVx2_ASAP7_75t_L g1330 ( .A(n_567), .Y(n_1330) );
INVx4_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_570), .A2(n_621), .B1(n_706), .B2(n_707), .C(n_708), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_577), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_573), .A2(n_575), .B1(n_985), .B2(n_986), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_573), .A2(n_807), .B1(n_1055), .B2(n_1059), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_573), .A2(n_807), .B1(n_1095), .B2(n_1098), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_573), .A2(n_1316), .B1(n_1319), .B2(n_1327), .Y(n_1326) );
OAI22xp33_ASAP7_75t_L g1358 ( .A1(n_573), .A2(n_699), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_575), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g1017 ( .A1(n_575), .A2(n_628), .B1(n_1001), .B2(n_1013), .Y(n_1017) );
INVx5_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx6_ASAP7_75t_L g1333 ( .A(n_576), .Y(n_1333) );
OAI33xp33_ASAP7_75t_L g607 ( .A1(n_578), .A2(n_608), .A3(n_610), .B1(n_616), .B2(n_620), .B3(n_627), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_578), .A2(n_705), .B(n_711), .Y(n_704) );
OAI33xp33_ASAP7_75t_L g1016 ( .A1(n_578), .A2(n_608), .A3(n_1017), .B1(n_1018), .B2(n_1019), .B3(n_1023), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g1334 ( .A(n_579), .Y(n_1334) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI33xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .A3(n_590), .B1(n_596), .B2(n_599), .B3(n_602), .Y(n_582) );
OAI33xp33_ASAP7_75t_L g999 ( .A1(n_583), .A2(n_1000), .A3(n_1003), .B1(n_1007), .B2(n_1011), .B3(n_1012), .Y(n_999) );
OAI33xp33_ASAP7_75t_L g1372 ( .A1(n_583), .A2(n_841), .A3(n_1373), .B1(n_1374), .B2(n_1376), .B3(n_1377), .Y(n_1372) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_585), .A2(n_1013), .B1(n_1014), .B2(n_1015), .Y(n_1012) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g635 ( .A(n_587), .Y(n_635) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g603 ( .A(n_589), .Y(n_603) );
INVx1_ASAP7_75t_L g646 ( .A(n_589), .Y(n_646) );
INVx2_ASAP7_75t_L g763 ( .A(n_589), .Y(n_763) );
INVx1_ASAP7_75t_L g1037 ( .A(n_589), .Y(n_1037) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_593), .A2(n_619), .B1(n_631), .B2(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_593), .A2(n_1004), .B1(n_1005), .B2(n_1006), .Y(n_1003) );
OAI22xp33_ASAP7_75t_SL g1311 ( .A1(n_593), .A2(n_1312), .B1(n_1313), .B2(n_1314), .Y(n_1311) );
OAI221xp5_ASAP7_75t_L g1650 ( .A1(n_593), .A2(n_1378), .B1(n_1651), .B2(n_1652), .C(n_1653), .Y(n_1650) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx8_ASAP7_75t_L g838 ( .A(n_597), .Y(n_838) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_597), .Y(n_1009) );
INVx5_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx3_ASAP7_75t_L g750 ( .A(n_598), .Y(n_750) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_598), .Y(n_938) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_598), .Y(n_1269) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_601), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_603), .A2(n_1049), .B1(n_1174), .B2(n_1184), .Y(n_1183) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_647), .C(n_658), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_632), .Y(n_606) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_614), .B2(n_615), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_611), .A2(n_623), .B1(n_634), .B2(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_614), .A2(n_626), .B1(n_634), .B2(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B1(n_624), .B2(n_626), .Y(n_620) );
OAI22xp5_ASAP7_75t_SL g1018 ( .A1(n_621), .A2(n_950), .B1(n_1004), .B2(n_1008), .Y(n_1018) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_624), .A2(n_911), .B1(n_917), .B2(n_918), .Y(n_916) );
OAI211xp5_ASAP7_75t_L g1643 ( .A1(n_624), .A2(n_1644), .B(n_1645), .C(n_1646), .Y(n_1643) );
INVx5_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_628), .A2(n_806), .B1(n_807), .B2(n_808), .C(n_809), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_628), .A2(n_909), .B1(n_1048), .B2(n_1061), .Y(n_1065) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_634), .A2(n_931), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVxp67_ASAP7_75t_SL g1014 ( .A(n_637), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g1102 ( .A(n_637), .Y(n_1102) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g1052 ( .A(n_638), .Y(n_1052) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_641), .B(n_857), .Y(n_1144) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g1375 ( .A(n_644), .Y(n_1375) );
OAI31xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .A3(n_654), .B(n_657), .Y(n_647) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI31xp33_ASAP7_75t_L g1335 ( .A1(n_657), .A2(n_1336), .A3(n_1339), .B(n_1343), .Y(n_1335) );
OAI31xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .A3(n_671), .B(n_674), .Y(n_658) );
OAI22xp5_ASAP7_75t_SL g974 ( .A1(n_661), .A2(n_975), .B1(n_976), .B2(n_977), .Y(n_974) );
NAND2xp5_ASAP7_75t_SL g1158 ( .A(n_661), .B(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g879 ( .A(n_662), .Y(n_879) );
INVx2_ASAP7_75t_L g980 ( .A(n_662), .Y(n_980) );
INVx2_ASAP7_75t_L g1022 ( .A(n_662), .Y(n_1022) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g1112 ( .A(n_664), .Y(n_1112) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx2_ASAP7_75t_L g1641 ( .A(n_666), .Y(n_1641) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI31xp33_ASAP7_75t_L g1024 ( .A1(n_674), .A2(n_1025), .A3(n_1026), .B(n_1032), .Y(n_1024) );
OAI31xp33_ASAP7_75t_L g1345 ( .A1(n_674), .A2(n_1346), .A3(n_1347), .B(n_1352), .Y(n_1345) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
XNOR2x1_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND4xp75_ASAP7_75t_L g679 ( .A(n_680), .B(n_690), .C(n_720), .D(n_727), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g815 ( .A(n_683), .B(n_816), .Y(n_815) );
AND2x4_ASAP7_75t_L g847 ( .A(n_684), .B(n_733), .Y(n_847) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI211x1_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_702), .B(n_704), .C(n_715), .Y(n_690) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g793 ( .A(n_693), .Y(n_793) );
BUFx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_695), .A2(n_1257), .B1(n_1277), .B2(n_1292), .C(n_1294), .Y(n_1291) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_699), .B2(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g905 ( .A(n_698), .Y(n_905) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g762 ( .A1(n_701), .A2(n_707), .B1(n_763), .B2(n_764), .C(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI33xp33_ASAP7_75t_L g1229 ( .A1(n_703), .A2(n_919), .A3(n_1230), .B1(n_1235), .B2(n_1236), .B3(n_1237), .Y(n_1229) );
OAI33xp33_ASAP7_75t_L g1325 ( .A1(n_703), .A2(n_1326), .A3(n_1328), .B1(n_1329), .B2(n_1332), .B3(n_1334), .Y(n_1325) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g1171 ( .A(n_710), .Y(n_1171) );
INVx2_ASAP7_75t_L g1633 ( .A(n_710), .Y(n_1633) );
INVx2_ASAP7_75t_SL g1636 ( .A(n_710), .Y(n_1636) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2x2_ASAP7_75t_L g716 ( .A(n_713), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g821 ( .A(n_719), .B(n_822), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_724), .B2(n_725), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_721), .A2(n_724), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx3_ASAP7_75t_L g1139 ( .A(n_722), .Y(n_1139) );
AND2x4_ASAP7_75t_L g725 ( .A(n_723), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g1145 ( .A(n_725), .Y(n_1145) );
OAI31xp67_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_746), .A3(n_761), .B(n_776), .Y(n_727) );
INVx4_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x6_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
AND2x2_ASAP7_75t_L g846 ( .A(n_731), .B(n_847), .Y(n_846) );
NAND2x1_ASAP7_75t_L g1149 ( .A(n_731), .B(n_847), .Y(n_1149) );
AND2x4_ASAP7_75t_SL g1274 ( .A(n_731), .B(n_847), .Y(n_1274) );
INVx3_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g736 ( .A(n_733), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g745 ( .A(n_733), .Y(n_745) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g851 ( .A(n_737), .Y(n_851) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_743), .C(n_744), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_L g775 ( .A(n_742), .Y(n_775) );
INVx2_ASAP7_75t_L g1262 ( .A(n_742), .Y(n_1262) );
INVx8_ASAP7_75t_L g1271 ( .A(n_742), .Y(n_1271) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_751), .B(n_757), .Y(n_746) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_755), .B2(n_756), .Y(n_751) );
BUFx3_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx5_ASAP7_75t_L g836 ( .A(n_754), .Y(n_836) );
BUFx3_ASAP7_75t_L g839 ( .A(n_754), .Y(n_839) );
BUFx12f_ASAP7_75t_L g1659 ( .A(n_754), .Y(n_1659) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI21xp5_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_767), .B(n_770), .Y(n_761) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_763), .Y(n_962) );
OAI22xp33_ASAP7_75t_L g1099 ( .A1(n_764), .A2(n_1100), .B1(n_1101), .B2(n_1102), .Y(n_1099) );
OAI22xp33_ASAP7_75t_L g1318 ( .A1(n_764), .A2(n_931), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x4_ASAP7_75t_L g859 ( .A(n_772), .B(n_860), .Y(n_859) );
INVx2_ASAP7_75t_SL g994 ( .A(n_772), .Y(n_994) );
INVx2_ASAP7_75t_SL g1187 ( .A(n_772), .Y(n_1187) );
INVx3_ASAP7_75t_L g1221 ( .A(n_772), .Y(n_1221) );
AOI31xp33_ASAP7_75t_L g1627 ( .A1(n_776), .A2(n_1628), .A3(n_1643), .B(n_1647), .Y(n_1627) );
BUFx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_1129), .B1(n_1130), .B2(n_1399), .Y(n_779) );
INVx1_ASAP7_75t_L g1399 ( .A(n_780), .Y(n_1399) );
OA22x2_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_943), .B1(n_944), .B2(n_1128), .Y(n_780) );
INVx1_ASAP7_75t_L g1128 ( .A(n_781), .Y(n_1128) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
XNOR2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_865), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_813), .C(n_826), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_800), .B(n_812), .Y(n_786) );
INVx2_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g1179 ( .A(n_802), .Y(n_1179) );
INVx4_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AOI21xp33_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_819), .B(n_820), .Y(n_813) );
INVx8_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g1264 ( .A(n_816), .Y(n_1264) );
OR2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_817), .Y(n_1058) );
INVx1_ASAP7_75t_L g857 ( .A(n_818), .Y(n_857) );
INVx1_ASAP7_75t_L g860 ( .A(n_818), .Y(n_860) );
INVx2_ASAP7_75t_L g1259 ( .A(n_822), .Y(n_1259) );
INVx5_ASAP7_75t_L g1280 ( .A(n_823), .Y(n_1280) );
INVx3_ASAP7_75t_L g1616 ( .A(n_823), .Y(n_1616) );
OR2x6_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_852), .C(n_861), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_828), .B(n_844), .Y(n_827) );
AOI33xp33_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .A3(n_834), .B1(n_837), .B2(n_840), .B3(n_842), .Y(n_828) );
BUFx3_ASAP7_75t_L g1191 ( .A(n_829), .Y(n_1191) );
NAND3xp33_ASAP7_75t_L g1253 ( .A(n_829), .B(n_1254), .C(n_1255), .Y(n_1253) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g1218 ( .A(n_838), .Y(n_1218) );
INVx1_ASAP7_75t_L g1313 ( .A(n_838), .Y(n_1313) );
NAND3xp33_ASAP7_75t_L g1266 ( .A(n_840), .B(n_1267), .C(n_1270), .Y(n_1266) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI33xp33_ASAP7_75t_L g987 ( .A1(n_841), .A2(n_988), .A3(n_989), .B1(n_991), .B2(n_993), .B3(n_995), .Y(n_987) );
OAI33xp33_ASAP7_75t_L g1046 ( .A1(n_841), .A2(n_988), .A3(n_1047), .B1(n_1053), .B2(n_1056), .B3(n_1060), .Y(n_1046) );
OAI33xp33_ASAP7_75t_L g1088 ( .A1(n_841), .A2(n_988), .A3(n_1089), .B1(n_1093), .B2(n_1096), .B3(n_1099), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_848), .B2(n_849), .Y(n_844) );
AND2x4_ASAP7_75t_L g849 ( .A(n_847), .B(n_850), .Y(n_849) );
AND2x4_ASAP7_75t_L g863 ( .A(n_847), .B(n_864), .Y(n_863) );
AND2x4_ASAP7_75t_SL g1276 ( .A(n_847), .B(n_850), .Y(n_1276) );
AOI221xp5_ASAP7_75t_L g1147 ( .A1(n_849), .A2(n_1148), .B1(n_1150), .B2(n_1151), .C(n_1152), .Y(n_1147) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
OR2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_856), .Y(n_853) );
INVx2_ASAP7_75t_SL g941 ( .A(n_854), .Y(n_941) );
OR2x6_ASAP7_75t_L g1140 ( .A(n_854), .B(n_856), .Y(n_1140) );
INVx2_ASAP7_75t_SL g854 ( .A(n_855), .Y(n_854) );
INVx3_ASAP7_75t_L g990 ( .A(n_855), .Y(n_990) );
INVxp67_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_859), .B(n_1257), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1261 ( .A(n_860), .B(n_1262), .Y(n_1261) );
INVx2_ASAP7_75t_SL g861 ( .A(n_862), .Y(n_861) );
OAI211xp5_ASAP7_75t_SL g1649 ( .A1(n_862), .A2(n_926), .B(n_1650), .C(n_1657), .Y(n_1649) );
INVx3_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_863), .A2(n_1274), .B1(n_1275), .B2(n_1276), .C(n_1277), .Y(n_1273) );
OAI221xp5_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B1(n_887), .B2(n_898), .C(n_899), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_876), .C(n_878), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
OAI211xp5_ASAP7_75t_L g1165 ( .A1(n_879), .A2(n_1166), .B(n_1167), .C(n_1170), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_881), .A2(n_884), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
BUFx3_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NOR3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_891), .C(n_895), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_925), .Y(n_899) );
OAI33xp33_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_902), .A3(n_910), .B1(n_916), .B2(n_919), .B3(n_922), .Y(n_900) );
OAI33xp33_ASAP7_75t_L g969 ( .A1(n_901), .A2(n_970), .A3(n_974), .B1(n_978), .B2(n_982), .B3(n_984), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B1(n_906), .B2(n_907), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_903), .A2(n_917), .B1(n_928), .B2(n_931), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_904), .A2(n_907), .B1(n_923), .B2(n_924), .Y(n_922) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_906), .A2(n_918), .B1(n_940), .B2(n_942), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_907), .A2(n_1211), .B1(n_1227), .B2(n_1231), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1237 ( .A1(n_907), .A2(n_1219), .B1(n_1223), .B2(n_1231), .Y(n_1237) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_909), .A2(n_971), .B1(n_972), .B2(n_973), .Y(n_970) );
OAI22xp33_ASAP7_75t_L g1106 ( .A1(n_909), .A2(n_972), .B1(n_1090), .B2(n_1100), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_913), .B1(n_914), .B2(n_915), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_911), .A2(n_914), .B1(n_1217), .B2(n_1222), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_911), .A2(n_914), .B1(n_1213), .B2(n_1228), .Y(n_1236) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_912), .Y(n_1021) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g1226 ( .A1(n_931), .A2(n_1212), .B1(n_1227), .B2(n_1228), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_931), .A2(n_990), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g1123 ( .A(n_932), .Y(n_1123) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
BUFx6f_ASAP7_75t_L g942 ( .A(n_933), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_933), .A2(n_973), .B1(n_981), .B2(n_990), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_935), .A2(n_1217), .B1(n_1218), .B2(n_1219), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_935), .A2(n_1221), .B1(n_1222), .B2(n_1223), .Y(n_1220) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g1212 ( .A(n_941), .Y(n_1212) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_1042), .B1(n_1126), .B2(n_1127), .Y(n_944) );
INVx1_ASAP7_75t_L g1126 ( .A(n_945), .Y(n_1126) );
XNOR2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_996), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_958), .C(n_968), .Y(n_947) );
INVx1_ASAP7_75t_L g1390 ( .A(n_956), .Y(n_1390) );
OAI31xp33_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_961), .A3(n_965), .B(n_967), .Y(n_958) );
OAI31xp33_ASAP7_75t_L g1077 ( .A1(n_967), .A2(n_1078), .A3(n_1080), .B(n_1083), .Y(n_1077) );
OAI31xp33_ASAP7_75t_SL g1118 ( .A1(n_967), .A2(n_1119), .A3(n_1120), .B(n_1122), .Y(n_1118) );
OAI31xp33_ASAP7_75t_L g1379 ( .A1(n_967), .A2(n_1380), .A3(n_1382), .B(n_1386), .Y(n_1379) );
NOR2xp33_ASAP7_75t_SL g968 ( .A(n_969), .B(n_987), .Y(n_968) );
OAI33xp33_ASAP7_75t_L g1103 ( .A1(n_982), .A2(n_1104), .A3(n_1105), .B1(n_1106), .B2(n_1107), .B3(n_1108), .Y(n_1103) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
BUFx4f_ASAP7_75t_SL g1049 ( .A(n_990), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_990), .A2(n_1061), .B1(n_1062), .B2(n_1063), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1373 ( .A1(n_990), .A2(n_1037), .B1(n_1359), .B2(n_1365), .Y(n_1373) );
OAI22xp33_ASAP7_75t_L g1376 ( .A1(n_990), .A2(n_1051), .B1(n_1360), .B2(n_1366), .Y(n_1376) );
NAND3xp33_ASAP7_75t_L g997 ( .A(n_998), .B(n_1024), .C(n_1033), .Y(n_997) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1016), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_1002), .A2(n_1015), .B1(n_1020), .B2(n_1022), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1321 ( .A1(n_1009), .A2(n_1322), .B1(n_1323), .B2(n_1324), .Y(n_1321) );
INVx4_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
OAI211xp5_ASAP7_75t_L g1173 ( .A1(n_1022), .A2(n_1174), .B(n_1175), .C(n_1177), .Y(n_1173) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1042), .Y(n_1127) );
XOR2xp5_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1084), .Y(n_1042) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1069), .C(n_1077), .Y(n_1044) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1064), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_1049), .A2(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1089) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1052), .Y(n_1092) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1062), .Y(n_1215) );
XNOR2xp5_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1086), .Y(n_1084) );
AND3x1_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1109), .C(n_1118), .Y(n_1086) );
NOR2xp33_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1103), .Y(n_1087) );
OAI31xp33_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1111), .A3(n_1116), .B(n_1117), .Y(n_1109) );
OAI31xp33_ASAP7_75t_SL g1387 ( .A1(n_1117), .A2(n_1388), .A3(n_1391), .B(n_1394), .Y(n_1387) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_1131), .A2(n_1247), .B1(n_1397), .B2(n_1398), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1397 ( .A(n_1132), .Y(n_1397) );
AO22x2_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1192), .B1(n_1193), .B2(n_1246), .Y(n_1132) );
INVx1_ASAP7_75t_SL g1246 ( .A(n_1133), .Y(n_1246) );
XNOR2x1_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
NOR2x1_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1146), .Y(n_1135) );
INVxp67_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_1138), .A2(n_1142), .B1(n_1618), .B2(n_1619), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1140), .Y(n_1138) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
NAND2x1_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1145), .Y(n_1142) );
INVx2_ASAP7_75t_SL g1143 ( .A(n_1144), .Y(n_1143) );
NAND3xp33_ASAP7_75t_SL g1146 ( .A(n_1147), .B(n_1153), .C(n_1181), .Y(n_1146) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_1150), .A2(n_1160), .B1(n_1161), .B2(n_1162), .Y(n_1159) );
OAI21xp5_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1178), .B(n_1180), .Y(n_1153) );
NAND3xp33_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1165), .C(n_1173), .Y(n_1154) );
A2O1A1Ixp33_ASAP7_75t_L g1155 ( .A1(n_1156), .A2(n_1157), .B(n_1158), .C(n_1164), .Y(n_1155) );
AOI22xp5_ASAP7_75t_L g1298 ( .A1(n_1160), .A2(n_1162), .B1(n_1260), .B2(n_1275), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1637 ( .A1(n_1162), .A2(n_1626), .B1(n_1638), .B2(n_1639), .C(n_1640), .Y(n_1637) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1164), .Y(n_1642) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1208), .C(n_1238), .Y(n_1195) );
NOR2xp33_ASAP7_75t_SL g1208 ( .A(n_1209), .B(n_1229), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1212), .B1(n_1213), .B2(n_1214), .Y(n_1210) );
INVx2_ASAP7_75t_SL g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx2_ASAP7_75t_SL g1232 ( .A(n_1233), .Y(n_1232) );
INVx3_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
BUFx6f_ASAP7_75t_L g1370 ( .A(n_1234), .Y(n_1370) );
OAI31xp33_ASAP7_75t_L g1238 ( .A1(n_1239), .A2(n_1240), .A3(n_1243), .B(n_1244), .Y(n_1238) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1247), .Y(n_1398) );
AOI22xp5_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1249), .B1(n_1306), .B2(n_1396), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
XNOR2x1_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1305), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1272), .Y(n_1251) );
NAND4xp25_ASAP7_75t_SL g1252 ( .A(n_1253), .B(n_1256), .C(n_1258), .D(n_1266), .Y(n_1252) );
AOI222xp33_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1260), .B1(n_1261), .B2(n_1263), .C1(n_1264), .C2(n_1265), .Y(n_1258) );
AOI22xp5_ASAP7_75t_L g1624 ( .A1(n_1259), .A2(n_1264), .B1(n_1625), .B2(n_1626), .Y(n_1624) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
NAND3xp33_ASAP7_75t_SL g1272 ( .A(n_1273), .B(n_1278), .C(n_1281), .Y(n_1272) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1274), .Y(n_1622) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1276), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1280), .Y(n_1278) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
OAI21xp5_ASAP7_75t_SL g1288 ( .A1(n_1289), .A2(n_1291), .B(n_1296), .Y(n_1288) );
INVxp67_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1306), .Y(n_1396) );
OA22x2_ASAP7_75t_L g1306 ( .A1(n_1307), .A2(n_1353), .B1(n_1354), .B2(n_1395), .Y(n_1306) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1307), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1335), .C(n_1345), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1325), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_1317), .A2(n_1320), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx2_ASAP7_75t_SL g1353 ( .A(n_1354), .Y(n_1353) );
NAND3xp33_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1379), .C(n_1387), .Y(n_1355) );
NOR2xp33_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1372), .Y(n_1356) );
INVx3_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
OAI221xp5_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1608), .B1(n_1610), .B2(n_1664), .C(n_1668), .Y(n_1400) );
AND4x1_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1563), .C(n_1581), .D(n_1597), .Y(n_1401) );
OAI33xp33_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1495), .A3(n_1513), .B1(n_1519), .B2(n_1531), .B3(n_1542), .Y(n_1402) );
OAI211xp5_ASAP7_75t_SL g1403 ( .A1(n_1404), .A2(n_1423), .B(n_1444), .C(n_1476), .Y(n_1403) );
INVx2_ASAP7_75t_L g1497 ( .A(n_1404), .Y(n_1497) );
AOI331xp33_ASAP7_75t_L g1520 ( .A1(n_1404), .A2(n_1425), .A3(n_1490), .B1(n_1518), .B2(n_1521), .B3(n_1523), .C1(n_1524), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1555 ( .A(n_1404), .B(n_1446), .Y(n_1555) );
NOR2xp33_ASAP7_75t_L g1598 ( .A(n_1404), .B(n_1426), .Y(n_1598) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1419), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1405), .B(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1405), .Y(n_1468) );
INVx2_ASAP7_75t_SL g1489 ( .A(n_1405), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1405), .B(n_1426), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1405), .B(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1413), .Y(n_1405) );
AND2x6_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1409), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1408), .B(n_1412), .Y(n_1411) );
AND2x4_ASAP7_75t_L g1414 ( .A(n_1408), .B(n_1415), .Y(n_1414) );
AND2x6_ASAP7_75t_L g1417 ( .A(n_1408), .B(n_1418), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1408), .B(n_1412), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1408), .B(n_1412), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1410), .B(n_1416), .Y(n_1415) );
OAI21xp5_ASAP7_75t_L g1674 ( .A1(n_1412), .A2(n_1675), .B(n_1676), .Y(n_1674) );
CKINVDCx5p33_ASAP7_75t_R g1461 ( .A(n_1419), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1419), .B(n_1468), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1485 ( .A(n_1419), .B(n_1427), .Y(n_1485) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1419), .B(n_1526), .Y(n_1525) );
AOI22xp5_ASAP7_75t_L g1532 ( .A1(n_1419), .A2(n_1511), .B1(n_1533), .B2(n_1536), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g1572 ( .A1(n_1419), .A2(n_1505), .B1(n_1573), .B2(n_1579), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1419), .B(n_1456), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1419), .B(n_1457), .Y(n_1607) );
AND2x4_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1422), .Y(n_1419) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1430), .Y(n_1424) );
O2A1O1Ixp33_ASAP7_75t_SL g1469 ( .A1(n_1425), .A2(n_1470), .B(n_1471), .C(n_1473), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1425), .B(n_1584), .Y(n_1583) );
CKINVDCx14_ASAP7_75t_R g1425 ( .A(n_1426), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1502 ( .A(n_1426), .B(n_1431), .Y(n_1502) );
NOR2xp33_ASAP7_75t_L g1504 ( .A(n_1426), .B(n_1505), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1426), .B(n_1465), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1426), .B(n_1497), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1534 ( .A(n_1426), .B(n_1535), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1426), .B(n_1430), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1426), .B(n_1489), .Y(n_1569) );
INVx3_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
CKINVDCx5p33_ASAP7_75t_R g1450 ( .A(n_1427), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1427), .B(n_1472), .Y(n_1471) );
OR2x2_ASAP7_75t_L g1499 ( .A(n_1427), .B(n_1500), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1427), .B(n_1432), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_1427), .B(n_1505), .Y(n_1529) );
AND2x4_ASAP7_75t_SL g1427 ( .A(n_1428), .B(n_1429), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1435), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1431), .B(n_1441), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1431), .B(n_1464), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1431), .B(n_1484), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1431), .B(n_1478), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1431), .B(n_1465), .Y(n_1546) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1431), .B(n_1436), .Y(n_1551) );
OR2x2_ASAP7_75t_L g1562 ( .A(n_1431), .B(n_1447), .Y(n_1562) );
OR2x2_ASAP7_75t_L g1591 ( .A(n_1431), .B(n_1509), .Y(n_1591) );
INVx2_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1432), .B(n_1447), .Y(n_1446) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1432), .B(n_1441), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1432), .B(n_1478), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1432), .B(n_1448), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1500 ( .A(n_1432), .B(n_1437), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1432), .B(n_1518), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1432), .B(n_1479), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1432), .B(n_1437), .Y(n_1578) );
NOR2xp33_ASAP7_75t_L g1593 ( .A(n_1432), .B(n_1594), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1434), .Y(n_1432) );
NOR2xp33_ASAP7_75t_L g1594 ( .A(n_1435), .B(n_1472), .Y(n_1594) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
OR2x2_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1440), .Y(n_1436) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1437), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1437), .B(n_1441), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1439), .Y(n_1437) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1441), .B(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1441), .Y(n_1479) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1441), .Y(n_1484) );
NAND2x1_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1443), .Y(n_1441) );
AOI221xp5_ASAP7_75t_L g1444 ( .A1(n_1445), .A2(n_1453), .B1(n_1462), .B2(n_1466), .C(n_1469), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1449), .Y(n_1445) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1446), .Y(n_1584) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1447), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1448), .B(n_1479), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1451), .Y(n_1449) );
OR2x2_ASAP7_75t_L g1515 ( .A(n_1450), .B(n_1452), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1450), .B(n_1478), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1450), .B(n_1487), .Y(n_1536) );
OR2x2_ASAP7_75t_L g1548 ( .A(n_1450), .B(n_1467), .Y(n_1548) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1450), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1450), .B(n_1528), .Y(n_1588) );
AOI22xp5_ASAP7_75t_L g1539 ( .A1(n_1451), .A2(n_1461), .B1(n_1506), .B2(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1453), .B(n_1462), .Y(n_1530) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1460), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1456), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1456), .B(n_1474), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1456), .B(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1457), .Y(n_1490) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1457), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1457), .B(n_1461), .Y(n_1523) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_1457), .B(n_1554), .Y(n_1553) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1457), .B(n_1569), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1459), .Y(n_1457) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1461), .B(n_1489), .Y(n_1488) );
OAI32xp33_ASAP7_75t_L g1501 ( .A1(n_1461), .A2(n_1470), .A3(n_1478), .B1(n_1502), .B2(n_1503), .Y(n_1501) );
HB1xp67_ASAP7_75t_SL g1514 ( .A(n_1461), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1461), .B(n_1508), .Y(n_1574) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1602 ( .A(n_1464), .B(n_1502), .Y(n_1602) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1465), .B(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1467), .Y(n_1596) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1468), .Y(n_1474) );
AOI31xp33_ASAP7_75t_L g1585 ( .A1(n_1468), .A2(n_1545), .A3(n_1586), .B(n_1587), .Y(n_1585) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1470), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1521 ( .A(n_1470), .B(n_1522), .Y(n_1521) );
OAI221xp5_ASAP7_75t_L g1531 ( .A1(n_1473), .A2(n_1490), .B1(n_1532), .B2(n_1537), .C(n_1539), .Y(n_1531) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1475), .Y(n_1473) );
OAI221xp5_ASAP7_75t_SL g1495 ( .A1(n_1474), .A2(n_1496), .B1(n_1508), .B2(n_1509), .C(n_1510), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1474), .B(n_1506), .Y(n_1580) );
AOI221xp5_ASAP7_75t_L g1476 ( .A1(n_1477), .A2(n_1480), .B1(n_1481), .B2(n_1490), .C(n_1491), .Y(n_1476) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1477), .Y(n_1604) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1478), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_1478), .B(n_1507), .Y(n_1576) );
OAI22xp33_ASAP7_75t_L g1481 ( .A1(n_1482), .A2(n_1485), .B1(n_1486), .B2(n_1488), .Y(n_1481) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVxp33_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1488), .Y(n_1535) );
INVx2_ASAP7_75t_L g1505 ( .A(n_1489), .Y(n_1505) );
O2A1O1Ixp33_ASAP7_75t_L g1513 ( .A1(n_1489), .A2(n_1514), .B(n_1515), .C(n_1516), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1489), .B(n_1506), .Y(n_1565) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1490), .Y(n_1564) );
AOI221xp5_ASAP7_75t_L g1597 ( .A1(n_1490), .A2(n_1584), .B1(n_1598), .B2(n_1599), .C(n_1603), .Y(n_1597) );
INVx3_ASAP7_75t_L g1556 ( .A(n_1491), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1494), .Y(n_1491) );
HB1xp67_ASAP7_75t_L g1609 ( .A(n_1493), .Y(n_1609) );
AOI211xp5_ASAP7_75t_L g1496 ( .A1(n_1497), .A2(n_1498), .B(n_1501), .C(n_1506), .Y(n_1496) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1505), .B(n_1523), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1512), .Y(n_1510) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1512), .Y(n_1567) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1530), .Y(n_1519) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1523), .Y(n_1559) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_1523), .A2(n_1574), .B1(n_1575), .B2(n_1577), .Y(n_1573) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
INVxp33_ASAP7_75t_SL g1605 ( .A(n_1526), .Y(n_1605) );
NOR2xp33_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1529), .Y(n_1526) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1536), .Y(n_1586) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
NAND3xp33_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1549), .C(n_1557), .Y(n_1542) );
INVxp67_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
AOI21xp33_ASAP7_75t_L g1544 ( .A1(n_1545), .A2(n_1547), .B(n_1548), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
NOR2xp33_ASAP7_75t_L g1570 ( .A(n_1546), .B(n_1571), .Y(n_1570) );
AOI211xp5_ASAP7_75t_L g1549 ( .A1(n_1550), .A2(n_1552), .B(n_1555), .C(n_1556), .Y(n_1549) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
NOR2xp33_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1560), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1562), .Y(n_1560) );
INVx2_ASAP7_75t_L g1571 ( .A(n_1562), .Y(n_1571) );
AOI211xp5_ASAP7_75t_L g1563 ( .A1(n_1564), .A2(n_1565), .B(n_1566), .C(n_1572), .Y(n_1563) );
AOI21xp33_ASAP7_75t_L g1566 ( .A1(n_1567), .A2(n_1568), .B(n_1570), .Y(n_1566) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVxp33_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
O2A1O1Ixp33_ASAP7_75t_L g1581 ( .A1(n_1582), .A2(n_1585), .B(n_1589), .C(n_1590), .Y(n_1581) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
AOI21xp5_ASAP7_75t_L g1590 ( .A1(n_1591), .A2(n_1592), .B(n_1595), .Y(n_1590) );
INVxp33_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVxp67_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
AOI21xp33_ASAP7_75t_L g1603 ( .A1(n_1604), .A2(n_1605), .B(n_1606), .Y(n_1603) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVx4_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
HB1xp67_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1613), .Y(n_1662) );
NAND3xp33_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1617), .C(n_1620), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
NOR3xp33_ASAP7_75t_SL g1620 ( .A(n_1621), .B(n_1627), .C(n_1649), .Y(n_1620) );
NAND2xp5_ASAP7_75t_L g1635 ( .A(n_1625), .B(n_1636), .Y(n_1635) );
AOI21xp5_ASAP7_75t_L g1628 ( .A1(n_1629), .A2(n_1632), .B(n_1634), .Y(n_1628) );
INVx2_ASAP7_75t_SL g1630 ( .A(n_1631), .Y(n_1630) );
AOI21xp5_ASAP7_75t_L g1634 ( .A1(n_1635), .A2(n_1637), .B(n_1642), .Y(n_1634) );
INVx2_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
HB1xp67_ASAP7_75t_L g1673 ( .A(n_1662), .Y(n_1673) );
INVx2_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
BUFx3_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
HB1xp67_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVxp33_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
endmodule