module fake_jpeg_5649_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx12_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_0),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_13),
.B(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_1),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_18),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_6),
.B1(n_9),
.B2(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_13),
.C(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_17),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_25),
.B1(n_22),
.B2(n_20),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_9),
.B1(n_16),
.B2(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_23),
.B1(n_24),
.B2(n_16),
.Y(n_28)
);

AOI322xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_29),
.A3(n_12),
.B1(n_27),
.B2(n_14),
.C1(n_7),
.C2(n_5),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_29),
.B(n_7),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_7),
.C2(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_2),
.C(n_3),
.Y(n_33)
);


endmodule