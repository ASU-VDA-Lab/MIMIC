module fake_jpeg_31836_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_0),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_48),
.B1(n_44),
.B2(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_47),
.B1(n_40),
.B2(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_68),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_44),
.B(n_48),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_41),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_39),
.C(n_49),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_1),
.C(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_4),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_6),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_44),
.B(n_20),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_14),
.B(n_15),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_80),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_21),
.C(n_37),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_4),
.B(n_5),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_26),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_95),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_23),
.B1(n_9),
.B2(n_10),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_98),
.B1(n_99),
.B2(n_29),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_8),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_100),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_19),
.B(n_24),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_30),
.C(n_33),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_27),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_106),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_109),
.C(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_114),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_104),
.B1(n_110),
.B2(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_113),
.B1(n_107),
.B2(n_111),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_116),
.C(n_101),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_35),
.C(n_36),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_119),
.Y(n_120)
);


endmodule