module fake_jpeg_11018_n_45 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_19),
.B1(n_20),
.B2(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_25),
.Y(n_26)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.C(n_8),
.Y(n_33)
);

BUFx24_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_30),
.Y(n_32)
);

AOI22x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_33),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_9),
.C(n_15),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_16),
.C(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_1),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_11),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_6),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_37),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_35),
.B1(n_4),
.B2(n_5),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_1),
.B(n_4),
.Y(n_45)
);


endmodule