module fake_jpeg_24822_n_166 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_2),
.C(n_3),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_3),
.Y(n_45)
);

OR2x4_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_48),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_29),
.B1(n_25),
.B2(n_15),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_22),
.B(n_19),
.C(n_30),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_50),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_29),
.B1(n_25),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_65),
.B1(n_19),
.B2(n_20),
.Y(n_87)
);

CKINVDCx11_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_52),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_58),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_21),
.B(n_24),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_21),
.B1(n_28),
.B2(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_19),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_7),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_23),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_91),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_64),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_87),
.B1(n_30),
.B2(n_20),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_19),
.B1(n_30),
.B2(n_20),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_49),
.B1(n_46),
.B2(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_55),
.C(n_60),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_16),
.C(n_10),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_96),
.B(n_85),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_54),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_109),
.Y(n_115)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_106),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_104),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_60),
.B(n_30),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_113),
.C(n_94),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_16),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_60),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_80),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_61),
.B1(n_20),
.B2(n_16),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_111),
.B1(n_83),
.B2(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_117),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_126),
.B1(n_109),
.B2(n_107),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_79),
.C(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_119),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_90),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_91),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_127),
.C(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_128),
.B(n_95),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_91),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_132),
.C(n_133),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_105),
.C(n_96),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_128),
.B1(n_108),
.B2(n_116),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_110),
.C(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_145),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_138),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_115),
.B1(n_111),
.B2(n_108),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_134),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_98),
.B(n_86),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_132),
.C(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

OAI321xp33_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_101),
.A3(n_84),
.B1(n_121),
.B2(n_73),
.C(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_153),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_148),
.C(n_144),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_129),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_157),
.C(n_158),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_146),
.B1(n_145),
.B2(n_143),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_148),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_74),
.C(n_11),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_150),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_157),
.A3(n_159),
.B1(n_103),
.B2(n_74),
.C1(n_13),
.C2(n_12),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.C(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_8),
.Y(n_166)
);


endmodule