module fake_jpeg_11486_n_387 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_58),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_50),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_59),
.Y(n_100)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_26),
.B(n_13),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_71),
.Y(n_115)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_13),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_33),
.B(n_11),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_10),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_10),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_82),
.Y(n_84)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_98),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_42),
.B1(n_21),
.B2(n_27),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_86),
.A2(n_97),
.B1(n_108),
.B2(n_118),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_53),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_21),
.B1(n_34),
.B2(n_24),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_94),
.B(n_121),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_42),
.B1(n_21),
.B2(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_52),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_18),
.B1(n_41),
.B2(n_38),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_119),
.B1(n_83),
.B2(n_5),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_42),
.B1(n_44),
.B2(n_23),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_44),
.B1(n_40),
.B2(n_41),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_113),
.B1(n_83),
.B2(n_2),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_44),
.B1(n_40),
.B2(n_36),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_17),
.B1(n_36),
.B2(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_129),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_17),
.B1(n_35),
.B2(n_31),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_47),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_61),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_123),
.B1(n_4),
.B2(n_5),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_60),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_71),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_0),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_72),
.B1(n_69),
.B2(n_81),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_133),
.A2(n_135),
.B1(n_142),
.B2(n_94),
.Y(n_184)
);

AOI222xp33_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_63),
.B1(n_54),
.B2(n_66),
.C1(n_65),
.C2(n_68),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_134),
.A2(n_109),
.B(n_101),
.C(n_90),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_72),
.B1(n_69),
.B2(n_62),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_138),
.Y(n_178)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_49),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_147),
.Y(n_199)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_1),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_149),
.C(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_10),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_3),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_83),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_155),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_3),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_4),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_167),
.Y(n_179)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_162),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_173),
.B1(n_143),
.B2(n_152),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_165),
.B1(n_95),
.B2(n_105),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_107),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_164),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_6),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_169),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_6),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_131),
.B(n_9),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_172),
.Y(n_210)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_9),
.B1(n_121),
.B2(n_117),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_114),
.B(n_122),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_92),
.C(n_125),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_176),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_107),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_181),
.B(n_188),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_191),
.B1(n_203),
.B2(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_130),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_198),
.B1(n_209),
.B2(n_91),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_130),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_212),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_100),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_215),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_131),
.B1(n_124),
.B2(n_126),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_148),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_194),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_197),
.B(n_200),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_149),
.A2(n_126),
.B1(n_124),
.B2(n_105),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_142),
.A2(n_92),
.B1(n_91),
.B2(n_109),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_206),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_168),
.B1(n_170),
.B2(n_134),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_112),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_112),
.Y(n_215)
);

CKINVDCx11_ASAP7_75t_R g216 ( 
.A(n_161),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_161),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_228),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_231),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_181),
.A2(n_159),
.B(n_170),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_154),
.B1(n_145),
.B2(n_141),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_225),
.B1(n_230),
.B2(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_166),
.B1(n_162),
.B2(n_172),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_90),
.B(n_157),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_237),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_214),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_139),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_187),
.C(n_200),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_234),
.C(n_180),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_151),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

AO22x1_ASAP7_75t_SL g237 ( 
.A1(n_184),
.A2(n_153),
.B1(n_146),
.B2(n_136),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_175),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_246),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_179),
.B1(n_191),
.B2(n_192),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_213),
.B1(n_183),
.B2(n_202),
.Y(n_268)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_177),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_196),
.A2(n_179),
.B1(n_199),
.B2(n_190),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_192),
.A2(n_104),
.B(n_125),
.C(n_102),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_247),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_125),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_102),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_189),
.B(n_99),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_189),
.B(n_9),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_218),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_270),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_249),
.A2(n_194),
.B1(n_193),
.B2(n_195),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_257),
.A2(n_227),
.B(n_229),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_259),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_220),
.A2(n_198),
.A3(n_180),
.B1(n_177),
.B2(n_208),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_195),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_226),
.B(n_214),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_274),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_218),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_183),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_216),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_222),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_202),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_227),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_202),
.B1(n_182),
.B2(n_204),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_280),
.B1(n_257),
.B2(n_236),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_247),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_251),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_223),
.A2(n_182),
.B1(n_204),
.B2(n_227),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_275),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_234),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_294),
.C(n_253),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_292),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_290),
.B1(n_301),
.B2(n_255),
.Y(n_310)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_252),
.A2(n_219),
.B1(n_241),
.B2(n_237),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_233),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_296),
.A2(n_303),
.B(n_261),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_246),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_248),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_228),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_304),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_255),
.B1(n_280),
.B2(n_276),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_260),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_302),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_249),
.B(n_245),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_233),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_306),
.C(n_315),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_307),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_310),
.A2(n_311),
.B1(n_314),
.B2(n_286),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_268),
.B1(n_261),
.B2(n_249),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_279),
.B1(n_277),
.B2(n_256),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_265),
.C(n_253),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_284),
.A2(n_278),
.B1(n_262),
.B2(n_256),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_320),
.B1(n_286),
.B2(n_285),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_284),
.A2(n_262),
.B1(n_259),
.B2(n_260),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_294),
.C(n_282),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_281),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_258),
.Y(n_322)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_322),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_300),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_283),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_332),
.B1(n_340),
.B2(n_225),
.Y(n_354)
);

A2O1A1O1Ixp25_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_309),
.B(n_317),
.C(n_289),
.D(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_326),
.B(n_330),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_327),
.A2(n_331),
.B1(n_312),
.B2(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_329),
.A2(n_333),
.B1(n_335),
.B2(n_339),
.Y(n_353)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_293),
.B(n_320),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_297),
.C(n_303),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_337),
.A2(n_338),
.B(n_287),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_322),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_310),
.A2(n_288),
.B1(n_296),
.B2(n_287),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_305),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_321),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_346),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_345),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_306),
.C(n_315),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_307),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_348),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_332),
.B(n_314),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_318),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_340),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_328),
.A2(n_329),
.B1(n_318),
.B2(n_336),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_350),
.B(n_352),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_351),
.A2(n_336),
.B(n_313),
.Y(n_355)
);

XOR2x1_ASAP7_75t_SL g352 ( 
.A(n_325),
.B(n_271),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_355),
.A2(n_349),
.B(n_347),
.Y(n_366)
);

AOI321xp33_ASAP7_75t_L g357 ( 
.A1(n_345),
.A2(n_326),
.A3(n_299),
.B1(n_291),
.B2(n_269),
.C(n_332),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_360),
.Y(n_365)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_273),
.Y(n_372)
);

BUFx4f_ASAP7_75t_SL g362 ( 
.A(n_353),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_348),
.Y(n_367)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_366),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_367),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_363),
.A2(n_354),
.B1(n_352),
.B2(n_237),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_369),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_363),
.A2(n_237),
.B1(n_269),
.B2(n_271),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_343),
.C(n_346),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_371),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_273),
.B1(n_239),
.B2(n_242),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_373),
.C(n_358),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_359),
.A2(n_239),
.B1(n_224),
.B2(n_235),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_378),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_365),
.A2(n_362),
.B(n_182),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_373),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_381),
.A2(n_379),
.B(n_366),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_374),
.A2(n_368),
.B1(n_369),
.B2(n_362),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_382),
.Y(n_384)
);

AOI321xp33_ASAP7_75t_L g385 ( 
.A1(n_383),
.A2(n_379),
.A3(n_380),
.B1(n_377),
.B2(n_382),
.C(n_370),
.Y(n_385)
);

O2A1O1Ixp33_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_384),
.B(n_371),
.C(n_204),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_204),
.Y(n_387)
);


endmodule