module fake_jpeg_13590_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_20),
.A2(n_0),
.B(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_42),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_27),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_24),
.B1(n_17),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_58),
.B1(n_26),
.B2(n_2),
.Y(n_74)
);

OR2x4_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_26),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_21),
.B1(n_17),
.B2(n_23),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_40),
.C(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_40),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_29),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_25),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_69),
.C(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_66),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_74),
.B(n_78),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_34),
.B1(n_26),
.B2(n_3),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_60),
.B1(n_49),
.B2(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_34),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_9),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_76),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_52),
.Y(n_73)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_43),
.C(n_55),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_55),
.C(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_45),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_67),
.B1(n_65),
.B2(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_96),
.B(n_97),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_99),
.B1(n_91),
.B2(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_75),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_88),
.B(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_68),
.B1(n_50),
.B2(n_78),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NOR4xp25_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_88),
.C(n_84),
.D(n_79),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_90),
.C(n_83),
.Y(n_110)
);

AOI21x1_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_107),
.B(n_110),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_105),
.B1(n_95),
.B2(n_84),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_90),
.C(n_80),
.Y(n_107)
);

NOR4xp25_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_84),
.C(n_97),
.D(n_83),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_106),
.A3(n_107),
.B1(n_88),
.B2(n_111),
.C1(n_109),
.C2(n_98),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_102),
.B1(n_94),
.B2(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_115),
.Y(n_118)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_86),
.B(n_77),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_114),
.C(n_112),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_114),
.C(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_86),
.Y(n_124)
);

OAI31xp33_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_121),
.A3(n_7),
.B(n_3),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_0),
.C(n_2),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_4),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_26),
.A3(n_5),
.B1(n_4),
.B2(n_125),
.C1(n_45),
.C2(n_49),
.Y(n_129)
);


endmodule