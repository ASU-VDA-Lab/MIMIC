module real_jpeg_12588_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_4),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_27),
.B1(n_63),
.B2(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_4),
.A2(n_27),
.B1(n_51),
.B2(n_52),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_5),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_160),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_5),
.A2(n_33),
.B1(n_37),
.B2(n_160),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_160),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_7),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_7),
.A2(n_33),
.B1(n_37),
.B2(n_164),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_164),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_8),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_8),
.A2(n_60),
.B(n_63),
.C(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_8),
.B(n_102),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_8),
.B(n_30),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_SL g231 ( 
.A1(n_8),
.A2(n_30),
.B(n_217),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_47),
.C(n_52),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_8),
.A2(n_33),
.B1(n_37),
.B2(n_157),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_8),
.A2(n_86),
.B1(n_87),
.B2(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_8),
.B(n_42),
.Y(n_266)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_10),
.A2(n_33),
.B1(n_37),
.B2(n_67),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_67),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_146),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_11),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_146),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_33),
.B1(n_37),
.B2(n_146),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_146),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_13),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_13),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_13),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_33),
.B1(n_37),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_114)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_103),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_19),
.B(n_103),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.C(n_84),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_20),
.B(n_74),
.CI(n_84),
.CON(n_148),
.SN(n_148)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_58),
.B2(n_73),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_43),
.B2(n_57),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_23),
.B(n_57),
.C(n_58),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_26),
.A2(n_42),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_28),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_SL g218 ( 
.A(n_28),
.B(n_35),
.C(n_37),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_61),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_31),
.A2(n_32),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_31),
.A2(n_32),
.B1(n_163),
.B2(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_31),
.A2(n_112),
.B(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_31),
.A2(n_32),
.B1(n_185),
.B2(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_31),
.A2(n_39),
.B(n_114),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_32),
.A2(n_82),
.B(n_115),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx5_ASAP7_75t_SL g37 ( 
.A(n_33),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_33),
.A2(n_36),
.B(n_216),
.C(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_33),
.B(n_240),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_40),
.B(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_42),
.B(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_43),
.A2(n_57),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_50),
.B(n_54),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_44),
.A2(n_54),
.B(n_96),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_44),
.A2(n_76),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_45),
.A2(n_77),
.B1(n_94),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_45),
.A2(n_77),
.B1(n_212),
.B2(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_45),
.A2(n_77),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_45),
.A2(n_77),
.B1(n_233),
.B2(n_243),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_50),
.A2(n_78),
.B(n_142),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_50),
.B(n_157),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_51),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_73),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_68),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_59),
.A2(n_62),
.B1(n_70),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_59),
.A2(n_70),
.B1(n_159),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_59),
.A2(n_70),
.B1(n_145),
.B2(n_190),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_71)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_69),
.A2(n_102),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_99),
.B(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_70),
.A2(n_145),
.B(n_147),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_74),
.A2(n_75),
.B(n_80),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_91),
.B(n_97),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_97),
.B1(n_98),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_85),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_85),
.A2(n_92),
.B1(n_93),
.B2(n_127),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_89),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_86),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_86),
.A2(n_87),
.B1(n_246),
.B2(n_254),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_86),
.A2(n_136),
.B(n_248),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_87),
.B(n_138),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_87),
.B(n_157),
.Y(n_252)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_90),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_88),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_88),
.A2(n_137),
.B(n_174),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_88),
.A2(n_173),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_90),
.A2(n_173),
.B(n_199),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_102),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_116),
.B2(n_117),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_149),
.B(n_311),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_148),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_124),
.B(n_148),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_129),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_125),
.B(n_128),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_129),
.A2(n_130),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_143),
.C(n_144),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_131),
.A2(n_132),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_133),
.A2(n_134),
.B1(n_139),
.B2(n_140),
.Y(n_283)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_143),
.B(n_144),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_148),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_305),
.B(n_310),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_293),
.B(n_304),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_201),
.B(n_279),
.C(n_292),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_186),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_153),
.B(n_186),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_169),
.C(n_179),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_166),
.C(n_168),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_170),
.B1(n_179),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_176),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_184),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_184),
.B(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_187),
.B(n_194),
.C(n_200),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_195),
.B(n_196),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_277),
.B(n_278),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_221),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_204),
.B(n_207),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_213),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_213),
.B1(n_214),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_219),
.B1(n_220),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_234),
.B(n_276),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_223),
.B(n_226),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_270),
.B(n_275),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_260),
.B(n_269),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_249),
.B(n_259),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_244),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_244),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_241),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_255),
.B(n_258),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_265),
.C(n_268),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_291),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.C(n_284),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_287),
.C(n_290),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_303),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_302),
.C(n_303),
.Y(n_309)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_309),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);


endmodule