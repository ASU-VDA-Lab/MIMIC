module fake_jpeg_20116_n_239 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_25),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_20),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_28),
.B1(n_30),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_71),
.B1(n_76),
.B2(n_0),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_23),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_75),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_36),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_21),
.B1(n_35),
.B2(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_35),
.B1(n_31),
.B2(n_33),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_78),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_81),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_47),
.B1(n_40),
.B2(n_26),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_88),
.Y(n_119)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_36),
.B(n_33),
.C(n_31),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_94),
.B(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_27),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_29),
.B1(n_1),
.B2(n_3),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_101),
.Y(n_127)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_104),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_3),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_10),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_52),
.C(n_61),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_52),
.C(n_51),
.Y(n_117)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_66),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_132),
.B1(n_94),
.B2(n_95),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_51),
.C(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_120),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_106),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_62),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_1),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_5),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_135),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_85),
.B1(n_81),
.B2(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_152),
.B1(n_127),
.B2(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_129),
.C(n_115),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_90),
.B1(n_101),
.B2(n_94),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_154),
.B1(n_110),
.B2(n_8),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_94),
.B1(n_107),
.B2(n_97),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_149),
.B(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

OAI21x1_ASAP7_75t_R g169 ( 
.A1(n_146),
.A2(n_151),
.B(n_128),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_112),
.A2(n_82),
.B(n_88),
.C(n_102),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_111),
.B(n_127),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_83),
.B(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_80),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_84),
.B1(n_99),
.B2(n_7),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_122),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_4),
.B(n_5),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_126),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_120),
.C(n_114),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_166),
.C(n_172),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_162),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_176),
.B1(n_148),
.B2(n_110),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NAND2x1_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_127),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_111),
.C(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_148),
.B1(n_133),
.B2(n_139),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_156),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_109),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_136),
.B1(n_152),
.B2(n_147),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_130),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_187),
.B1(n_189),
.B2(n_164),
.Y(n_195)
);

OAI321xp33_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_155),
.A3(n_147),
.B1(n_144),
.B2(n_154),
.C(n_148),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_192),
.B1(n_194),
.B2(n_174),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_190),
.B1(n_121),
.B2(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_170),
.B(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_167),
.B(n_165),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_205),
.B(n_108),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_204),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_172),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_199),
.C(n_201),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_165),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_206),
.B1(n_193),
.B2(n_187),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_157),
.C(n_173),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_173),
.B(n_176),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_171),
.B1(n_161),
.B2(n_169),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_182),
.Y(n_211)
);

AOI221xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_185),
.B1(n_180),
.B2(n_183),
.C(n_191),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_11),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_185),
.B1(n_169),
.B2(n_130),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_216),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_203),
.B1(n_199),
.B2(n_207),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_203),
.Y(n_220)
);

AOI31xp67_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_224),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_222),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_198),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_217),
.C(n_212),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_214),
.B(n_213),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_SL g230 ( 
.A(n_225),
.B(n_209),
.C(n_210),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_215),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_216),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_227),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_223),
.C(n_219),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_232),
.B(n_233),
.Y(n_236)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_12),
.B(n_11),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_12),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_9),
.B1(n_233),
.B2(n_236),
.Y(n_238)
);


endmodule