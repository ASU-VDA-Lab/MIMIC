module real_jpeg_2697_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_1),
.B(n_96),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_35),
.B(n_50),
.C(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_1),
.B(n_52),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_1),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_62),
.C(n_65),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_1),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_1),
.B(n_84),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_1),
.B(n_119),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_62),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_2),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_62),
.B1(n_66),
.B2(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_30),
.B1(n_35),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_58),
.B1(n_62),
.B2(n_66),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_10),
.A2(n_62),
.B1(n_66),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_10),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_30),
.B1(n_35),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_48),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_12),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_12),
.A2(n_48),
.B1(n_62),
.B2(n_66),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_13),
.A2(n_62),
.B1(n_66),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_13),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_81),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_14),
.A2(n_28),
.B1(n_62),
.B2(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_125),
.B1(n_202),
.B2(n_203),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_18),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_99),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_99),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_88),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_21),
.B(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_44),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_22),
.B(n_46),
.C(n_59),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_25),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_38),
.B(n_39),
.C(n_41),
.Y(n_37)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_26),
.A2(n_33),
.A3(n_35),
.B1(n_40),
.B2(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_29),
.A2(n_108),
.B(n_110),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_30),
.B(n_36),
.Y(n_77)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_50),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_38),
.A2(n_53),
.B(n_56),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_38),
.A2(n_121),
.B(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_52),
.B2(n_57),
.Y(n_46)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_93),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_54),
.B(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_67),
.B(n_70),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_61),
.A2(n_70),
.B(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_61),
.A2(n_133),
.B1(n_151),
.B2(n_163),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_62),
.B(n_181),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_71),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_71),
.A2(n_132),
.B(n_134),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_74),
.B(n_88),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_82),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_82),
.A2(n_83),
.B1(n_155),
.B2(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_83),
.A2(n_98),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_83),
.B(n_142),
.Y(n_157)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_86),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_84),
.A2(n_141),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.C(n_97),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_112),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_104),
.A2(n_106),
.B(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_145),
.B(n_201),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_143),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_143),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.C(n_136),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_136),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_163),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_196),
.B(n_200),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_165),
.B(n_195),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_158),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_158),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_153),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_154),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_177),
.B(n_194),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_188),
.B(n_193),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_183),
.B(n_187),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_186),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_199),
.Y(n_200)
);


endmodule