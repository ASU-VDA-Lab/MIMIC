module fake_jpeg_5586_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx11_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_6),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_3),
.A2(n_4),
.B1(n_6),
.B2(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_9),
.B1(n_8),
.B2(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_1),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_22),
.B(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_10),
.B(n_2),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_24),
.B(n_14),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.C(n_2),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_8),
.C(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_0),
.B(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_28),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_12),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.C(n_33),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_17),
.B1(n_9),
.B2(n_21),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_20),
.A2(n_12),
.B(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_24),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_16),
.B1(n_8),
.B2(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_33),
.B(n_26),
.Y(n_43)
);

NOR2xp67_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_41),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_34),
.B1(n_39),
.B2(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_45),
.B(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_43),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);


endmodule