module fake_jpeg_22281_n_239 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_40),
.B1(n_37),
.B2(n_25),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_29),
.C(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_55),
.B(n_63),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_16),
.B1(n_27),
.B2(n_21),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_64),
.B1(n_24),
.B2(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_26),
.B1(n_31),
.B2(n_22),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_26),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_2),
.B(n_3),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_17),
.B1(n_22),
.B2(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_75),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_76),
.B1(n_64),
.B2(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_18),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_2),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_94),
.B(n_83),
.Y(n_109)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_91),
.Y(n_128)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_97),
.Y(n_115)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_101),
.Y(n_117)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_43),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_66),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_54),
.B1(n_45),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_107),
.B1(n_33),
.B2(n_81),
.Y(n_126)
);

CKINVDCx10_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_38),
.B1(n_35),
.B2(n_49),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_80),
.B1(n_75),
.B2(n_76),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_113),
.B1(n_118),
.B2(n_124),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_112),
.B(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_119),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_123),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_72),
.B(n_57),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_45),
.B1(n_57),
.B2(n_38),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_79),
.B1(n_85),
.B2(n_38),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_125),
.B1(n_129),
.B2(n_95),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_48),
.B1(n_46),
.B2(n_60),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_49),
.C(n_78),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_33),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_46),
.B1(n_65),
.B2(n_60),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_53),
.B1(n_65),
.B2(n_29),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_81),
.B1(n_20),
.B2(n_15),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_90),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_29),
.B1(n_20),
.B2(n_15),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_99),
.B1(n_104),
.B2(n_94),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_99),
.B(n_96),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_137),
.B(n_149),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_100),
.A3(n_95),
.B1(n_86),
.B2(n_33),
.C1(n_101),
.C2(n_97),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_140),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_100),
.B(n_98),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_150),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_145),
.B1(n_147),
.B2(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_101),
.B1(n_81),
.B2(n_33),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_148),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_20),
.B(n_24),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_125),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_108),
.B1(n_126),
.B2(n_113),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_144),
.B1(n_151),
.B2(n_147),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_114),
.B(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_120),
.C(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_122),
.C(n_129),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_167),
.B(n_170),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_134),
.C(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_119),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_122),
.C(n_24),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_148),
.C(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_136),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_186),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_183),
.B1(n_3),
.B2(n_6),
.Y(n_202)
);

CKINVDCx11_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_179),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_181),
.C(n_185),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_137),
.C(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_164),
.B(n_5),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_149),
.B1(n_141),
.B2(n_140),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_143),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_188),
.C(n_159),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_3),
.C(n_4),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_165),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_14),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_155),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_180),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_153),
.C(n_169),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_192),
.C(n_199),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_171),
.C(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_183),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_185),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_154),
.C(n_155),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_156),
.B1(n_164),
.B2(n_6),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_200),
.A2(n_202),
.B1(n_176),
.B2(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_212),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_191),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_182),
.B1(n_176),
.B2(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_193),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_175),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_217),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_218),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_220),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_192),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_189),
.B(n_195),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_203),
.B(n_211),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_179),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_222),
.B(n_224),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_203),
.B(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_212),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_217),
.B1(n_207),
.B2(n_205),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_231),
.A3(n_227),
.B1(n_229),
.B2(n_10),
.C1(n_11),
.C2(n_8),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_7),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_9),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_8),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_233),
.C(n_12),
.Y(n_235)
);

O2A1O1Ixp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_234),
.A2(n_12),
.B(n_13),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_14),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_238),
.Y(n_239)
);


endmodule