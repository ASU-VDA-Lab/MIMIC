module fake_aes_8623_n_646 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_646);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_646;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_18), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_6), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_19), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_11), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_41), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_72), .Y(n_78) );
INVx1_ASAP7_75t_SL g79 ( .A(n_52), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_12), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_65), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_44), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_49), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_43), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_16), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_66), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_33), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_50), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_24), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_61), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_17), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_18), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_42), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_67), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_9), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_39), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_37), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_68), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_58), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_1), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_70), .Y(n_102) );
INVxp33_ASAP7_75t_SL g103 ( .A(n_45), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_25), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_20), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_48), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_35), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_23), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_26), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_22), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_60), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_38), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_51), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_46), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_19), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_36), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_0), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_100), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_89), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
NOR2xp33_ASAP7_75t_R g126 ( .A(n_111), .B(n_29), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_90), .Y(n_127) );
INVx6_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_95), .A2(n_114), .B(n_81), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_91), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_91), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_94), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_109), .B(n_1), .Y(n_134) );
NAND2xp33_ASAP7_75t_R g135 ( .A(n_94), .B(n_30), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
AND3x2_ASAP7_75t_L g141 ( .A(n_88), .B(n_2), .C(n_3), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_107), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_84), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_99), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_107), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_73), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_99), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_108), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_110), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_76), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_110), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_113), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_103), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_88), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_113), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_115), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_128), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_159), .B(n_112), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_121), .B(n_98), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
INVxp67_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_137), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_160), .B(n_93), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
INVxp67_ASAP7_75t_L g177 ( .A(n_131), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_128), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_162), .B(n_93), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_162), .B(n_118), .Y(n_182) );
NOR2xp33_ASAP7_75t_R g183 ( .A(n_132), .B(n_85), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_139), .B(n_115), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_137), .Y(n_185) );
XNOR2xp5_ASAP7_75t_L g186 ( .A(n_156), .B(n_92), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_121), .A2(n_116), .B(n_119), .C(n_117), .Y(n_187) );
INVxp67_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_124), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_125), .B(n_97), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_124), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_145), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_146), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_139), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_144), .B(n_102), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_124), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_124), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_134), .B(n_118), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_149), .B(n_106), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_124), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_146), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_125), .B(n_119), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_129), .B(n_120), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_122), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_145), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_129), .B(n_105), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_148), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_145), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_122), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_123), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_122), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_138), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_148), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_161), .B(n_74), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_138), .B(n_104), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_126), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_140), .B(n_117), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_140), .B(n_116), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_142), .B(n_101), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_175), .B(n_161), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_170), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_206), .B(n_158), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_217), .B(n_158), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_175), .B(n_143), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_175), .B(n_141), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_167), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_183), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_170), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_184), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_172), .B(n_143), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_224), .Y(n_237) );
AND2x6_ASAP7_75t_L g238 ( .A(n_169), .B(n_154), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
INVx4_ASAP7_75t_L g240 ( .A(n_210), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_184), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_163), .Y(n_242) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_181), .B(n_154), .Y(n_243) );
BUFx3_ASAP7_75t_L g244 ( .A(n_163), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_170), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_181), .B(n_153), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_169), .Y(n_247) );
OR2x6_ASAP7_75t_L g248 ( .A(n_224), .B(n_153), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_224), .A2(n_135), .B1(n_151), .B2(n_147), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_166), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_164), .B(n_142), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_198), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_206), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_195), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_201), .A2(n_151), .B1(n_147), .B2(n_155), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_219), .B(n_80), .Y(n_259) );
NAND2xp33_ASAP7_75t_L g260 ( .A(n_223), .B(n_157), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
NOR3xp33_ASAP7_75t_SL g262 ( .A(n_215), .B(n_75), .C(n_96), .Y(n_262) );
INVx5_ASAP7_75t_L g263 ( .A(n_210), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_195), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_207), .B(n_157), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_219), .B(n_157), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_204), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_181), .B(n_155), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_182), .B(n_155), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_204), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_205), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_201), .B(n_79), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_197), .B(n_87), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_205), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
BUFx12f_ASAP7_75t_L g277 ( .A(n_215), .Y(n_277) );
NOR2xp33_ASAP7_75t_R g278 ( .A(n_186), .B(n_2), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_165), .Y(n_279) );
INVx4_ASAP7_75t_L g280 ( .A(n_210), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_182), .B(n_136), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_165), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_219), .A2(n_78), .B1(n_136), .B2(n_127), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_209), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_218), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_177), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_202), .A2(n_127), .B1(n_4), .B2(n_5), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_171), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_250), .B(n_188), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_286), .B(n_207), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_228), .A2(n_194), .B(n_196), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g294 ( .A1(n_243), .A2(n_221), .B1(n_182), .B2(n_222), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_225), .B(n_213), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_243), .A2(n_194), .B1(n_213), .B2(n_220), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_259), .A2(n_213), .B1(n_212), .B2(n_168), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_286), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_267), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_237), .B(n_179), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_267), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_225), .B(n_211), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_248), .A2(n_192), .B1(n_187), .B2(n_208), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_236), .B(n_216), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_248), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_237), .B(n_179), .Y(n_306) );
AOI22x1_ASAP7_75t_L g307 ( .A1(n_228), .A2(n_200), .B1(n_193), .B2(n_190), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_232), .A2(n_189), .B(n_180), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_232), .A2(n_179), .B(n_171), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_248), .A2(n_216), .B1(n_214), .B2(n_208), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_248), .A2(n_214), .B1(n_178), .B2(n_191), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_265), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_236), .B(n_186), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_277), .B(n_178), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_265), .B(n_191), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_239), .B(n_203), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_239), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_231), .B(n_3), .Y(n_319) );
INVx5_ASAP7_75t_L g320 ( .A(n_239), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_239), .Y(n_321) );
INVx5_ASAP7_75t_L g322 ( .A(n_239), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_247), .A2(n_227), .B(n_260), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_238), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_231), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_247), .A2(n_200), .B(n_193), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_231), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_259), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_238), .Y(n_329) );
INVx5_ASAP7_75t_L g330 ( .A(n_241), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_273), .B(n_4), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_256), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_227), .A2(n_185), .B(n_180), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_255), .A2(n_203), .B1(n_199), .B2(n_190), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_238), .B(n_185), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_257), .A2(n_189), .B1(n_199), .B2(n_190), .C(n_203), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_259), .B(n_5), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_238), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g340 ( .A1(n_294), .A2(n_262), .B1(n_251), .B2(n_287), .C(n_283), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_291), .B(n_258), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_305), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_305), .B(n_261), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_320), .B(n_241), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_298), .A2(n_233), .B1(n_230), .B2(n_249), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_333), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_314), .A2(n_266), .B1(n_278), .B2(n_274), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_313), .B(n_256), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_302), .B(n_264), .Y(n_349) );
NAND3xp33_ASAP7_75t_SL g350 ( .A(n_290), .B(n_278), .C(n_229), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_235), .B1(n_241), .B2(n_246), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_308), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_327), .B(n_235), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g355 ( .A1(n_319), .A2(n_241), .B1(n_269), .B2(n_270), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_320), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_319), .A2(n_241), .B1(n_252), .B2(n_253), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_332), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_295), .Y(n_359) );
NOR2xp67_ASAP7_75t_SL g360 ( .A(n_324), .B(n_238), .Y(n_360) );
NAND2x1_ASAP7_75t_L g361 ( .A(n_324), .B(n_238), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g362 ( .A1(n_315), .A2(n_260), .B1(n_264), .B2(n_271), .Y(n_362) );
NAND3x1_ASAP7_75t_L g363 ( .A(n_331), .B(n_288), .C(n_285), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_324), .B(n_271), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_320), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_322), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_328), .A2(n_252), .B1(n_253), .B2(n_272), .Y(n_367) );
OAI211xp5_ASAP7_75t_L g368 ( .A1(n_297), .A2(n_245), .B(n_254), .C(n_226), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_338), .B(n_268), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_316), .B(n_275), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_323), .A2(n_284), .B(n_276), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_341), .B(n_293), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_340), .A2(n_339), .B1(n_329), .B2(n_315), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_349), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_340), .A2(n_301), .B1(n_299), .B2(n_315), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_349), .B(n_322), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_358), .B(n_303), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_350), .A2(n_310), .B1(n_325), .B2(n_312), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_353), .A2(n_307), .B(n_317), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_296), .B1(n_312), .B2(n_316), .Y(n_380) );
OA21x2_ASAP7_75t_L g381 ( .A1(n_353), .A2(n_337), .B(n_292), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_347), .A2(n_252), .B1(n_234), .B2(n_322), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_341), .B(n_306), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_358), .B(n_330), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_359), .A2(n_330), .B1(n_322), .B2(n_280), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_342), .B(n_321), .Y(n_386) );
INVx4_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_359), .A2(n_330), .B1(n_240), .B2(n_280), .Y(n_388) );
AOI22xp5_ASAP7_75t_SL g389 ( .A1(n_342), .A2(n_343), .B1(n_352), .B2(n_351), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_370), .B(n_330), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_352), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_351), .A2(n_329), .B1(n_339), .B2(n_321), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_355), .A2(n_280), .B1(n_240), .B2(n_318), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_369), .A2(n_339), .B1(n_329), .B2(n_311), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_362), .A2(n_300), .B1(n_306), .B2(n_318), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_370), .B(n_300), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_343), .A2(n_240), .B1(n_244), .B2(n_242), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_346), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_395), .A2(n_353), .B(n_371), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_397), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_375), .A2(n_343), .B1(n_363), .B2(n_354), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_348), .B1(n_343), .B2(n_369), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_397), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_391), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_395), .B(n_356), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_399), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_379), .A2(n_371), .B(n_361), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_389), .A2(n_366), .B1(n_365), .B2(n_356), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_374), .B(n_348), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_374), .B(n_368), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_394), .A2(n_335), .B(n_361), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_396), .B(n_365), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_373), .A2(n_365), .B1(n_356), .B2(n_357), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_389), .A2(n_363), .B1(n_364), .B2(n_366), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_399), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_396), .B(n_344), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_387), .B(n_364), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_379), .A2(n_309), .B(n_326), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_387), .B(n_364), .Y(n_421) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_383), .A2(n_364), .B1(n_360), .B2(n_263), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_378), .B(n_367), .C(n_190), .Y(n_423) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_377), .A2(n_360), .B1(n_279), .B2(n_282), .C1(n_289), .C2(n_242), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g425 ( .A1(n_377), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_9), .B3(n_10), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_372), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_372), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_390), .B(n_364), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
OAI211xp5_ASAP7_75t_SL g431 ( .A1(n_382), .A2(n_334), .B(n_336), .C(n_10), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_384), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_390), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_380), .A2(n_336), .B1(n_289), .B2(n_282), .C(n_279), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_427), .B(n_376), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_427), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_417), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_404), .B(n_376), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_417), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_411), .B(n_380), .C(n_392), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_416), .B(n_387), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_416), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_401), .B(n_386), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_405), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_407), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_408), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_433), .B(n_387), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_419), .Y(n_450) );
INVx4_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_408), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_430), .B(n_432), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
XOR2xp5_ASAP7_75t_L g455 ( .A(n_418), .B(n_391), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_426), .B(n_381), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_428), .B(n_381), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_411), .B(n_414), .C(n_423), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_410), .B(n_386), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_403), .B(n_381), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_409), .Y(n_465) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_403), .A2(n_391), .A3(n_393), .B(n_385), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_402), .A2(n_392), .B1(n_388), .B2(n_398), .C(n_203), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_419), .B(n_7), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_413), .B(n_8), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_421), .B(n_11), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_421), .B(n_12), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_429), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_421), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_414), .B(n_13), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_420), .B(n_13), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_422), .B(n_14), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_412), .B(n_15), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_424), .B(n_15), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
AOI33xp33_ASAP7_75t_L g481 ( .A1(n_434), .A2(n_16), .A3(n_17), .B1(n_21), .B2(n_27), .B3(n_28), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_404), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_404), .B(n_190), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_404), .B(n_203), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_456), .B(n_199), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_453), .B(n_199), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_436), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_445), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_441), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_443), .Y(n_493) );
NOR3xp33_ASAP7_75t_SL g494 ( .A(n_462), .B(n_31), .C(n_32), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_443), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_482), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_472), .B(n_199), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_472), .B(n_176), .Y(n_498) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_462), .B(n_34), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_482), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_435), .B(n_176), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_456), .B(n_176), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_458), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_446), .Y(n_504) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_442), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_435), .B(n_176), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_456), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_457), .B(n_176), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_442), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_435), .B(n_174), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_457), .B(n_174), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_174), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_174), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_464), .B(n_174), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_464), .B(n_173), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_453), .B(n_173), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_475), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_453), .B(n_173), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_451), .B(n_53), .Y(n_521) );
INVx5_ASAP7_75t_L g522 ( .A(n_476), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_438), .B(n_173), .Y(n_523) );
AND2x2_ASAP7_75t_SL g524 ( .A(n_451), .B(n_54), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_450), .B(n_173), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_437), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_437), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_437), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_458), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_439), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_450), .B(n_460), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_438), .B(n_55), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_438), .B(n_56), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g534 ( .A(n_480), .B(n_244), .C(n_59), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_469), .B(n_57), .Y(n_535) );
NAND2xp33_ASAP7_75t_SL g536 ( .A(n_468), .B(n_62), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_463), .B(n_63), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g538 ( .A1(n_490), .A2(n_465), .B(n_480), .Y(n_538) );
NOR2xp67_ASAP7_75t_SL g539 ( .A(n_522), .B(n_476), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_508), .B(n_473), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_536), .A2(n_440), .B1(n_535), .B2(n_467), .C(n_534), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_524), .A2(n_479), .B1(n_455), .B2(n_476), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_505), .B(n_451), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_524), .A2(n_479), .B1(n_474), .B2(n_480), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_504), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_532), .A2(n_479), .B1(n_474), .B2(n_480), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g547 ( .A1(n_514), .A2(n_471), .B1(n_470), .B2(n_468), .C1(n_477), .C2(n_478), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_504), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_510), .B(n_470), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_507), .B(n_444), .Y(n_550) );
OAI32xp33_ASAP7_75t_L g551 ( .A1(n_531), .A2(n_469), .A3(n_470), .B1(n_471), .B2(n_455), .Y(n_551) );
OAI32xp33_ASAP7_75t_L g552 ( .A1(n_531), .A2(n_471), .A3(n_477), .B1(n_478), .B2(n_444), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_499), .B(n_481), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_507), .B(n_448), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_492), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_487), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_532), .Y(n_557) );
OAI21xp33_ASAP7_75t_L g558 ( .A1(n_494), .A2(n_449), .B(n_454), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g559 ( .A1(n_537), .A2(n_466), .B1(n_449), .B2(n_454), .C(n_448), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_533), .A2(n_484), .B1(n_483), .B2(n_461), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
AO21x1_ASAP7_75t_L g562 ( .A1(n_521), .A2(n_466), .B(n_483), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_521), .Y(n_563) );
OAI221xp5_ASAP7_75t_SL g564 ( .A1(n_519), .A2(n_461), .B1(n_459), .B2(n_452), .C(n_447), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_522), .B(n_459), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_522), .B(n_447), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
OAI322xp33_ASAP7_75t_L g568 ( .A1(n_519), .A2(n_439), .A3(n_447), .B1(n_452), .B2(n_64), .C1(n_69), .C2(n_71), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_495), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_487), .Y(n_570) );
OA22x2_ASAP7_75t_L g571 ( .A1(n_521), .A2(n_263), .B1(n_452), .B2(n_533), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_522), .B(n_263), .Y(n_572) );
OA21x2_ASAP7_75t_SL g573 ( .A1(n_522), .A2(n_263), .B(n_486), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_497), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_500), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_500), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_491), .B(n_263), .Y(n_577) );
AOI322xp5_ASAP7_75t_L g578 ( .A1(n_491), .A2(n_496), .A3(n_517), .B1(n_516), .B2(n_515), .C1(n_485), .C2(n_530), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_550), .B(n_512), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_570), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_553), .A2(n_520), .B(n_518), .C(n_498), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_554), .B(n_513), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_540), .B(n_513), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_562), .B(n_498), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_543), .Y(n_585) );
XNOR2x1_ASAP7_75t_L g586 ( .A(n_542), .B(n_523), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_549), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_556), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_574), .B(n_509), .Y(n_589) );
AOI211xp5_ASAP7_75t_L g590 ( .A1(n_551), .A2(n_516), .B(n_515), .C(n_517), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_545), .B(n_509), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_571), .B(n_525), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_548), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_541), .B(n_525), .C(n_523), .Y(n_594) );
XNOR2x2_ASAP7_75t_L g595 ( .A(n_544), .B(n_502), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_555), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_559), .B(n_538), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_561), .B(n_502), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_567), .B(n_503), .Y(n_599) );
XNOR2x1_ASAP7_75t_L g600 ( .A(n_544), .B(n_511), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_575), .B(n_503), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_576), .Y(n_603) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_572), .B(n_488), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_568), .B(n_488), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_552), .B(n_529), .Y(n_606) );
XOR2x2_ASAP7_75t_L g607 ( .A(n_546), .B(n_501), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_590), .B(n_578), .Y(n_608) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_584), .A2(n_546), .B(n_547), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_604), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_584), .A2(n_557), .B1(n_563), .B2(n_560), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_580), .Y(n_612) );
XNOR2x1_ASAP7_75t_L g613 ( .A(n_586), .B(n_572), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_580), .B(n_573), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_597), .A2(n_564), .B(n_558), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_594), .A2(n_565), .B(n_566), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g617 ( .A1(n_592), .A2(n_539), .B(n_577), .C(n_501), .Y(n_617) );
OAI21xp33_ASAP7_75t_SL g618 ( .A1(n_606), .A2(n_530), .B(n_528), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_609), .A2(n_587), .B1(n_581), .B2(n_596), .C(n_601), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_612), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_615), .A2(n_600), .B1(n_605), .B2(n_585), .C(n_607), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_618), .B(n_595), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_610), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_612), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_611), .B(n_588), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_611), .A2(n_589), .B(n_579), .C(n_583), .Y(n_626) );
INVx5_ASAP7_75t_L g627 ( .A(n_617), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_614), .A2(n_582), .B1(n_591), .B2(n_598), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_614), .B(n_603), .Y(n_629) );
AOI21xp33_ASAP7_75t_L g630 ( .A1(n_608), .A2(n_593), .B(n_599), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_616), .B(n_602), .C(n_506), .D(n_511), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_613), .A2(n_489), .B1(n_526), .B2(n_527), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_612), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g634 ( .A1(n_615), .A2(n_609), .B(n_611), .C(n_608), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_634), .B(n_619), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_623), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_630), .B(n_628), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_620), .B(n_633), .Y(n_638) );
NAND4xp25_ASAP7_75t_SL g639 ( .A(n_635), .B(n_621), .C(n_626), .D(n_632), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_637), .A2(n_622), .B1(n_625), .B2(n_627), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_638), .A2(n_627), .B1(n_629), .B2(n_631), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_640), .B(n_624), .Y(n_642) );
INVx8_ASAP7_75t_L g643 ( .A(n_639), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_642), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_644), .B(n_641), .C(n_636), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_645), .A2(n_643), .B(n_627), .Y(n_646) );
endmodule