module fake_jpeg_31264_n_153 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_1),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_55),
.C(n_58),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_48),
.B1(n_46),
.B2(n_51),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_4),
.Y(n_117)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_92),
.Y(n_107)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_97),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_60),
.B1(n_47),
.B2(n_46),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_100),
.B1(n_19),
.B2(n_41),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_87),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_20),
.B1(n_44),
.B2(n_42),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_2),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_85),
.C(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_108),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_17),
.B(n_40),
.C(n_38),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_116),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_3),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_4),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_123),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_5),
.CI(n_6),
.CON(n_118),
.SN(n_118)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_6),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_7),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_133),
.B(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_22),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_132),
.B1(n_134),
.B2(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_106),
.B(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_146),
.C(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_145),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_136),
.Y(n_149)
);

AOI322xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_132),
.A3(n_141),
.B1(n_124),
.B2(n_139),
.C1(n_125),
.C2(n_128),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_R g151 ( 
.A(n_150),
.B(n_143),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_127),
.Y(n_153)
);


endmodule