module fake_jpeg_6125_n_238 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_39),
.B(n_59),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_44),
.Y(n_66)
);

NAND2x1_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_10),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_41),
.A2(n_26),
.B(n_20),
.C(n_19),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_54),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_58),
.Y(n_74)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_70),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_30),
.B1(n_33),
.B2(n_26),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_90),
.B1(n_27),
.B2(n_36),
.Y(n_116)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_20),
.B1(n_30),
.B2(n_33),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_16),
.B(n_14),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_28),
.B1(n_24),
.B2(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_24),
.B1(n_36),
.B2(n_27),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_86),
.B1(n_71),
.B2(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_124),
.B1(n_93),
.B2(n_81),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_103),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_36),
.B1(n_27),
.B2(n_17),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_89),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_112),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_119),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_16),
.C(n_15),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_13),
.C(n_12),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_62),
.B1(n_81),
.B2(n_93),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_4),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_92),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_137),
.C(n_2),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_132),
.Y(n_165)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_61),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_62),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_119),
.B1(n_100),
.B2(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_1),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_1),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_117),
.B1(n_121),
.B2(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_68),
.B1(n_82),
.B2(n_94),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_146),
.A2(n_124),
.B1(n_107),
.B2(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_2),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_9),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_158),
.B1(n_160),
.B2(n_164),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_108),
.B(n_110),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_174),
.B(n_150),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_161),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_121),
.B1(n_120),
.B2(n_113),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_168),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_97),
.C(n_103),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_141),
.C(n_145),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_111),
.B1(n_3),
.B2(n_4),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_172),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_133),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_127),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_128),
.A2(n_146),
.B1(n_140),
.B2(n_138),
.Y(n_172)
);

NAND2xp67_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_140),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_180),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_144),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_150),
.B(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_164),
.B1(n_169),
.B2(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_159),
.C(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_148),
.B(n_136),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_154),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_199),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_184),
.A3(n_180),
.B1(n_183),
.B2(n_181),
.C1(n_178),
.C2(n_179),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_206),
.C(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_189),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_184),
.B1(n_180),
.B2(n_177),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_182),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_187),
.C(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_210),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_186),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_202),
.B(n_198),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_213),
.B1(n_197),
.B2(n_200),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_214),
.C(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_185),
.B1(n_170),
.B2(n_173),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_153),
.C(n_170),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_156),
.B1(n_130),
.B2(n_136),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.C(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_209),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_197),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_227),
.B(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_211),
.B1(n_194),
.B2(n_193),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_220),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_230),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_232),
.A2(n_233),
.B(n_208),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_217),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_231),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_234),
.Y(n_238)
);


endmodule