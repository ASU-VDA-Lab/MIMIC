module fake_netlist_5_2332_n_762 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_762);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_762;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_728;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_52),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_77),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_1),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_30),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_117),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_26),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_45),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_89),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_9),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_28),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_53),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_10),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_40),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_111),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_59),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_87),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_18),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_74),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_17),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_82),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_63),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_42),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_65),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_115),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_73),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_38),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_131),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_103),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_22),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_196),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_178),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_155),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_158),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_183),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_204),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_163),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_177),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_0),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_167),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_168),
.B(n_0),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_213),
.B(n_187),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_165),
.B(n_173),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_175),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_218),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_179),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_157),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_208),
.B(n_181),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_165),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_182),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_206),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_185),
.Y(n_278)
);

CKINVDCx8_ASAP7_75t_R g279 ( 
.A(n_237),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_190),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_245),
.A2(n_203),
.B(n_200),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

CKINVDCx8_ASAP7_75t_R g283 ( 
.A(n_232),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_199),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_229),
.B(n_192),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_229),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_207),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_193),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_195),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_197),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_162),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_274),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_198),
.Y(n_304)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_247),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_278),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_292),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_278),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g311 ( 
.A(n_281),
.B(n_286),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_284),
.A2(n_256),
.B1(n_265),
.B2(n_246),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_246),
.B(n_164),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_170),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_271),
.B(n_226),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_23),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_281),
.A2(n_226),
.B1(n_220),
.B2(n_207),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_256),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_24),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_257),
.B(n_220),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_281),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_250),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_250),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_258),
.B(n_2),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_276),
.B(n_25),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

NAND2x1p5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_251),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_268),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_262),
.B(n_27),
.Y(n_337)
);

NAND3x1_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_4),
.C(n_5),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_247),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_268),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_276),
.Y(n_341)
);

INVx4_ASAP7_75t_SL g342 ( 
.A(n_268),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_268),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_343)
);

OAI221xp5_ASAP7_75t_L g344 ( 
.A1(n_253),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_275),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_252),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_283),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_260),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_252),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_252),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_266),
.B(n_29),
.Y(n_352)
);

CKINVDCx8_ASAP7_75t_R g353 ( 
.A(n_289),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_283),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_248),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_347),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_324),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_345),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_296),
.B(n_285),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_316),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_293),
.B(n_253),
.Y(n_364)
);

AO22x2_ASAP7_75t_L g365 ( 
.A1(n_319),
.A2(n_288),
.B1(n_285),
.B2(n_292),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_309),
.Y(n_366)
);

AO22x2_ASAP7_75t_L g367 ( 
.A1(n_319),
.A2(n_288),
.B1(n_287),
.B2(n_291),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_311),
.A2(n_266),
.B1(n_260),
.B2(n_251),
.Y(n_368)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_336),
.B(n_291),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_294),
.B(n_254),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_266),
.B1(n_260),
.B2(n_257),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

NAND2x1p5_ASAP7_75t_L g373 ( 
.A(n_310),
.B(n_289),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_302),
.B(n_266),
.Y(n_374)
);

OR2x6_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_291),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_289),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

OR2x6_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_291),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_297),
.A2(n_254),
.B1(n_289),
.B2(n_15),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_297),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_308),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

OAI221xp5_ASAP7_75t_L g388 ( 
.A1(n_355),
.A2(n_270),
.B1(n_272),
.B2(n_249),
.C(n_252),
.Y(n_388)
);

AO22x2_ASAP7_75t_L g389 ( 
.A1(n_322),
.A2(n_289),
.B1(n_14),
.B2(n_15),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_331),
.A2(n_260),
.B1(n_270),
.B2(n_272),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_354),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_304),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

OR2x6_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_290),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

AO22x2_ASAP7_75t_L g400 ( 
.A1(n_336),
.A2(n_289),
.B1(n_14),
.B2(n_16),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_333),
.Y(n_401)
);

AO22x2_ASAP7_75t_L g402 ( 
.A1(n_343),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_402)
);

OAI221xp5_ASAP7_75t_L g403 ( 
.A1(n_328),
.A2(n_249),
.B1(n_279),
.B2(n_20),
.C(n_21),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_279),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_313),
.A2(n_268),
.B1(n_92),
.B2(n_93),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_300),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_341),
.B(n_268),
.Y(n_408)
);

AO22x2_ASAP7_75t_L g409 ( 
.A1(n_343),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_346),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

NAND2x1p5_ASAP7_75t_L g414 ( 
.A(n_325),
.B(n_31),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_332),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_332),
.B(n_33),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_348),
.B(n_34),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

AO22x2_ASAP7_75t_L g420 ( 
.A1(n_344),
.A2(n_352),
.B1(n_332),
.B2(n_320),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_334),
.A2(n_19),
.B1(n_21),
.B2(n_35),
.Y(n_421)
);

AO22x2_ASAP7_75t_L g422 ( 
.A1(n_352),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_337),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_SL g424 ( 
.A(n_405),
.B(n_353),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_348),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_360),
.B(n_323),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_SL g427 ( 
.A(n_407),
.B(n_323),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_359),
.B(n_334),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_392),
.B(n_323),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_SL g430 ( 
.A(n_378),
.B(n_340),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_383),
.B(n_340),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_303),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_363),
.B(n_340),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_385),
.B(n_342),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_397),
.B(n_342),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_303),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_364),
.B(n_342),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_SL g438 ( 
.A(n_366),
.B(n_339),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_391),
.B(n_339),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_369),
.B(n_306),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_356),
.B(n_306),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_417),
.B(n_306),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_417),
.B(n_306),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_372),
.B(n_303),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g445 ( 
.A(n_358),
.B(n_312),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_364),
.B(n_312),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_370),
.B(n_312),
.Y(n_447)
);

AND2x2_ASAP7_75t_SL g448 ( 
.A(n_421),
.B(n_314),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_370),
.B(n_314),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_314),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_376),
.B(n_329),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_361),
.B(n_329),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_377),
.B(n_305),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_381),
.B(n_330),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_384),
.B(n_330),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_386),
.B(n_393),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_401),
.B(n_305),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_390),
.B(n_41),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_414),
.B(n_305),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_394),
.B(n_44),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_365),
.B(n_398),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g462 ( 
.A(n_394),
.B(n_46),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_373),
.B(n_47),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_395),
.B(n_48),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_395),
.B(n_49),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_371),
.B(n_50),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_396),
.B(n_51),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_396),
.B(n_54),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_406),
.B(n_56),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_374),
.B(n_57),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_368),
.B(n_58),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_410),
.B(n_60),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_SL g473 ( 
.A(n_418),
.B(n_61),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_SL g474 ( 
.A(n_400),
.B(n_64),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_SL g475 ( 
.A(n_400),
.B(n_66),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_413),
.B(n_67),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_68),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_416),
.B(n_69),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_419),
.B(n_70),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_442),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_465),
.B(n_436),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_428),
.B(n_398),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g483 ( 
.A1(n_423),
.A2(n_408),
.B(n_422),
.Y(n_483)
);

AO21x2_ASAP7_75t_L g484 ( 
.A1(n_477),
.A2(n_388),
.B(n_357),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_375),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_440),
.B(n_420),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_387),
.B(n_411),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_450),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_432),
.A2(n_379),
.B(n_422),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_365),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_443),
.A2(n_409),
.B(n_402),
.Y(n_492)
);

AOI221x1_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_367),
.B1(n_382),
.B2(n_389),
.C(n_402),
.Y(n_493)
);

NOR3xp33_ASAP7_75t_L g494 ( 
.A(n_424),
.B(n_403),
.C(n_367),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_466),
.A2(n_382),
.B(n_389),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_454),
.A2(n_71),
.B(n_72),
.Y(n_496)
);

OAI21x1_ASAP7_75t_SL g497 ( 
.A1(n_425),
.A2(n_409),
.B(n_380),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

AOI21x1_ASAP7_75t_SL g499 ( 
.A1(n_453),
.A2(n_380),
.B(n_375),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_455),
.A2(n_75),
.B(n_76),
.Y(n_500)
);

O2A1O1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_451),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_447),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_437),
.B(n_83),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_431),
.A2(n_84),
.B(n_85),
.Y(n_505)
);

AO31x2_ASAP7_75t_L g506 ( 
.A1(n_448),
.A2(n_86),
.A3(n_88),
.B(n_91),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_94),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_434),
.B(n_95),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_449),
.B(n_96),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_433),
.A2(n_97),
.B(n_98),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_426),
.A2(n_99),
.B(n_100),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_461),
.B(n_101),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_459),
.A2(n_104),
.B(n_105),
.Y(n_513)
);

AO31x2_ASAP7_75t_L g514 ( 
.A1(n_475),
.A2(n_106),
.A3(n_107),
.B(n_108),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_109),
.C(n_110),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_439),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_427),
.B(n_112),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_435),
.B(n_114),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_441),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_430),
.A2(n_116),
.B(n_118),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_469),
.B(n_119),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_121),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_457),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_458),
.A2(n_122),
.B(n_123),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_479),
.B(n_126),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_486),
.B(n_429),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_494),
.A2(n_445),
.B1(n_460),
.B2(n_462),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_482),
.A2(n_493),
.B1(n_516),
.B2(n_491),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_504),
.B(n_498),
.Y(n_529)
);

BUFx4f_ASAP7_75t_L g530 ( 
.A(n_498),
.Y(n_530)
);

BUFx2_ASAP7_75t_R g531 ( 
.A(n_491),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_481),
.A2(n_479),
.B(n_467),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_487),
.A2(n_468),
.B(n_463),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_478),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_510),
.A2(n_476),
.B(n_472),
.Y(n_535)
);

AO31x2_ASAP7_75t_L g536 ( 
.A1(n_483),
.A2(n_473),
.A3(n_452),
.B(n_130),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_502),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_511),
.A2(n_127),
.B(n_129),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_134),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_485),
.B(n_135),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_517),
.A2(n_136),
.B(n_138),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_498),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_487),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_492),
.B(n_140),
.Y(n_544)
);

CKINVDCx6p67_ASAP7_75t_R g545 ( 
.A(n_489),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_496),
.A2(n_142),
.B(n_143),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_500),
.A2(n_513),
.B(n_490),
.Y(n_548)
);

OAI221xp5_ASAP7_75t_L g549 ( 
.A1(n_521),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.C(n_148),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_520),
.A2(n_150),
.B(n_151),
.Y(n_550)
);

AO21x2_ASAP7_75t_L g551 ( 
.A1(n_484),
.A2(n_152),
.B(n_497),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_504),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_519),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_480),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_499),
.A2(n_488),
.B(n_524),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_522),
.A2(n_505),
.B(n_495),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_507),
.B(n_523),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_484),
.A2(n_515),
.B(n_522),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_SL g560 ( 
.A1(n_507),
.A2(n_525),
.B1(n_521),
.B2(n_515),
.Y(n_560)
);

OA21x2_ASAP7_75t_L g561 ( 
.A1(n_508),
.A2(n_509),
.B(n_518),
.Y(n_561)
);

AO21x2_ASAP7_75t_L g562 ( 
.A1(n_508),
.A2(n_509),
.B(n_518),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_506),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_501),
.A2(n_506),
.B(n_514),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_506),
.B(n_514),
.Y(n_565)
);

CKINVDCx8_ASAP7_75t_R g566 ( 
.A(n_514),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_486),
.A2(n_391),
.B1(n_359),
.B2(n_315),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_557),
.B(n_552),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_563),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_559),
.Y(n_570)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_560),
.A2(n_527),
.B(n_544),
.C(n_541),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_563),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_548),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_543),
.B(n_546),
.Y(n_574)
);

OA21x2_ASAP7_75t_L g575 ( 
.A1(n_564),
.A2(n_565),
.B(n_548),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_547),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_543),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_565),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_546),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_551),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_547),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_554),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_551),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_555),
.A2(n_532),
.B(n_538),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_537),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_551),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_566),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_539),
.A2(n_549),
.B1(n_534),
.B2(n_526),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_566),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_536),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_553),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_542),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_550),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_550),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_534),
.B(n_539),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_567),
.B(n_533),
.C(n_528),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_555),
.A2(n_532),
.B(n_538),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_531),
.A2(n_529),
.B1(n_530),
.B2(n_545),
.Y(n_600)
);

AOI21x1_ASAP7_75t_L g601 ( 
.A1(n_564),
.A2(n_556),
.B(n_561),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_556),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_561),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_536),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_536),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_561),
.B(n_535),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_530),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_558),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_536),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_562),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_535),
.A2(n_540),
.B(n_536),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_594),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_574),
.B(n_529),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

CKINVDCx8_ASAP7_75t_R g617 ( 
.A(n_582),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_559),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_SL g619 ( 
.A(n_607),
.B(n_529),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_597),
.B(n_545),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_574),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_577),
.B(n_562),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_570),
.B(n_530),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_585),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_585),
.B(n_597),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_582),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_570),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_R g628 ( 
.A(n_589),
.B(n_591),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_590),
.B(n_598),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_R g630 ( 
.A(n_607),
.B(n_589),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_579),
.B(n_593),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_588),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_R g633 ( 
.A(n_591),
.B(n_578),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_R g634 ( 
.A(n_575),
.B(n_593),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_579),
.B(n_578),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_579),
.B(n_571),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_569),
.B(n_572),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_R g638 ( 
.A(n_575),
.B(n_576),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_R g639 ( 
.A(n_601),
.B(n_604),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_613),
.B(n_610),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_569),
.B(n_572),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_592),
.B(n_605),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_592),
.B(n_605),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_R g644 ( 
.A(n_575),
.B(n_576),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_R g645 ( 
.A(n_575),
.B(n_576),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_611),
.B(n_612),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_611),
.B(n_612),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_604),
.B(n_610),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_611),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_606),
.B(n_596),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_622),
.B(n_612),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_617),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_635),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_622),
.B(n_603),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_625),
.B(n_603),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_625),
.B(n_586),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_637),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_646),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_650),
.B(n_602),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_626),
.B(n_609),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_649),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_636),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_642),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_629),
.B(n_595),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_637),
.B(n_586),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_636),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_650),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_641),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_639),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_643),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_641),
.B(n_586),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_631),
.B(n_609),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_648),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_631),
.B(n_609),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_633),
.A2(n_587),
.B1(n_580),
.B2(n_583),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_624),
.B(n_608),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_654),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_654),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_663),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_616),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_668),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_655),
.B(n_640),
.Y(n_682)
);

INVxp33_ASAP7_75t_SL g683 ( 
.A(n_652),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_652),
.B(n_632),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_676),
.B(n_608),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_655),
.B(n_647),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_651),
.B(n_580),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_657),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_667),
.B(n_624),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_663),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_682),
.B(n_667),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_683),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_677),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_677),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_683),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_680),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_679),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_678),
.B(n_676),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_681),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_678),
.A2(n_662),
.B1(n_666),
.B2(n_628),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_696),
.B(n_686),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_L g702 ( 
.A1(n_692),
.A2(n_662),
.B1(n_666),
.B2(n_652),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_695),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_L g704 ( 
.A1(n_691),
.A2(n_684),
.B1(n_664),
.B2(n_620),
.C(n_618),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_698),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_704),
.A2(n_700),
.B(n_691),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_702),
.A2(n_662),
.B1(n_666),
.B2(n_699),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_703),
.A2(n_662),
.B1(n_666),
.B2(n_699),
.Y(n_708)
);

XNOR2x1_ASAP7_75t_L g709 ( 
.A(n_701),
.B(n_627),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_705),
.B(n_689),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_705),
.Y(n_711)
);

O2A1O1Ixp5_ASAP7_75t_L g712 ( 
.A1(n_706),
.A2(n_697),
.B(n_688),
.C(n_690),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_711),
.B(n_689),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_709),
.B(n_694),
.Y(n_714)
);

AOI32xp33_ASAP7_75t_L g715 ( 
.A1(n_708),
.A2(n_669),
.A3(n_675),
.B1(n_689),
.B2(n_686),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_714),
.B(n_707),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_713),
.B(n_710),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_715),
.B(n_693),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_716),
.B(n_712),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_718),
.B(n_717),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_716),
.B(n_698),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_716),
.B(n_688),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_720),
.B(n_614),
.Y(n_723)
);

NAND4xp75_ASAP7_75t_L g724 ( 
.A(n_719),
.B(n_623),
.C(n_667),
.D(n_660),
.Y(n_724)
);

AO21x1_ASAP7_75t_L g725 ( 
.A1(n_721),
.A2(n_619),
.B(n_634),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_722),
.B(n_668),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_721),
.Y(n_727)
);

AND5x1_ASAP7_75t_L g728 ( 
.A(n_719),
.B(n_630),
.C(n_669),
.D(n_675),
.E(n_645),
.Y(n_728)
);

NOR4xp25_ASAP7_75t_L g729 ( 
.A(n_719),
.B(n_658),
.C(n_660),
.D(n_587),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_727),
.A2(n_583),
.B(n_661),
.C(n_657),
.Y(n_730)
);

XNOR2x1_ASAP7_75t_L g731 ( 
.A(n_724),
.B(n_615),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_723),
.B(n_668),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_726),
.A2(n_668),
.B1(n_685),
.B2(n_621),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_725),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_729),
.A2(n_613),
.B(n_658),
.Y(n_735)
);

AOI221xp5_ASAP7_75t_L g736 ( 
.A1(n_728),
.A2(n_661),
.B1(n_653),
.B2(n_687),
.C(n_659),
.Y(n_736)
);

INVxp33_ASAP7_75t_L g737 ( 
.A(n_731),
.Y(n_737)
);

OR3x2_ASAP7_75t_L g738 ( 
.A(n_734),
.B(n_685),
.C(n_653),
.Y(n_738)
);

XOR2x1_ASAP7_75t_L g739 ( 
.A(n_732),
.B(n_615),
.Y(n_739)
);

NAND4xp75_ASAP7_75t_L g740 ( 
.A(n_736),
.B(n_687),
.C(n_671),
.D(n_665),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_733),
.B(n_671),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_730),
.B(n_673),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_735),
.A2(n_659),
.B1(n_665),
.B2(n_673),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_R g744 ( 
.A(n_737),
.B(n_644),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_743),
.B(n_659),
.Y(n_745)
);

XNOR2xp5_ASAP7_75t_L g746 ( 
.A(n_739),
.B(n_656),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_742),
.B(n_659),
.Y(n_747)
);

XNOR2xp5_ASAP7_75t_L g748 ( 
.A(n_740),
.B(n_656),
.Y(n_748)
);

XNOR2xp5_ASAP7_75t_L g749 ( 
.A(n_746),
.B(n_741),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_744),
.B(n_738),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_748),
.Y(n_751)
);

OAI211xp5_ASAP7_75t_L g752 ( 
.A1(n_747),
.A2(n_670),
.B(n_595),
.C(n_596),
.Y(n_752)
);

AO21x1_ASAP7_75t_L g753 ( 
.A1(n_750),
.A2(n_745),
.B(n_638),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_SL g754 ( 
.A1(n_749),
.A2(n_670),
.B(n_672),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_751),
.B1(n_752),
.B2(n_606),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_753),
.Y(n_756)
);

AOI31xp33_ASAP7_75t_L g757 ( 
.A1(n_756),
.A2(n_674),
.A3(n_672),
.B(n_651),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_757),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_758),
.A2(n_755),
.B(n_576),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_759),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_581),
.B1(n_608),
.B2(n_602),
.C(n_573),
.Y(n_761)
);

AOI211xp5_ASAP7_75t_L g762 ( 
.A1(n_761),
.A2(n_584),
.B(n_599),
.C(n_674),
.Y(n_762)
);


endmodule