module fake_jpeg_2026_n_212 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_25),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_26),
.B1(n_21),
.B2(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_56),
.B1(n_69),
.B2(n_44),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_26),
.B1(n_21),
.B2(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_29),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_35),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_71),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_25),
.B1(n_28),
.B2(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_23),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_50),
.C(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_21),
.B1(n_34),
.B2(n_32),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_70),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_27),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_46),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_80),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_81),
.Y(n_116)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_98),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_97),
.B1(n_65),
.B2(n_68),
.Y(n_114)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_35),
.B(n_31),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_70),
.C(n_27),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_50),
.B1(n_40),
.B2(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_63),
.B(n_70),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_118),
.B(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_125),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_61),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_84),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_97),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_67),
.B1(n_54),
.B2(n_66),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_51),
.B(n_18),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_14),
.Y(n_125)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_131),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_77),
.B(n_97),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_110),
.B(n_113),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_133),
.B(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_77),
.C(n_85),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_118),
.C(n_115),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_92),
.B1(n_101),
.B2(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_79),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_87),
.C(n_102),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_141),
.B(n_144),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_96),
.B(n_51),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_66),
.B1(n_55),
.B2(n_76),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_96),
.B(n_55),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_147),
.B(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_159),
.C(n_160),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_123),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_116),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_115),
.C(n_105),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_161),
.B(n_164),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_116),
.A3(n_112),
.B1(n_117),
.B2(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_145),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_144),
.B(n_143),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_124),
.C(n_110),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_173),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_133),
.B1(n_129),
.B2(n_143),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_172),
.B1(n_175),
.B2(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_141),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_140),
.B1(n_139),
.B2(n_127),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_119),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_147),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_145),
.B1(n_142),
.B2(n_124),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_159),
.C(n_176),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_182),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_156),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_183),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_161),
.C(n_150),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_148),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_148),
.C(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_165),
.B1(n_152),
.B2(n_172),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_162),
.B(n_153),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_8),
.B(n_12),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_16),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_12),
.B(n_13),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_189),
.B(n_180),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_178),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_203),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_196),
.A3(n_194),
.B1(n_184),
.B2(n_181),
.C1(n_183),
.C2(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_206),
.B(n_195),
.CI(n_13),
.CON(n_208),
.SN(n_208)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_207),
.B(n_14),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_6),
.A3(n_15),
.B1(n_16),
.B2(n_208),
.C1(n_209),
.C2(n_199),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_15),
.Y(n_212)
);


endmodule