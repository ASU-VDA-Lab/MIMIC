module fake_ibex_1156_n_5977 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_974, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_960, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_979, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_983, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_5977);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_974;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_960;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_979;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_983;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_5977;

wire n_4557;
wire n_5285;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_5591;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_5673;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_1865;
wire n_5033;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_5612;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_5252;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_5099;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_5719;
wire n_5157;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_5959;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_3339;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_5566;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_1072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_3096;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5824;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_5403;
wire n_985;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_4686;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_4733;
wire n_5368;
wire n_987;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4797;
wire n_4493;
wire n_1082;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_1012;
wire n_4412;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_5506;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_5319;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5543;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_5796;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_5854;
wire n_4067;
wire n_4997;
wire n_5906;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_5828;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3788;
wire n_3448;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_1312;
wire n_5844;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_5294;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_3394;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_4991;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_3703;
wire n_5116;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_5953;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_998;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_5193;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_5153;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_5399;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_5096;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_5778;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_5208;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_5644;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_1442;
wire n_2168;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_5940;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_5324;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_5184;
wire n_5747;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_5618;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3819;
wire n_3334;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_5464;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_5688;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_5804;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_5123;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_1003;
wire n_2708;
wire n_5164;
wire n_2748;
wire n_5359;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_1076;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_3284;
wire n_2875;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_994;
wire n_5136;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_1839;
wire n_5160;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_5313;
wire n_2108;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_5744;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_5715;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_5558;
wire n_2157;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_5708;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_5853;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_5592;
wire n_5484;
wire n_4982;
wire n_5418;
wire n_5432;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_3989;
wire n_5565;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_5293;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5533;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_4912;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_5479;
wire n_5598;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_4311;
wire n_5766;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_5279;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_5613;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_5897;
wire n_5331;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_3624;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1464;
wire n_1566;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_2252;
wire n_1982;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_1009;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2991;
wire n_2699;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5819;
wire n_5855;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_2990;
wire n_3449;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5105;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_5846;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2187;
wire n_2105;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_4149;
wire n_3930;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_993;
wire n_5409;
wire n_2581;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_1088;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_5761;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_5298;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_4811;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_5965;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4595;
wire n_4418;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_5507;
wire n_1164;
wire n_3749;
wire n_5470;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_5963;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_37),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_413),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_517),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_240),
.Y(n_987)
);

CKINVDCx16_ASAP7_75t_R g988 ( 
.A(n_864),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_736),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_983),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_880),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_253),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_115),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_367),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_275),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_220),
.Y(n_996)
);

BUFx10_ASAP7_75t_L g997 ( 
.A(n_473),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_900),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_751),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_41),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_446),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_930),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_525),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_664),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_660),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_433),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_242),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_935),
.Y(n_1008)
);

CKINVDCx14_ASAP7_75t_R g1009 ( 
.A(n_258),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_349),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_656),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_707),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_499),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_344),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_337),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_542),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_641),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_297),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_541),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_471),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_856),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_277),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_693),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_707),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_438),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_146),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_455),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_936),
.Y(n_1028)
);

CKINVDCx16_ASAP7_75t_R g1029 ( 
.A(n_519),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_678),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_973),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_559),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_760),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_852),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_425),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_244),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_9),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_164),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_585),
.Y(n_1039)
);

CKINVDCx14_ASAP7_75t_R g1040 ( 
.A(n_903),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_174),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_931),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_871),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_426),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_290),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_676),
.Y(n_1046)
);

BUFx10_ASAP7_75t_L g1047 ( 
.A(n_649),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_361),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_419),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_845),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_932),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_512),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_58),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_256),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_910),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_883),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_115),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_534),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_159),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_645),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_541),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_886),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_920),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_926),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_656),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_927),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_898),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_704),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_74),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_275),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_948),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_812),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_26),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_756),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_954),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_885),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_964),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_602),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_102),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_228),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_174),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_928),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_575),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_488),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_689),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_849),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_866),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_420),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_853),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_242),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_158),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_62),
.Y(n_1092)
);

BUFx10_ASAP7_75t_L g1093 ( 
.A(n_855),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_413),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_837),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_301),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_125),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_885),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_854),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_757),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_612),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_965),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_202),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_521),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_755),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_879),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_54),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_783),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_983),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_850),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_943),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_348),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_893),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_717),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_57),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_664),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_810),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_864),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_665),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_742),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_851),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_770),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_354),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_54),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_103),
.Y(n_1125)
);

BUFx2_ASAP7_75t_SL g1126 ( 
.A(n_937),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_901),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_965),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_661),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_480),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_423),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_571),
.Y(n_1132)
);

INVxp33_ASAP7_75t_R g1133 ( 
.A(n_289),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_842),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_403),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_915),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_929),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_877),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_887),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_272),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_547),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_484),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_65),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_128),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_937),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_891),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_336),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_817),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_970),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_963),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_324),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_899),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_212),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_659),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_181),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_972),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_197),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_102),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_665),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_413),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_366),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_297),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_967),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_433),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_683),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_746),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_724),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_223),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_555),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_284),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_725),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_402),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_891),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_614),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_982),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_960),
.Y(n_1176)
);

BUFx2_ASAP7_75t_SL g1177 ( 
.A(n_834),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_447),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_25),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_635),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_266),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_250),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_386),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_893),
.Y(n_1184)
);

BUFx8_ASAP7_75t_SL g1185 ( 
.A(n_889),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_248),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_414),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_972),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_591),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_803),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_946),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_938),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_493),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_884),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_799),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_907),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_312),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_481),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_780),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_8),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_906),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_897),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_744),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_89),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_690),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_386),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_781),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_757),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_667),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_905),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_941),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_919),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_424),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_592),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_951),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_556),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_941),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_456),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_869),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_47),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_680),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_104),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_464),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_909),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_101),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_528),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_331),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_982),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_341),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_508),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_111),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_188),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_888),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_890),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_842),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_21),
.Y(n_1236)
);

INVxp67_ASAP7_75t_SL g1237 ( 
.A(n_427),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_754),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_260),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_969),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_636),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_491),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_158),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_265),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_415),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_876),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_673),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_576),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_327),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_7),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_27),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_347),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_156),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_736),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_841),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_718),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_870),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_330),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_25),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_54),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_563),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_325),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_769),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_956),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_632),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_107),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_814),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_959),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_291),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_685),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_132),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_506),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_276),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_79),
.Y(n_1274)
);

BUFx10_ASAP7_75t_L g1275 ( 
.A(n_774),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_290),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_178),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_860),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_836),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_632),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_925),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_208),
.Y(n_1282)
);

CKINVDCx14_ASAP7_75t_R g1283 ( 
.A(n_255),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_923),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_508),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_369),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_878),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_968),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_256),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_144),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_943),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_300),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_550),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_750),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_659),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_192),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_811),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_192),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_698),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_847),
.Y(n_1300)
);

BUFx8_ASAP7_75t_SL g1301 ( 
.A(n_724),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_555),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_582),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_952),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_206),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_892),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_731),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_296),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_482),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_439),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_322),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_550),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_666),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_921),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_539),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_517),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_530),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_536),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_623),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_551),
.Y(n_1320)
);

BUFx8_ASAP7_75t_SL g1321 ( 
.A(n_450),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_28),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_36),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_569),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_862),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_874),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_928),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_942),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_825),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_729),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_698),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_258),
.Y(n_1332)
);

CKINVDCx16_ASAP7_75t_R g1333 ( 
.A(n_130),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_240),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_763),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_73),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_970),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_433),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_795),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_657),
.Y(n_1340)
);

CKINVDCx16_ASAP7_75t_R g1341 ( 
.A(n_227),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_135),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_214),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_615),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_670),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_371),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_23),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_60),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_914),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_902),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_848),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_272),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_833),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_979),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_681),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_509),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_588),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_349),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_374),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_594),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_87),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_0),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_684),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_846),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_355),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_663),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_525),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_828),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_19),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_57),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_157),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_916),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_541),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_772),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_124),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_726),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_875),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_955),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_51),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_182),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_677),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_678),
.Y(n_1382)
);

BUFx10_ASAP7_75t_L g1383 ( 
.A(n_945),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_185),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_168),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_957),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_625),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_699),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_909),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_980),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_895),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_77),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_119),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_798),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_674),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_482),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_766),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_745),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_963),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_873),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_555),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_861),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_978),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_859),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_545),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_370),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_939),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_922),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_279),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_211),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_718),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_644),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_949),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_855),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_740),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_160),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_315),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_679),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_959),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_239),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_460),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_281),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_460),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_609),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_657),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_512),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_453),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_597),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_561),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_241),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_953),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_9),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_507),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_819),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_960),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_326),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_722),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_694),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_911),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_872),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_114),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_253),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_491),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_503),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_140),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_826),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_19),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_311),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_940),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_734),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_917),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_916),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_616),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_406),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_418),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_935),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_849),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_723),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_899),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_583),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_882),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_313),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_913),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_950),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_868),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_426),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_585),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_976),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_389),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_857),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_562),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_434),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_904),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_923),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_384),
.Y(n_1475)
);

BUFx10_ASAP7_75t_L g1476 ( 
.A(n_24),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_206),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_776),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_449),
.Y(n_1479)
);

CKINVDCx14_ASAP7_75t_R g1480 ( 
.A(n_931),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_273),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_858),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_5),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_971),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_964),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_958),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_213),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_11),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_449),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_934),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_195),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_215),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_690),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_37),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_980),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_472),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_850),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_61),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_658),
.Y(n_1499)
);

BUFx2_ASAP7_75t_SL g1500 ( 
.A(n_277),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_142),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_874),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_384),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_73),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_587),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_902),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_908),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_667),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_870),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_643),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_513),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_282),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_383),
.Y(n_1513)
);

BUFx8_ASAP7_75t_SL g1514 ( 
.A(n_160),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_624),
.Y(n_1515)
);

BUFx10_ASAP7_75t_L g1516 ( 
.A(n_39),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_51),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_468),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_346),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_962),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_591),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_241),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_646),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_922),
.Y(n_1524)
);

BUFx5_ASAP7_75t_L g1525 ( 
.A(n_947),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_799),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_268),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_88),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_5),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_402),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_514),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_865),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_141),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_815),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_816),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_826),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_802),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_788),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_918),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_0),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_961),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_725),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_131),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_348),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_357),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_197),
.Y(n_1546)
);

CKINVDCx16_ASAP7_75t_R g1547 ( 
.A(n_720),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_58),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_486),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_181),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_641),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_809),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_350),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_52),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_22),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_827),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_876),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_714),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_711),
.Y(n_1559)
);

BUFx5_ASAP7_75t_L g1560 ( 
.A(n_318),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_30),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_881),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_178),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_543),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_975),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_62),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_867),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_914),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_912),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_924),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_329),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_944),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_232),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_188),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_801),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_894),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_953),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_966),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_575),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_816),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_377),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_933),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_627),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_253),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_703),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_480),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_368),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_791),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_308),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_968),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_401),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_199),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_554),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_974),
.Y(n_1594)
);

BUFx8_ASAP7_75t_SL g1595 ( 
.A(n_896),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_863),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_145),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_371),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_398),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_574),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_927),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1009),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1009),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_989),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1321),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_989),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1085),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_984),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1085),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1223),
.Y(n_1610)
);

CKINVDCx16_ASAP7_75t_R g1611 ( 
.A(n_1029),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1155),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1491),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1522),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_997),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1548),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1311),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1519),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_985),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_985),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1230),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1321),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1296),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1283),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1322),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_994),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1525),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_995),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1283),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1079),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_991),
.B(n_0),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1010),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1020),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1022),
.Y(n_1634)
);

CKINVDCx16_ASAP7_75t_R g1635 ( 
.A(n_1049),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1525),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1079),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1384),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1032),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1038),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1053),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1091),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1097),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1103),
.Y(n_1644)
);

BUFx10_ASAP7_75t_L g1645 ( 
.A(n_1137),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1112),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1525),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1384),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1115),
.Y(n_1649)
);

CKINVDCx16_ASAP7_75t_R g1650 ( 
.A(n_1200),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1143),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1051),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1147),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1158),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1161),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1561),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1170),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1181),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1514),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1514),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1116),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1183),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_1561),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1573),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1186),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1213),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1225),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1227),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1525),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1573),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1232),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1525),
.Y(n_1672)
);

INVxp33_ASAP7_75t_L g1673 ( 
.A(n_1478),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1242),
.Y(n_1674)
);

INVxp67_ASAP7_75t_SL g1675 ( 
.A(n_1057),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1248),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1019),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1333),
.Y(n_1678)
);

INVxp33_ASAP7_75t_SL g1679 ( 
.A(n_992),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1249),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_997),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1250),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1260),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1525),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1040),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1261),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1266),
.Y(n_1687)
);

INVxp33_ASAP7_75t_L g1688 ( 
.A(n_1004),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1057),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1480),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1272),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1094),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1341),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1094),
.Y(n_1694)
);

INVxp67_ASAP7_75t_SL g1695 ( 
.A(n_1140),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1276),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1140),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1285),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1298),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1308),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1310),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1525),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1027),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1315),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1193),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1316),
.Y(n_1706)
);

BUFx2_ASAP7_75t_SL g1707 ( 
.A(n_997),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1318),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1040),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1324),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1334),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1342),
.Y(n_1712)
);

INVxp33_ASAP7_75t_SL g1713 ( 
.A(n_993),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1193),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1050),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1346),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1352),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1560),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1361),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1367),
.Y(n_1720)
);

INVxp33_ASAP7_75t_SL g1721 ( 
.A(n_996),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1369),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1027),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1370),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1371),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1409),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1480),
.Y(n_1727)
);

INVxp33_ASAP7_75t_SL g1728 ( 
.A(n_1000),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1106),
.B(n_1),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1560),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1422),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1432),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1560),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1436),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1447),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1615),
.A2(n_1677),
.B1(n_1693),
.B2(n_1678),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1630),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1630),
.Y(n_1738)
);

AND2x6_ASAP7_75t_L g1739 ( 
.A(n_1615),
.B(n_1050),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1715),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1627),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1637),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1637),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1718),
.A2(n_1320),
.B(n_1309),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1645),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1648),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1648),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1608),
.B(n_1069),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1629),
.B(n_1407),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1730),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1611),
.A2(n_1006),
.B1(n_1007),
.B2(n_1001),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1679),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1608),
.B(n_1069),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1645),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1681),
.B(n_1570),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1733),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1677),
.A2(n_1338),
.B1(n_1359),
.B2(n_1271),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1604),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1606),
.Y(n_1759)
);

OAI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1636),
.A2(n_1320),
.B(n_1309),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1713),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1659),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1647),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1607),
.Y(n_1764)
);

BUFx8_ASAP7_75t_L g1765 ( 
.A(n_1621),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1721),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1670),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1681),
.B(n_1013),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1612),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1609),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1669),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1672),
.A2(n_1362),
.B(n_1348),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1684),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1702),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1670),
.Y(n_1775)
);

INVx6_ASAP7_75t_L g1776 ( 
.A(n_1635),
.Y(n_1776)
);

CKINVDCx6p67_ASAP7_75t_R g1777 ( 
.A(n_1650),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1619),
.Y(n_1778)
);

BUFx12f_ASAP7_75t_L g1779 ( 
.A(n_1602),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1610),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1603),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1613),
.Y(n_1782)
);

OA21x2_ASAP7_75t_L g1783 ( 
.A1(n_1638),
.A2(n_1362),
.B(n_1348),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1614),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1638),
.Y(n_1785)
);

OA21x2_ASAP7_75t_L g1786 ( 
.A1(n_1656),
.A2(n_1483),
.B(n_1441),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1656),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1612),
.B(n_1069),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1620),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1663),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1616),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1626),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1628),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1664),
.Y(n_1794)
);

BUFx12f_ASAP7_75t_L g1795 ( 
.A(n_1624),
.Y(n_1795)
);

OA21x2_ASAP7_75t_L g1796 ( 
.A1(n_1735),
.A2(n_1483),
.B(n_1441),
.Y(n_1796)
);

INVx4_ASAP7_75t_L g1797 ( 
.A(n_1685),
.Y(n_1797)
);

BUFx12f_ASAP7_75t_L g1798 ( 
.A(n_1690),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1623),
.B(n_1135),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1632),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1633),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1675),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1617),
.B(n_1241),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1728),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1634),
.A2(n_1498),
.B(n_1487),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1639),
.Y(n_1806)
);

INVx5_ASAP7_75t_L g1807 ( 
.A(n_1707),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1640),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1641),
.Y(n_1809)
);

BUFx8_ASAP7_75t_SL g1810 ( 
.A(n_1605),
.Y(n_1810)
);

OA21x2_ASAP7_75t_L g1811 ( 
.A1(n_1642),
.A2(n_1498),
.B(n_1487),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1643),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1644),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1689),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1692),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1652),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1646),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1694),
.B(n_1695),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1697),
.B(n_1016),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1618),
.B(n_1412),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1625),
.B(n_1661),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1705),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1703),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1714),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1709),
.B(n_1439),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1673),
.B(n_1135),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1649),
.Y(n_1827)
);

OAI22x1_ASAP7_75t_SL g1828 ( 
.A1(n_1723),
.A2(n_1338),
.B1(n_1359),
.B2(n_1271),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1651),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1727),
.B(n_1560),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1653),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1622),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1654),
.Y(n_1833)
);

BUFx12f_ASAP7_75t_L g1834 ( 
.A(n_1660),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1655),
.B(n_1018),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1657),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1658),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1662),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_L g1839 ( 
.A(n_1665),
.B(n_1560),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1688),
.Y(n_1840)
);

INVx4_ASAP7_75t_L g1841 ( 
.A(n_1666),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1667),
.B(n_1025),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1668),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1671),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1674),
.Y(n_1845)
);

NAND2x1p5_ASAP7_75t_L g1846 ( 
.A(n_1676),
.B(n_1082),
.Y(n_1846)
);

CKINVDCx16_ASAP7_75t_R g1847 ( 
.A(n_1631),
.Y(n_1847)
);

INVx5_ASAP7_75t_L g1848 ( 
.A(n_1729),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1680),
.B(n_1464),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1682),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1683),
.B(n_1135),
.Y(n_1851)
);

BUFx12f_ASAP7_75t_L g1852 ( 
.A(n_1734),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1686),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1687),
.B(n_1507),
.Y(n_1854)
);

OAI22x1_ASAP7_75t_R g1855 ( 
.A1(n_1691),
.A2(n_987),
.B1(n_1096),
.B2(n_1014),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_1696),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1698),
.Y(n_1857)
);

CKINVDCx16_ASAP7_75t_R g1858 ( 
.A(n_1699),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1700),
.Y(n_1859)
);

INVx4_ASAP7_75t_L g1860 ( 
.A(n_1701),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1704),
.A2(n_1708),
.B1(n_1710),
.B2(n_1706),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1711),
.Y(n_1862)
);

BUFx12f_ASAP7_75t_L g1863 ( 
.A(n_1732),
.Y(n_1863)
);

BUFx8_ASAP7_75t_SL g1864 ( 
.A(n_1712),
.Y(n_1864)
);

CKINVDCx6p67_ASAP7_75t_R g1865 ( 
.A(n_1716),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1717),
.A2(n_1035),
.B1(n_1036),
.B2(n_1026),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1719),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1720),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1722),
.A2(n_1041),
.B1(n_1044),
.B2(n_1037),
.Y(n_1869)
);

XNOR2x2_ASAP7_75t_L g1870 ( 
.A(n_1724),
.B(n_986),
.Y(n_1870)
);

OAI21x1_ASAP7_75t_L g1871 ( 
.A1(n_1725),
.A2(n_1528),
.B(n_1504),
.Y(n_1871)
);

INVx5_ASAP7_75t_L g1872 ( 
.A(n_1726),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1731),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1630),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1629),
.B(n_1045),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1629),
.B(n_1048),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1715),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1630),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1715),
.Y(n_1879)
);

INVx5_ASAP7_75t_L g1880 ( 
.A(n_1645),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1608),
.B(n_1476),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1659),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1629),
.B(n_988),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1630),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1715),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1629),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1715),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1611),
.A2(n_1054),
.B1(n_1058),
.B2(n_1052),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1645),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1608),
.B(n_1476),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1645),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1611),
.A2(n_1061),
.B1(n_1070),
.B2(n_1059),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1715),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1615),
.A2(n_1080),
.B1(n_1083),
.B2(n_1073),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1718),
.A2(n_1528),
.B(n_1504),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1630),
.Y(n_1896)
);

INVx5_ASAP7_75t_L g1897 ( 
.A(n_1645),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1715),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1629),
.B(n_1084),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1678),
.Y(n_1900)
);

BUFx8_ASAP7_75t_SL g1901 ( 
.A(n_1605),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1629),
.B(n_1088),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1645),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1715),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1715),
.Y(n_1905)
);

BUFx12f_ASAP7_75t_L g1906 ( 
.A(n_1659),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1715),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1630),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1629),
.B(n_1090),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1630),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1703),
.A2(n_1172),
.B1(n_1178),
.B2(n_1132),
.Y(n_1911)
);

INVx2_ASAP7_75t_SL g1912 ( 
.A(n_1629),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1715),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1608),
.B(n_1476),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1630),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1715),
.Y(n_1916)
);

BUFx6f_ASAP7_75t_L g1917 ( 
.A(n_1715),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1659),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1715),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1630),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1715),
.Y(n_1921)
);

OA21x2_ASAP7_75t_L g1922 ( 
.A1(n_1718),
.A2(n_1471),
.B(n_1462),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1629),
.B(n_1092),
.Y(n_1923)
);

INVx5_ASAP7_75t_L g1924 ( 
.A(n_1645),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1715),
.Y(n_1925)
);

AND2x2_ASAP7_75t_SL g1926 ( 
.A(n_1611),
.B(n_998),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1645),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1715),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1715),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1715),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1629),
.B(n_1104),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1645),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1629),
.Y(n_1933)
);

BUFx8_ASAP7_75t_L g1934 ( 
.A(n_1629),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1629),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1715),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1630),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1615),
.B(n_1516),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1715),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1629),
.B(n_1547),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1645),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1615),
.A2(n_1123),
.B1(n_1124),
.B2(n_1107),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1630),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1703),
.A2(n_1251),
.B1(n_1252),
.B2(n_1220),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1629),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1703),
.A2(n_1410),
.B1(n_1420),
.B2(n_1259),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1630),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1629),
.B(n_1082),
.Y(n_1948)
);

BUFx8_ASAP7_75t_L g1949 ( 
.A(n_1629),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1715),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1715),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1715),
.Y(n_1952)
);

INVx5_ASAP7_75t_L g1953 ( 
.A(n_1645),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1715),
.Y(n_1954)
);

INVx5_ASAP7_75t_L g1955 ( 
.A(n_1645),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1629),
.Y(n_1956)
);

CKINVDCx6p67_ASAP7_75t_R g1957 ( 
.A(n_1611),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1659),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1630),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1629),
.B(n_1130),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1715),
.Y(n_1961)
);

INVx6_ASAP7_75t_L g1962 ( 
.A(n_1645),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1826),
.B(n_1516),
.Y(n_1963)
);

CKINVDCx8_ASAP7_75t_R g1964 ( 
.A(n_1832),
.Y(n_1964)
);

AOI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1799),
.A2(n_1851),
.B1(n_1845),
.B2(n_1837),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1865),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1851),
.B(n_1516),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1865),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1853),
.B(n_1144),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1740),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1782),
.Y(n_1971)
);

BUFx8_ASAP7_75t_L g1972 ( 
.A(n_1834),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1740),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1841),
.B(n_1216),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1799),
.B(n_1089),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1852),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1863),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1871),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1796),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1805),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1885),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1885),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1784),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_1840),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1791),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1818),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1857),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1748),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1748),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1858),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1826),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1811),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1760),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1860),
.B(n_1269),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1831),
.B(n_1873),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1753),
.Y(n_1996)
);

INVx4_ASAP7_75t_L g1997 ( 
.A(n_1807),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1753),
.B(n_1047),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1893),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1788),
.Y(n_2000)
);

OAI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1895),
.A2(n_1477),
.B(n_1475),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1788),
.Y(n_2002)
);

AND2x6_ASAP7_75t_L g2003 ( 
.A(n_1881),
.B(n_1890),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1881),
.B(n_1047),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1890),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1772),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1744),
.Y(n_2007)
);

OA21x2_ASAP7_75t_L g2008 ( 
.A1(n_1750),
.A2(n_1488),
.B(n_1481),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1914),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1833),
.B(n_1406),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1914),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1838),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1893),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1777),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1816),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1905),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1900),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1783),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1745),
.B(n_1131),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1933),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1802),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1814),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1786),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1815),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_SL g2025 ( 
.A1(n_1823),
.A2(n_1911),
.B1(n_1946),
.B2(n_1944),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1819),
.B(n_1560),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1905),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1886),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1822),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1824),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1807),
.B(n_1089),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1821),
.B(n_1047),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1778),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1768),
.B(n_1141),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1785),
.B(n_1560),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1778),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1758),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1759),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1764),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1770),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1787),
.B(n_1769),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1922),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_1935),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1737),
.B(n_1142),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_1945),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1738),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1907),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1742),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1866),
.A2(n_1869),
.B1(n_1755),
.B2(n_1894),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1743),
.B(n_1151),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1746),
.B(n_1153),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1956),
.B(n_1093),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1747),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1907),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_1752),
.Y(n_2055)
);

INVx4_ASAP7_75t_L g2056 ( 
.A(n_1880),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1761),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1767),
.B(n_1775),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1874),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1916),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1766),
.B(n_1093),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1878),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_1916),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1793),
.Y(n_2064)
);

BUFx6f_ASAP7_75t_L g2065 ( 
.A(n_1917),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1884),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1896),
.Y(n_2067)
);

INVxp67_ASAP7_75t_L g2068 ( 
.A(n_1938),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_1917),
.Y(n_2069)
);

HB1xp67_ASAP7_75t_L g2070 ( 
.A(n_1864),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1908),
.B(n_1157),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1910),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1793),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1942),
.B(n_1160),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1915),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1912),
.B(n_1164),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1801),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1749),
.B(n_1093),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1736),
.B(n_1196),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1920),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1937),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1777),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1928),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1928),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_1804),
.Y(n_2085)
);

INVxp67_ASAP7_75t_L g2086 ( 
.A(n_1765),
.Y(n_2086)
);

AND2x6_ASAP7_75t_L g2087 ( 
.A(n_1943),
.B(n_1003),
.Y(n_2087)
);

OAI21x1_ASAP7_75t_L g2088 ( 
.A1(n_1830),
.A2(n_1517),
.B(n_1511),
.Y(n_2088)
);

BUFx3_ASAP7_75t_L g2089 ( 
.A(n_1929),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1947),
.B(n_1168),
.Y(n_2090)
);

AND2x6_ASAP7_75t_L g2091 ( 
.A(n_1959),
.B(n_1003),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1801),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1957),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1754),
.B(n_1169),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1806),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1929),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_SL g2097 ( 
.A(n_1797),
.B(n_1179),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1806),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_1889),
.B(n_1182),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1808),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1808),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1812),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1812),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_1776),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1817),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1817),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1829),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1829),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1844),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1844),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1930),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1856),
.Y(n_2112)
);

INVxp67_ASAP7_75t_L g2113 ( 
.A(n_1934),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1949),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1856),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1930),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_SL g2117 ( 
.A(n_1751),
.B(n_1185),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1859),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1859),
.Y(n_2119)
);

INVx3_ASAP7_75t_L g2120 ( 
.A(n_1936),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_1912),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1877),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1879),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_1739),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1790),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1794),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1936),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1789),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1780),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1792),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1887),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1898),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1883),
.B(n_1196),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1800),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1835),
.B(n_1187),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_1957),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1809),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1813),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1827),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_1951),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1904),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1888),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1836),
.Y(n_2143)
);

BUFx6f_ASAP7_75t_L g2144 ( 
.A(n_1951),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1940),
.B(n_1196),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1781),
.B(n_1275),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1952),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1913),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1843),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1842),
.B(n_1197),
.Y(n_2150)
);

OAI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_1847),
.A2(n_1204),
.B1(n_1206),
.B2(n_1198),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1850),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_L g2153 ( 
.A(n_1952),
.Y(n_2153)
);

BUFx6f_ASAP7_75t_L g2154 ( 
.A(n_1880),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1892),
.B(n_1275),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_1962),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1897),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1891),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_1897),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1919),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1924),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1868),
.B(n_1218),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_1875),
.Y(n_2163)
);

AND2x6_ASAP7_75t_L g2164 ( 
.A(n_1825),
.B(n_1903),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1862),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1867),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1921),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1876),
.B(n_1222),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1925),
.Y(n_2169)
);

CKINVDCx20_ASAP7_75t_R g2170 ( 
.A(n_1855),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1939),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1950),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1954),
.Y(n_2173)
);

BUFx8_ASAP7_75t_L g2174 ( 
.A(n_1906),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1961),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1924),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1741),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_1810),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1849),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1854),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1899),
.B(n_1226),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_1953),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1861),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_1902),
.Y(n_2184)
);

CKINVDCx8_ASAP7_75t_R g2185 ( 
.A(n_1762),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1846),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1872),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1872),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1803),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1741),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1820),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_1909),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_1923),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1926),
.B(n_1275),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_1927),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_1931),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1948),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1870),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_SL g2199 ( 
.A1(n_1757),
.A2(n_1023),
.B1(n_1284),
.B2(n_1024),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1960),
.B(n_1229),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_1739),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1763),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1870),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1953),
.B(n_1231),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1739),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1763),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1932),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1771),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_1941),
.B(n_1236),
.Y(n_2209)
);

INVx3_ASAP7_75t_L g2210 ( 
.A(n_1955),
.Y(n_2210)
);

INVxp67_ASAP7_75t_L g2211 ( 
.A(n_1828),
.Y(n_2211)
);

XNOR2xp5_ASAP7_75t_L g2212 ( 
.A(n_1882),
.B(n_1442),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1756),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1955),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_1779),
.Y(n_2215)
);

NAND2xp33_ASAP7_75t_SL g2216 ( 
.A(n_1918),
.B(n_1239),
.Y(n_2216)
);

INVx6_ASAP7_75t_L g2217 ( 
.A(n_1795),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1771),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1839),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1773),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1773),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1848),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1774),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1848),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1774),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1798),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1958),
.Y(n_2227)
);

OA21x2_ASAP7_75t_L g2228 ( 
.A1(n_1901),
.A2(n_1529),
.B(n_1527),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_1745),
.B(n_1243),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1865),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1865),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1871),
.Y(n_2232)
);

BUFx2_ASAP7_75t_L g2233 ( 
.A(n_1865),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1865),
.Y(n_2234)
);

AND2x6_ASAP7_75t_L g2235 ( 
.A(n_1851),
.B(n_1003),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_1840),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1865),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1871),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1865),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1865),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1837),
.B(n_1244),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1871),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_1799),
.B(n_1102),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_1840),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_1826),
.B(n_1383),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1871),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1871),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1865),
.Y(n_2248)
);

CKINVDCx8_ASAP7_75t_R g2249 ( 
.A(n_1832),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1865),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1865),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_1837),
.B(n_1245),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1865),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_1840),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1865),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1871),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_1865),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1826),
.B(n_1383),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_1865),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1871),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1865),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1865),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_1840),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1871),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1871),
.Y(n_2265)
);

OA21x2_ASAP7_75t_L g2266 ( 
.A1(n_1871),
.A2(n_1531),
.B(n_1530),
.Y(n_2266)
);

INVx5_ASAP7_75t_L g2267 ( 
.A(n_1968),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1986),
.B(n_1253),
.Y(n_2268)
);

BUFx3_ASAP7_75t_L g2269 ( 
.A(n_1972),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2017),
.B(n_1544),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_1968),
.B(n_1258),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1992),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2001),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_2259),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2042),
.Y(n_2275)
);

INVx3_ASAP7_75t_L g2276 ( 
.A(n_2259),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1979),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2192),
.B(n_1262),
.Y(n_2278)
);

INVx2_ASAP7_75t_SL g2279 ( 
.A(n_2020),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1979),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_2154),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2003),
.A2(n_1500),
.B1(n_1574),
.B2(n_1571),
.Y(n_2282)
);

INVx4_ASAP7_75t_L g2283 ( 
.A(n_2154),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1980),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2196),
.B(n_1273),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_1972),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1980),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_2157),
.Y(n_2288)
);

AND2x6_ASAP7_75t_L g2289 ( 
.A(n_1966),
.B(n_1003),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2018),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2021),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2023),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2003),
.B(n_1274),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2022),
.Y(n_2294)
);

BUFx3_ASAP7_75t_L g2295 ( 
.A(n_2114),
.Y(n_2295)
);

INVx4_ASAP7_75t_L g2296 ( 
.A(n_2157),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2240),
.B(n_2257),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2003),
.B(n_1277),
.Y(n_2298)
);

BUFx3_ASAP7_75t_L g2299 ( 
.A(n_2114),
.Y(n_2299)
);

BUFx4f_ASAP7_75t_L g2300 ( 
.A(n_2215),
.Y(n_2300)
);

INVx5_ASAP7_75t_L g2301 ( 
.A(n_2233),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2262),
.B(n_1282),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2233),
.B(n_1286),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2024),
.Y(n_2304)
);

BUFx10_ASAP7_75t_L g2305 ( 
.A(n_2217),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2029),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1963),
.B(n_1289),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2030),
.Y(n_2308)
);

NAND2x1_ASAP7_75t_L g2309 ( 
.A(n_2266),
.B(n_1125),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2128),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1988),
.B(n_1290),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2230),
.B(n_1292),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2008),
.Y(n_2313)
);

AOI22xp33_ASAP7_75t_L g2314 ( 
.A1(n_2198),
.A2(n_1579),
.B1(n_1326),
.B2(n_1461),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2231),
.B(n_2234),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2008),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2237),
.B(n_1293),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_2174),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2046),
.Y(n_2319)
);

BUFx2_ASAP7_75t_L g2320 ( 
.A(n_1984),
.Y(n_2320)
);

INVx4_ASAP7_75t_L g2321 ( 
.A(n_2161),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_2239),
.B(n_1237),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1989),
.B(n_1302),
.Y(n_2323)
);

AOI22xp33_ASAP7_75t_L g2324 ( 
.A1(n_2203),
.A2(n_1326),
.B1(n_1461),
.B2(n_1102),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2048),
.Y(n_2325)
);

AOI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_1991),
.A2(n_1312),
.B1(n_1317),
.B2(n_1305),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2053),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_1996),
.B(n_1323),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_1978),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2000),
.B(n_1332),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2015),
.B(n_1023),
.Y(n_2331)
);

OR2x6_ASAP7_75t_L g2332 ( 
.A(n_2217),
.B(n_1133),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2059),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_2161),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2244),
.B(n_1185),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2002),
.B(n_1336),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2232),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2055),
.B(n_1024),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2238),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_2174),
.Y(n_2340)
);

AOI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2005),
.A2(n_1542),
.B1(n_1552),
.B2(n_1537),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2236),
.B(n_1284),
.Y(n_2342)
);

AND2x4_ASAP7_75t_L g2343 ( 
.A(n_2248),
.B(n_999),
.Y(n_2343)
);

BUFx10_ASAP7_75t_L g2344 ( 
.A(n_2215),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2062),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2242),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2250),
.B(n_2251),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2066),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2246),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_1990),
.B(n_1015),
.Y(n_2350)
);

OAI22xp33_ASAP7_75t_L g2351 ( 
.A1(n_2117),
.A2(n_1366),
.B1(n_1066),
.B2(n_1075),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_2176),
.Y(n_2352)
);

OR2x2_ASAP7_75t_L g2353 ( 
.A(n_2254),
.B(n_1081),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2067),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2009),
.B(n_1343),
.Y(n_2355)
);

INVx4_ASAP7_75t_SL g2356 ( 
.A(n_2235),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2247),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2072),
.Y(n_2358)
);

XNOR2xp5_ASAP7_75t_L g2359 ( 
.A(n_2199),
.B(n_1366),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2011),
.B(n_1347),
.Y(n_2360)
);

NAND2xp33_ASAP7_75t_SL g2361 ( 
.A(n_2253),
.B(n_1017),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2256),
.Y(n_2362)
);

INVxp33_ASAP7_75t_SL g2363 ( 
.A(n_2212),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2075),
.Y(n_2364)
);

INVx1_ASAP7_75t_SL g2365 ( 
.A(n_2020),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2176),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2260),
.Y(n_2367)
);

INVx4_ASAP7_75t_L g2368 ( 
.A(n_2182),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_2182),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2265),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2080),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2255),
.B(n_1358),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2081),
.Y(n_2373)
);

INVx5_ASAP7_75t_L g2374 ( 
.A(n_2087),
.Y(n_2374)
);

CKINVDCx6p67_ASAP7_75t_R g2375 ( 
.A(n_2136),
.Y(n_2375)
);

INVx1_ASAP7_75t_SL g2376 ( 
.A(n_2043),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2178),
.Y(n_2377)
);

INVx1_ASAP7_75t_SL g2378 ( 
.A(n_2043),
.Y(n_2378)
);

AOI22xp33_ASAP7_75t_L g2379 ( 
.A1(n_1987),
.A2(n_1542),
.B1(n_1552),
.B2(n_1537),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2125),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_1965),
.B(n_2163),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2245),
.A2(n_1373),
.B1(n_1375),
.B2(n_1365),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2184),
.B(n_1379),
.Y(n_2383)
);

INVx4_ASAP7_75t_L g2384 ( 
.A(n_2214),
.Y(n_2384)
);

AND2x6_ASAP7_75t_L g2385 ( 
.A(n_2261),
.B(n_1125),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2126),
.Y(n_2386)
);

AND2x2_ASAP7_75t_SL g2387 ( 
.A(n_2070),
.B(n_1301),
.Y(n_2387)
);

CKINVDCx20_ASAP7_75t_R g2388 ( 
.A(n_2185),
.Y(n_2388)
);

INVx6_ASAP7_75t_L g2389 ( 
.A(n_2214),
.Y(n_2389)
);

INVx1_ASAP7_75t_SL g2390 ( 
.A(n_2263),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2193),
.B(n_1385),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2058),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1971),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1983),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2258),
.A2(n_2049),
.B1(n_1998),
.B2(n_2004),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_2121),
.B(n_1301),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1985),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_1969),
.B(n_1392),
.Y(n_2398)
);

OR2x2_ASAP7_75t_SL g2399 ( 
.A(n_2085),
.B(n_1595),
.Y(n_2399)
);

BUFx10_ASAP7_75t_L g2400 ( 
.A(n_2014),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2056),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2028),
.B(n_1383),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2057),
.B(n_1087),
.Y(n_2403)
);

CKINVDCx16_ASAP7_75t_R g2404 ( 
.A(n_2212),
.Y(n_2404)
);

BUFx10_ASAP7_75t_L g2405 ( 
.A(n_2082),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2068),
.B(n_1421),
.Y(n_2406)
);

BUFx10_ASAP7_75t_L g2407 ( 
.A(n_2093),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2142),
.A2(n_1396),
.B1(n_1405),
.B2(n_1393),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2266),
.Y(n_2409)
);

NAND2xp33_ASAP7_75t_L g2410 ( 
.A(n_2235),
.B(n_1426),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2130),
.Y(n_2411)
);

INVx8_ASAP7_75t_L g2412 ( 
.A(n_2235),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_1975),
.B(n_2243),
.Y(n_2413)
);

BUFx3_ASAP7_75t_L g2414 ( 
.A(n_2089),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2264),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2045),
.B(n_1173),
.Y(n_2416)
);

INVx4_ASAP7_75t_L g2417 ( 
.A(n_1997),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_1975),
.B(n_1589),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2134),
.Y(n_2419)
);

HB1xp67_ASAP7_75t_L g2420 ( 
.A(n_2104),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2052),
.B(n_2079),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2243),
.B(n_1592),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2137),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2135),
.B(n_1593),
.Y(n_2424)
);

HB1xp67_ASAP7_75t_L g2425 ( 
.A(n_2151),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2138),
.Y(n_2426)
);

INVx1_ASAP7_75t_SL g2427 ( 
.A(n_2031),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2150),
.B(n_1597),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2159),
.Y(n_2429)
);

AND2x4_ASAP7_75t_L g2430 ( 
.A(n_2186),
.B(n_1008),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2264),
.Y(n_2431)
);

INVx3_ASAP7_75t_L g2432 ( 
.A(n_1970),
.Y(n_2432)
);

INVx4_ASAP7_75t_L g2433 ( 
.A(n_1976),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2162),
.B(n_1598),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2010),
.B(n_1599),
.Y(n_2435)
);

AND3x2_ASAP7_75t_L g2436 ( 
.A(n_2086),
.B(n_1595),
.C(n_1424),
.Y(n_2436)
);

AO22x2_ASAP7_75t_L g2437 ( 
.A1(n_2211),
.A2(n_2183),
.B1(n_2155),
.B2(n_2025),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2006),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2139),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_1977),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_2156),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2074),
.A2(n_1417),
.B1(n_1423),
.B2(n_1416),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2143),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_1970),
.Y(n_2444)
);

OAI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_1964),
.A2(n_1176),
.B1(n_1460),
.B2(n_1446),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2149),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2097),
.B(n_1469),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2152),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2146),
.B(n_1532),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2168),
.B(n_1584),
.Y(n_2450)
);

NAND2xp33_ASAP7_75t_SL g2451 ( 
.A(n_2124),
.B(n_1580),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2165),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2124),
.B(n_1600),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2181),
.B(n_1427),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_SL g2455 ( 
.A(n_1995),
.B(n_1472),
.Y(n_2455)
);

OR2x2_ASAP7_75t_L g2456 ( 
.A(n_2032),
.B(n_1591),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2166),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2037),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2200),
.B(n_1501),
.Y(n_2459)
);

INVx3_ASAP7_75t_L g2460 ( 
.A(n_1973),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2007),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_1974),
.B(n_1513),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2061),
.B(n_1429),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2122),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_2113),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2038),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_2249),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2123),
.Y(n_2468)
);

INVx3_ASAP7_75t_L g2469 ( 
.A(n_1973),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2133),
.B(n_1430),
.Y(n_2470)
);

BUFx4f_ASAP7_75t_L g2471 ( 
.A(n_2226),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_1994),
.B(n_1479),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2041),
.B(n_1433),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2039),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_1999),
.Y(n_2475)
);

NAND2xp33_ASAP7_75t_L g2476 ( 
.A(n_2087),
.B(n_1443),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2145),
.B(n_1444),
.Y(n_2477)
);

INVx6_ASAP7_75t_L g2478 ( 
.A(n_1999),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_SL g2479 ( 
.A(n_2164),
.Y(n_2479)
);

BUFx4f_ASAP7_75t_L g2480 ( 
.A(n_2164),
.Y(n_2480)
);

BUFx2_ASAP7_75t_L g2481 ( 
.A(n_2087),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2076),
.B(n_1445),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_2241),
.B(n_1448),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2252),
.B(n_1454),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2047),
.Y(n_2485)
);

INVx1_ASAP7_75t_SL g2486 ( 
.A(n_2031),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_SL g2487 ( 
.A(n_2201),
.B(n_2044),
.Y(n_2487)
);

INVxp33_ASAP7_75t_L g2488 ( 
.A(n_2078),
.Y(n_2488)
);

XOR2xp5_ASAP7_75t_L g2489 ( 
.A(n_2170),
.B(n_1455),
.Y(n_2489)
);

INVx4_ASAP7_75t_L g2490 ( 
.A(n_2047),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2050),
.B(n_1466),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2040),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_2091),
.Y(n_2493)
);

BUFx3_ASAP7_75t_L g2494 ( 
.A(n_2060),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2194),
.B(n_1489),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2131),
.Y(n_2496)
);

AND2x6_ASAP7_75t_L g2497 ( 
.A(n_2205),
.B(n_1125),
.Y(n_2497)
);

OR2x6_ASAP7_75t_L g2498 ( 
.A(n_2227),
.B(n_1126),
.Y(n_2498)
);

AND2x6_ASAP7_75t_L g2499 ( 
.A(n_2012),
.B(n_1125),
.Y(n_2499)
);

INVx2_ASAP7_75t_SL g2500 ( 
.A(n_2060),
.Y(n_2500)
);

OR2x2_ASAP7_75t_L g2501 ( 
.A(n_2216),
.B(n_1162),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2019),
.B(n_1492),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_L g2503 ( 
.A(n_1967),
.B(n_2197),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2034),
.B(n_1494),
.Y(n_2504)
);

BUFx6f_ASAP7_75t_L g2505 ( 
.A(n_2065),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2051),
.B(n_1496),
.Y(n_2506)
);

INVx4_ASAP7_75t_L g2507 ( 
.A(n_2065),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2035),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2132),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2179),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_L g2511 ( 
.A(n_2094),
.B(n_1503),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2083),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2180),
.Y(n_2513)
);

BUFx6f_ASAP7_75t_L g2514 ( 
.A(n_2083),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2071),
.B(n_1512),
.Y(n_2515)
);

NAND3xp33_ASAP7_75t_L g2516 ( 
.A(n_2099),
.B(n_1533),
.C(n_1518),
.Y(n_2516)
);

AND2x4_ASAP7_75t_L g2517 ( 
.A(n_2222),
.B(n_1011),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2141),
.Y(n_2518)
);

HB1xp67_ASAP7_75t_L g2519 ( 
.A(n_2228),
.Y(n_2519)
);

AOI22xp33_ASAP7_75t_L g2520 ( 
.A1(n_2090),
.A2(n_1546),
.B1(n_1550),
.B2(n_1545),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2209),
.B(n_2229),
.Y(n_2521)
);

BUFx2_ASAP7_75t_L g2522 ( 
.A(n_2091),
.Y(n_2522)
);

INVx2_ASAP7_75t_SL g2523 ( 
.A(n_2096),
.Y(n_2523)
);

INVx5_ASAP7_75t_L g2524 ( 
.A(n_2091),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2167),
.Y(n_2525)
);

INVxp67_ASAP7_75t_SL g2526 ( 
.A(n_2210),
.Y(n_2526)
);

OR2x2_ASAP7_75t_L g2527 ( 
.A(n_2204),
.B(n_1356),
.Y(n_2527)
);

AND2x2_ASAP7_75t_SL g2528 ( 
.A(n_2228),
.B(n_1586),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_SL g2529 ( 
.A(n_2164),
.B(n_1553),
.Y(n_2529)
);

BUFx10_ASAP7_75t_L g2530 ( 
.A(n_2096),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2148),
.Y(n_2531)
);

OAI22xp33_ASAP7_75t_L g2532 ( 
.A1(n_2189),
.A2(n_1555),
.B1(n_1566),
.B2(n_1380),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2160),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2169),
.Y(n_2534)
);

INVx4_ASAP7_75t_L g2535 ( 
.A(n_2111),
.Y(n_2535)
);

INVx4_ASAP7_75t_L g2536 ( 
.A(n_2111),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_2129),
.B(n_1002),
.Y(n_2537)
);

AND2x2_ASAP7_75t_SL g2538 ( 
.A(n_2116),
.B(n_1540),
.Y(n_2538)
);

INVxp67_ASAP7_75t_SL g2539 ( 
.A(n_2116),
.Y(n_2539)
);

OAI22xp33_ASAP7_75t_L g2540 ( 
.A1(n_2191),
.A2(n_1601),
.B1(n_1005),
.B2(n_1028),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_1993),
.Y(n_2541)
);

AND2x6_ASAP7_75t_L g2542 ( 
.A(n_2224),
.B(n_1401),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2158),
.Y(n_2543)
);

INVxp67_ASAP7_75t_L g2544 ( 
.A(n_2195),
.Y(n_2544)
);

OR2x6_ASAP7_75t_L g2545 ( 
.A(n_2207),
.B(n_1177),
.Y(n_2545)
);

BUFx3_ASAP7_75t_L g2546 ( 
.A(n_2127),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2171),
.Y(n_2547)
);

BUFx8_ASAP7_75t_SL g2548 ( 
.A(n_2127),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2026),
.A2(n_1021),
.B1(n_1039),
.B2(n_1031),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2172),
.B(n_2173),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2175),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2144),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2213),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2187),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2188),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2115),
.B(n_1581),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2144),
.Y(n_2557)
);

INVx3_ASAP7_75t_L g2558 ( 
.A(n_2153),
.Y(n_2558)
);

OR2x2_ASAP7_75t_L g2559 ( 
.A(n_1981),
.B(n_990),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2153),
.B(n_1159),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2115),
.B(n_1587),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2036),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2219),
.B(n_1543),
.Y(n_2563)
);

AOI22xp33_ASAP7_75t_L g2564 ( 
.A1(n_2095),
.A2(n_1549),
.B1(n_1563),
.B2(n_1554),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_1982),
.B(n_1564),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_L g2566 ( 
.A(n_2013),
.B(n_1043),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2098),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2088),
.Y(n_2568)
);

NAND2xp33_ASAP7_75t_SL g2569 ( 
.A(n_2103),
.B(n_1055),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2106),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2016),
.B(n_1295),
.Y(n_2571)
);

NAND2x1p5_ASAP7_75t_L g2572 ( 
.A(n_2027),
.B(n_1327),
.Y(n_2572)
);

BUFx3_ASAP7_75t_L g2573 ( 
.A(n_2054),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2064),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2107),
.Y(n_2575)
);

AND2x2_ASAP7_75t_SL g2576 ( 
.A(n_2063),
.B(n_1101),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2073),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_L g2578 ( 
.A(n_2069),
.B(n_1056),
.Y(n_2578)
);

OA22x2_ASAP7_75t_L g2579 ( 
.A1(n_2084),
.A2(n_1063),
.B1(n_1064),
.B2(n_1060),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2112),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2077),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2092),
.Y(n_2582)
);

OAI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2100),
.A2(n_1030),
.B1(n_1033),
.B2(n_1012),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2101),
.Y(n_2584)
);

INVx3_ASAP7_75t_L g2585 ( 
.A(n_2120),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2102),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2140),
.Y(n_2587)
);

INVx4_ASAP7_75t_L g2588 ( 
.A(n_2147),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2105),
.A2(n_1401),
.B1(n_1042),
.B2(n_1046),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_2108),
.B(n_1067),
.Y(n_2590)
);

INVxp67_ASAP7_75t_L g2591 ( 
.A(n_2109),
.Y(n_2591)
);

CKINVDCx20_ASAP7_75t_R g2592 ( 
.A(n_2033),
.Y(n_2592)
);

INVxp67_ASAP7_75t_SL g2593 ( 
.A(n_2110),
.Y(n_2593)
);

NAND2xp33_ASAP7_75t_L g2594 ( 
.A(n_2118),
.B(n_1068),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2119),
.B(n_1071),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2225),
.B(n_1072),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2177),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2190),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2202),
.B(n_1074),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2206),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_SL g2601 ( 
.A(n_2208),
.B(n_1078),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2218),
.B(n_1086),
.Y(n_2602)
);

INVxp67_ASAP7_75t_L g2603 ( 
.A(n_2223),
.Y(n_2603)
);

HB1xp67_ASAP7_75t_L g2604 ( 
.A(n_2220),
.Y(n_2604)
);

OAI22xp5_ASAP7_75t_L g2605 ( 
.A1(n_2221),
.A2(n_1062),
.B1(n_1065),
.B2(n_1034),
.Y(n_2605)
);

INVx4_ASAP7_75t_SL g2606 ( 
.A(n_1968),
.Y(n_2606)
);

BUFx8_ASAP7_75t_SL g2607 ( 
.A(n_2114),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_1992),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_1986),
.B(n_1095),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_1986),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_1968),
.B(n_1099),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1986),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_1991),
.B(n_1100),
.Y(n_2613)
);

AND2x4_ASAP7_75t_L g2614 ( 
.A(n_2233),
.B(n_1076),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_1991),
.B(n_1105),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_1991),
.B(n_1108),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_2003),
.A2(n_1401),
.B1(n_1098),
.B2(n_1114),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_1968),
.Y(n_2618)
);

INVx2_ASAP7_75t_SL g2619 ( 
.A(n_1968),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_1986),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_1986),
.Y(n_2621)
);

BUFx3_ASAP7_75t_L g2622 ( 
.A(n_1972),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_1972),
.Y(n_2623)
);

NAND3xp33_ASAP7_75t_SL g2624 ( 
.A(n_2055),
.B(n_1486),
.C(n_1465),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1986),
.Y(n_2625)
);

HB1xp67_ASAP7_75t_L g2626 ( 
.A(n_1984),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_1991),
.B(n_1110),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_SL g2628 ( 
.A(n_1968),
.B(n_1109),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_1992),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_1992),
.Y(n_2630)
);

INVx6_ASAP7_75t_L g2631 ( 
.A(n_1972),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_1991),
.B(n_1113),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_1986),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_1986),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_1992),
.Y(n_2635)
);

OR2x2_ASAP7_75t_L g2636 ( 
.A(n_2055),
.B(n_1499),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_1986),
.B(n_1111),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_1986),
.B(n_1117),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_1968),
.B(n_1118),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2003),
.A2(n_1401),
.B1(n_1128),
.B2(n_1136),
.Y(n_2640)
);

BUFx4f_ASAP7_75t_L g2641 ( 
.A(n_2215),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_1992),
.Y(n_2642)
);

INVx4_ASAP7_75t_L g2643 ( 
.A(n_1968),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2233),
.B(n_1077),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_1968),
.Y(n_2645)
);

BUFx4f_ASAP7_75t_L g2646 ( 
.A(n_2215),
.Y(n_2646)
);

INVx1_ASAP7_75t_SL g2647 ( 
.A(n_2055),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_1972),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_SL g2649 ( 
.A(n_2647),
.B(n_1583),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2610),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2488),
.B(n_1120),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2392),
.B(n_1121),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2612),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2381),
.A2(n_1127),
.B1(n_1134),
.B2(n_1122),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2620),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_2444),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2621),
.Y(n_2657)
);

O2A1O1Ixp33_ASAP7_75t_L g2658 ( 
.A1(n_2521),
.A2(n_1577),
.B(n_1567),
.C(n_1139),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2625),
.Y(n_2659)
);

NAND3x1_ASAP7_75t_L g2660 ( 
.A(n_2338),
.B(n_1582),
.C(n_1568),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2633),
.B(n_1145),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_R g2662 ( 
.A(n_2623),
.B(n_1149),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2390),
.B(n_2529),
.Y(n_2663)
);

NOR3xp33_ASAP7_75t_L g2664 ( 
.A(n_2624),
.B(n_1590),
.C(n_1585),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2634),
.B(n_1154),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2320),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_SL g2667 ( 
.A(n_2412),
.B(n_1165),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2277),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2320),
.B(n_1576),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2280),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2270),
.B(n_1167),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2291),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2395),
.B(n_1171),
.Y(n_2673)
);

AOI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2437),
.A2(n_1175),
.B1(n_1184),
.B2(n_1174),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2284),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2294),
.B(n_1188),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2304),
.B(n_1189),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_SL g2678 ( 
.A(n_2538),
.B(n_1556),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2425),
.B(n_1190),
.Y(n_2679)
);

BUFx2_ASAP7_75t_L g2680 ( 
.A(n_2626),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2306),
.B(n_1191),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2449),
.B(n_1195),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2287),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2308),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2365),
.B(n_2376),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2437),
.A2(n_2421),
.B1(n_2528),
.B2(n_2477),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2495),
.B(n_1199),
.Y(n_2687)
);

A2O1A1Ixp33_ASAP7_75t_L g2688 ( 
.A1(n_2508),
.A2(n_1150),
.B(n_1152),
.C(n_1138),
.Y(n_2688)
);

NAND2x1p5_ASAP7_75t_L g2689 ( 
.A(n_2267),
.B(n_1119),
.Y(n_2689)
);

XNOR2xp5_ASAP7_75t_L g2690 ( 
.A(n_2332),
.B(n_2359),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2403),
.B(n_1201),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2331),
.B(n_1202),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2310),
.Y(n_2693)
);

NOR2xp67_ASAP7_75t_L g2694 ( 
.A(n_2648),
.B(n_1),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2378),
.B(n_1588),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2301),
.B(n_1156),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2380),
.B(n_1203),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2415),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2386),
.B(n_1205),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2319),
.B(n_1207),
.Y(n_2700)
);

BUFx6f_ASAP7_75t_L g2701 ( 
.A(n_2444),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2431),
.Y(n_2702)
);

NAND3x1_ASAP7_75t_L g2703 ( 
.A(n_2399),
.B(n_1594),
.C(n_1558),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_SL g2704 ( 
.A(n_2532),
.B(n_1539),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2342),
.B(n_1209),
.Y(n_2705)
);

A2O1A1Ixp33_ASAP7_75t_L g2706 ( 
.A1(n_2511),
.A2(n_1166),
.B(n_1180),
.C(n_1163),
.Y(n_2706)
);

INVx4_ASAP7_75t_L g2707 ( 
.A(n_2267),
.Y(n_2707)
);

AND2x6_ASAP7_75t_SL g2708 ( 
.A(n_2332),
.B(n_1192),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2313),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2470),
.B(n_1210),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2267),
.B(n_1569),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2325),
.B(n_1211),
.Y(n_2712)
);

NOR2x1p5_ASAP7_75t_L g2713 ( 
.A(n_2318),
.B(n_1215),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2340),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2327),
.B(n_2333),
.Y(n_2715)
);

NOR2xp67_ASAP7_75t_L g2716 ( 
.A(n_2269),
.B(n_1),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2345),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2348),
.B(n_2354),
.Y(n_2718)
);

AND2x4_ASAP7_75t_L g2719 ( 
.A(n_2301),
.B(n_1208),
.Y(n_2719)
);

AOI22xp33_ASAP7_75t_L g2720 ( 
.A1(n_2463),
.A2(n_1221),
.B1(n_1228),
.B2(n_1217),
.Y(n_2720)
);

INVx2_ASAP7_75t_SL g2721 ( 
.A(n_2344),
.Y(n_2721)
);

OAI221xp5_ASAP7_75t_L g2722 ( 
.A1(n_2282),
.A2(n_2408),
.B1(n_2382),
.B2(n_2456),
.C(n_2307),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_SL g2723 ( 
.A(n_2279),
.B(n_1535),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_SL g2724 ( 
.A(n_2301),
.B(n_1572),
.Y(n_2724)
);

INVxp67_ASAP7_75t_SL g2725 ( 
.A(n_2445),
.Y(n_2725)
);

INVx2_ASAP7_75t_SL g2726 ( 
.A(n_2344),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2358),
.B(n_1234),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2364),
.B(n_1235),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2353),
.B(n_1247),
.Y(n_2729)
);

NAND2xp33_ASAP7_75t_SL g2730 ( 
.A(n_2479),
.B(n_1254),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2416),
.B(n_1256),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2371),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2451),
.B(n_1559),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2373),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2393),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2383),
.B(n_2391),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2278),
.B(n_1257),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_L g2738 ( 
.A(n_2396),
.B(n_1263),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2316),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2268),
.B(n_1270),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2394),
.Y(n_2741)
);

INVxp33_ASAP7_75t_L g2742 ( 
.A(n_2350),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2275),
.A2(n_1281),
.B1(n_1287),
.B2(n_1280),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_SL g2744 ( 
.A(n_2361),
.B(n_1288),
.Y(n_2744)
);

A2O1A1Ixp33_ASAP7_75t_L g2745 ( 
.A1(n_2519),
.A2(n_1214),
.B(n_1219),
.C(n_1212),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2272),
.A2(n_1297),
.B1(n_1299),
.B2(n_1291),
.Y(n_2746)
);

BUFx10_ASAP7_75t_L g2747 ( 
.A(n_2631),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2281),
.B(n_1541),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2473),
.B(n_1303),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2281),
.B(n_1557),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2475),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2502),
.B(n_1304),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2285),
.B(n_1319),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2636),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2527),
.B(n_1328),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2290),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2491),
.B(n_1329),
.Y(n_2757)
);

NAND3xp33_ASAP7_75t_L g2758 ( 
.A(n_2324),
.B(n_1278),
.C(n_1119),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2402),
.B(n_1337),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2397),
.Y(n_2760)
);

NOR3xp33_ASAP7_75t_L g2761 ( 
.A(n_2351),
.B(n_1233),
.C(n_1224),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_L g2762 ( 
.A(n_2614),
.B(n_1340),
.Y(n_2762)
);

OAI22xp5_ASAP7_75t_SL g2763 ( 
.A1(n_2359),
.A2(n_1524),
.B1(n_1526),
.B2(n_1523),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2614),
.B(n_1345),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2411),
.Y(n_2765)
);

BUFx3_ASAP7_75t_L g2766 ( 
.A(n_2548),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2311),
.A2(n_1355),
.B1(n_1357),
.B2(n_1351),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2419),
.Y(n_2768)
);

BUFx6f_ASAP7_75t_L g2769 ( 
.A(n_2475),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2506),
.B(n_1364),
.Y(n_2770)
);

AOI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_2430),
.A2(n_1372),
.B1(n_1377),
.B2(n_1368),
.Y(n_2771)
);

NAND2xp33_ASAP7_75t_L g2772 ( 
.A(n_2412),
.B(n_1378),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_2420),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2423),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_2334),
.B(n_1382),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2426),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2439),
.Y(n_2777)
);

INVx2_ASAP7_75t_SL g2778 ( 
.A(n_2305),
.Y(n_2778)
);

INVx2_ASAP7_75t_SL g2779 ( 
.A(n_2305),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2430),
.A2(n_1388),
.B1(n_1389),
.B2(n_1386),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2443),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_2607),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2515),
.B(n_1391),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_SL g2784 ( 
.A(n_2334),
.B(n_1565),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2505),
.B(n_1575),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2292),
.Y(n_2786)
);

OR2x2_ASAP7_75t_L g2787 ( 
.A(n_2404),
.B(n_1394),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2446),
.Y(n_2788)
);

INVxp67_ASAP7_75t_L g2789 ( 
.A(n_2286),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2450),
.B(n_1395),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2448),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2295),
.Y(n_2792)
);

AOI22xp33_ASAP7_75t_L g2793 ( 
.A1(n_2322),
.A2(n_1399),
.B1(n_1400),
.B2(n_1397),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2622),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_L g2795 ( 
.A1(n_2322),
.A2(n_1413),
.B1(n_1414),
.B2(n_1411),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_SL g2796 ( 
.A(n_2374),
.B(n_1428),
.Y(n_2796)
);

AOI221xp5_ASAP7_75t_L g2797 ( 
.A1(n_2398),
.A2(n_1264),
.B1(n_1265),
.B2(n_1246),
.C(n_1240),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2323),
.A2(n_1434),
.B1(n_1435),
.B2(n_1431),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2328),
.A2(n_1449),
.B1(n_1450),
.B2(n_1440),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2452),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2644),
.B(n_1451),
.Y(n_2801)
);

AND2x6_ASAP7_75t_L g2802 ( 
.A(n_2505),
.B(n_1101),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_L g2803 ( 
.A(n_2644),
.B(n_1452),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_SL g2804 ( 
.A(n_2514),
.B(n_1456),
.Y(n_2804)
);

NAND3xp33_ASAP7_75t_L g2805 ( 
.A(n_2314),
.B(n_1278),
.C(n_1119),
.Y(n_2805)
);

AOI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2330),
.A2(n_1467),
.B1(n_1470),
.B2(n_1457),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2326),
.B(n_1473),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_SL g2808 ( 
.A(n_2374),
.B(n_1482),
.Y(n_2808)
);

AO221x1_ASAP7_75t_L g2809 ( 
.A1(n_2481),
.A2(n_1339),
.B1(n_1398),
.B2(n_1278),
.C(n_1119),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2514),
.Y(n_2810)
);

BUFx4_ASAP7_75t_L g2811 ( 
.A(n_2631),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2300),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2501),
.B(n_1484),
.Y(n_2813)
);

NAND2x1p5_ASAP7_75t_L g2814 ( 
.A(n_2643),
.B(n_1278),
.Y(n_2814)
);

NOR3xp33_ASAP7_75t_L g2815 ( 
.A(n_2335),
.B(n_1520),
.C(n_1515),
.Y(n_2815)
);

AOI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2336),
.A2(n_1490),
.B1(n_1493),
.B2(n_1485),
.Y(n_2816)
);

AOI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2355),
.A2(n_2360),
.B1(n_2343),
.B2(n_2517),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2613),
.B(n_1495),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2454),
.B(n_1510),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2424),
.B(n_1534),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2608),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2428),
.B(n_1562),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2434),
.B(n_1578),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2609),
.B(n_1267),
.Y(n_2824)
);

NOR2xp67_ASAP7_75t_L g2825 ( 
.A(n_2467),
.B(n_2),
.Y(n_2825)
);

AND2x2_ASAP7_75t_L g2826 ( 
.A(n_2615),
.B(n_1268),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2606),
.B(n_1279),
.Y(n_2827)
);

NOR2xp67_ASAP7_75t_L g2828 ( 
.A(n_2433),
.B(n_2),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2375),
.B(n_1294),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2637),
.B(n_1497),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2638),
.B(n_1505),
.Y(n_2831)
);

INVxp67_ASAP7_75t_L g2832 ( 
.A(n_2299),
.Y(n_2832)
);

INVx3_ASAP7_75t_L g2833 ( 
.A(n_2530),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2510),
.B(n_1506),
.Y(n_2834)
);

INVx2_ASAP7_75t_SL g2835 ( 
.A(n_2641),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2513),
.B(n_2435),
.Y(n_2836)
);

INVxp67_ASAP7_75t_SL g2837 ( 
.A(n_2410),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2457),
.Y(n_2838)
);

AND2x4_ASAP7_75t_L g2839 ( 
.A(n_2606),
.B(n_1300),
.Y(n_2839)
);

INVxp67_ASAP7_75t_L g2840 ( 
.A(n_2560),
.Y(n_2840)
);

INVx2_ASAP7_75t_SL g2841 ( 
.A(n_2646),
.Y(n_2841)
);

INVx2_ASAP7_75t_SL g2842 ( 
.A(n_2530),
.Y(n_2842)
);

OR2x6_ASAP7_75t_L g2843 ( 
.A(n_2572),
.B(n_1129),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2629),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2413),
.B(n_1508),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2520),
.B(n_1521),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2458),
.B(n_1536),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2630),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2466),
.B(n_1306),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2474),
.B(n_1307),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2635),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2492),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_SL g2853 ( 
.A(n_2576),
.B(n_1339),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2427),
.B(n_1313),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_SL g2855 ( 
.A(n_2540),
.B(n_1339),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2552),
.B(n_1339),
.Y(n_2856)
);

NAND3xp33_ASAP7_75t_L g2857 ( 
.A(n_2617),
.B(n_1403),
.C(n_1398),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2343),
.B(n_1314),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2616),
.B(n_1325),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2565),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2627),
.B(n_1330),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2480),
.B(n_1398),
.Y(n_2862)
);

INVx2_ASAP7_75t_SL g2863 ( 
.A(n_2389),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_2486),
.B(n_1419),
.Y(n_2864)
);

AOI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2517),
.A2(n_1335),
.B1(n_1344),
.B2(n_1331),
.Y(n_2865)
);

INVx2_ASAP7_75t_SL g2866 ( 
.A(n_2389),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2619),
.B(n_1398),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2632),
.B(n_1458),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2525),
.B(n_1459),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2303),
.B(n_1463),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2553),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2418),
.B(n_1349),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2534),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2547),
.B(n_2551),
.Y(n_2874)
);

INVx3_ASAP7_75t_R g2875 ( 
.A(n_2465),
.Y(n_2875)
);

NAND2xp33_ASAP7_75t_L g2876 ( 
.A(n_2289),
.B(n_1403),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2504),
.B(n_1350),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2550),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2642),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2482),
.B(n_1353),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2579),
.A2(n_1363),
.B1(n_1374),
.B2(n_1354),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_L g2882 ( 
.A1(n_2422),
.A2(n_1381),
.B1(n_1387),
.B2(n_1376),
.Y(n_2882)
);

AOI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2273),
.A2(n_1404),
.B(n_1390),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2442),
.B(n_1418),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2563),
.B(n_2459),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2329),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2556),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2561),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2464),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2337),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2339),
.Y(n_2891)
);

BUFx6f_ASAP7_75t_L g2892 ( 
.A(n_2374),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2498),
.B(n_1425),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2483),
.B(n_1437),
.Y(n_2894)
);

INVx2_ASAP7_75t_SL g2895 ( 
.A(n_2471),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2484),
.B(n_2503),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2468),
.Y(n_2897)
);

INVx4_ASAP7_75t_L g2898 ( 
.A(n_2478),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_2645),
.B(n_1403),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2496),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2564),
.B(n_1438),
.Y(n_2901)
);

NOR3xp33_ASAP7_75t_L g2902 ( 
.A(n_2516),
.B(n_1453),
.C(n_1415),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2509),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2640),
.B(n_1408),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2293),
.B(n_1129),
.Y(n_2905)
);

HB1xp67_ASAP7_75t_L g2906 ( 
.A(n_2440),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2298),
.B(n_1146),
.Y(n_2907)
);

HB1xp67_ASAP7_75t_L g2908 ( 
.A(n_2498),
.Y(n_2908)
);

AND2x4_ASAP7_75t_L g2909 ( 
.A(n_2315),
.B(n_1146),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2518),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2543),
.B(n_1403),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2462),
.B(n_1148),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2531),
.Y(n_2913)
);

NOR3xp33_ASAP7_75t_L g2914 ( 
.A(n_2447),
.B(n_1194),
.C(n_1148),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2533),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_SL g2916 ( 
.A(n_2524),
.B(n_1194),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2472),
.B(n_2549),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_SL g2918 ( 
.A(n_2524),
.B(n_1238),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2455),
.B(n_1238),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2481),
.B(n_1538),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2346),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2349),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2341),
.B(n_1255),
.Y(n_2923)
);

INVx8_ASAP7_75t_L g2924 ( 
.A(n_2289),
.Y(n_2924)
);

AND2x4_ASAP7_75t_L g2925 ( 
.A(n_2347),
.B(n_2554),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2438),
.A2(n_2461),
.B1(n_2409),
.B2(n_2362),
.Y(n_2926)
);

INVx4_ASAP7_75t_L g2927 ( 
.A(n_2478),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2357),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2312),
.B(n_1255),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2493),
.B(n_1538),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2367),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2317),
.B(n_1360),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_SL g2933 ( 
.A1(n_2363),
.A2(n_1402),
.B1(n_1468),
.B2(n_1360),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2571),
.B(n_1402),
.Y(n_2934)
);

INVx3_ASAP7_75t_L g2935 ( 
.A(n_2494),
.Y(n_2935)
);

NOR2xp67_ASAP7_75t_L g2936 ( 
.A(n_2377),
.B(n_2),
.Y(n_2936)
);

INVx8_ASAP7_75t_L g2937 ( 
.A(n_2289),
.Y(n_2937)
);

INVxp67_ASAP7_75t_L g2938 ( 
.A(n_2559),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_2400),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2370),
.A2(n_1474),
.B1(n_1502),
.B2(n_1468),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2583),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_SL g2942 ( 
.A(n_2524),
.B(n_1474),
.Y(n_2942)
);

INVx2_ASAP7_75t_SL g2943 ( 
.A(n_2400),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2372),
.B(n_1502),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2302),
.B(n_1509),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2379),
.B(n_2555),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2406),
.B(n_1509),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2274),
.B(n_1596),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2545),
.B(n_1596),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2276),
.B(n_3),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2541),
.Y(n_2951)
);

OAI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2592),
.A2(n_1551),
.B1(n_1538),
.B2(n_5),
.Y(n_2952)
);

OR2x2_ASAP7_75t_L g2953 ( 
.A(n_2283),
.B(n_3),
.Y(n_2953)
);

AOI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2605),
.A2(n_1551),
.B1(n_1538),
.B2(n_6),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2618),
.B(n_3),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2537),
.B(n_4),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2487),
.B(n_4),
.Y(n_2957)
);

INVxp67_ASAP7_75t_L g2958 ( 
.A(n_2545),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2562),
.Y(n_2959)
);

AOI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2569),
.A2(n_1551),
.B1(n_7),
.B2(n_4),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_2493),
.B(n_1551),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2522),
.B(n_7),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2567),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2453),
.B(n_6),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2544),
.B(n_6),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2296),
.B(n_8),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2522),
.B(n_9),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2570),
.Y(n_2968)
);

INVx8_ASAP7_75t_L g2969 ( 
.A(n_2385),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2356),
.B(n_10),
.Y(n_2970)
);

NOR3xp33_ASAP7_75t_L g2971 ( 
.A(n_2271),
.B(n_11),
.C(n_10),
.Y(n_2971)
);

INVxp67_ASAP7_75t_L g2972 ( 
.A(n_2546),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2526),
.B(n_8),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2441),
.B(n_2401),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_SL g2975 ( 
.A(n_2356),
.B(n_11),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2575),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2580),
.Y(n_2977)
);

INVx2_ASAP7_75t_SL g2978 ( 
.A(n_2405),
.Y(n_2978)
);

NAND2xp33_ASAP7_75t_L g2979 ( 
.A(n_2385),
.B(n_12),
.Y(n_2979)
);

INVxp67_ASAP7_75t_L g2980 ( 
.A(n_2557),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2321),
.B(n_10),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2429),
.B(n_12),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2596),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2599),
.B(n_2602),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2500),
.B(n_12),
.Y(n_2985)
);

OR2x2_ASAP7_75t_L g2986 ( 
.A(n_2368),
.B(n_13),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2568),
.Y(n_2987)
);

INVxp67_ASAP7_75t_L g2988 ( 
.A(n_2566),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2523),
.B(n_2578),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2384),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2288),
.B(n_13),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2574),
.Y(n_2992)
);

O2A1O1Ixp33_ASAP7_75t_L g2993 ( 
.A1(n_2594),
.A2(n_2628),
.B(n_2639),
.C(n_2611),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2352),
.B(n_14),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2297),
.B(n_14),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2366),
.B(n_15),
.Y(n_2996)
);

NOR3xp33_ASAP7_75t_L g2997 ( 
.A(n_2590),
.B(n_17),
.C(n_16),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2369),
.B(n_15),
.Y(n_2998)
);

NAND2xp33_ASAP7_75t_SL g2999 ( 
.A(n_2388),
.B(n_16),
.Y(n_2999)
);

AOI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2589),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2577),
.Y(n_3001)
);

INVx2_ASAP7_75t_SL g3002 ( 
.A(n_2405),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2604),
.Y(n_3003)
);

AND2x6_ASAP7_75t_SL g3004 ( 
.A(n_2489),
.B(n_18),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2490),
.B(n_18),
.Y(n_3005)
);

INVx3_ASAP7_75t_L g3006 ( 
.A(n_2507),
.Y(n_3006)
);

NOR3xp33_ASAP7_75t_L g3007 ( 
.A(n_2595),
.B(n_20),
.C(n_19),
.Y(n_3007)
);

INVx4_ASAP7_75t_L g3008 ( 
.A(n_2535),
.Y(n_3008)
);

NAND2xp33_ASAP7_75t_L g3009 ( 
.A(n_2385),
.B(n_20),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2601),
.B(n_17),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2536),
.B(n_21),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2581),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_SL g3013 ( 
.A(n_2417),
.B(n_21),
.Y(n_3013)
);

O2A1O1Ixp33_ASAP7_75t_L g3014 ( 
.A1(n_2476),
.A2(n_23),
.B(n_20),
.C(n_22),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2414),
.B(n_22),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2432),
.B(n_23),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_SL g3017 ( 
.A(n_2407),
.B(n_25),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2582),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2407),
.B(n_26),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2584),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2387),
.B(n_24),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2460),
.B(n_24),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2573),
.B(n_26),
.Y(n_3023)
);

INVx2_ASAP7_75t_SL g3024 ( 
.A(n_2436),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_SL g3025 ( 
.A(n_2469),
.B(n_28),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2586),
.Y(n_3026)
);

INVx2_ASAP7_75t_SL g3027 ( 
.A(n_2587),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2485),
.Y(n_3028)
);

OAI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2309),
.A2(n_27),
.B(n_28),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2512),
.B(n_27),
.Y(n_3030)
);

NOR3xp33_ASAP7_75t_L g3031 ( 
.A(n_2588),
.B(n_31),
.C(n_30),
.Y(n_3031)
);

BUFx6f_ASAP7_75t_L g3032 ( 
.A(n_2499),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2558),
.Y(n_3033)
);

INVx3_ASAP7_75t_L g3034 ( 
.A(n_2585),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2597),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2539),
.B(n_29),
.Y(n_3036)
);

INVx2_ASAP7_75t_SL g3037 ( 
.A(n_2489),
.Y(n_3037)
);

AOI22xp33_ASAP7_75t_L g3038 ( 
.A1(n_2598),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_3038)
);

BUFx2_ASAP7_75t_L g3039 ( 
.A(n_2499),
.Y(n_3039)
);

INVx3_ASAP7_75t_L g3040 ( 
.A(n_2499),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2591),
.B(n_29),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2600),
.Y(n_3042)
);

AND2x2_ASAP7_75t_L g3043 ( 
.A(n_2603),
.B(n_31),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2593),
.B(n_32),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_SL g3045 ( 
.A(n_2542),
.B(n_33),
.Y(n_3045)
);

BUFx3_ASAP7_75t_L g3046 ( 
.A(n_2542),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2542),
.B(n_32),
.Y(n_3047)
);

BUFx6f_ASAP7_75t_L g3048 ( 
.A(n_2309),
.Y(n_3048)
);

OAI22xp5_ASAP7_75t_L g3049 ( 
.A1(n_2497),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2497),
.B(n_34),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2497),
.B(n_33),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2610),
.Y(n_3052)
);

INVx1_ASAP7_75t_SL g3053 ( 
.A(n_2647),
.Y(n_3053)
);

O2A1O1Ixp33_ASAP7_75t_L g3054 ( 
.A1(n_2521),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_3054)
);

AO22x2_ASAP7_75t_L g3055 ( 
.A1(n_2647),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2488),
.B(n_35),
.Y(n_3056)
);

NAND2xp33_ASAP7_75t_SL g3057 ( 
.A(n_2392),
.B(n_38),
.Y(n_3057)
);

NOR3xp33_ASAP7_75t_L g3058 ( 
.A(n_2624),
.B(n_40),
.C(n_39),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2488),
.B(n_38),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2392),
.B(n_38),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2392),
.B(n_39),
.Y(n_3061)
);

BUFx8_ASAP7_75t_L g3062 ( 
.A(n_2318),
.Y(n_3062)
);

INVx2_ASAP7_75t_SL g3063 ( 
.A(n_2344),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2610),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2610),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2392),
.B(n_40),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2392),
.B(n_40),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2647),
.B(n_42),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2647),
.B(n_42),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2610),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2610),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2647),
.B(n_42),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2392),
.B(n_41),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2610),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2392),
.B(n_41),
.Y(n_3075)
);

INVx3_ASAP7_75t_L g3076 ( 
.A(n_2444),
.Y(n_3076)
);

AND2x4_ASAP7_75t_L g3077 ( 
.A(n_2392),
.B(n_43),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2610),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2610),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2392),
.B(n_43),
.Y(n_3080)
);

NAND2x1p5_ASAP7_75t_L g3081 ( 
.A(n_2267),
.B(n_43),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2647),
.B(n_45),
.Y(n_3082)
);

BUFx3_ASAP7_75t_L g3083 ( 
.A(n_2548),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2647),
.B(n_44),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2488),
.B(n_44),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2610),
.Y(n_3086)
);

INVx3_ASAP7_75t_L g3087 ( 
.A(n_2444),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2610),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2392),
.B(n_44),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2392),
.B(n_45),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2444),
.Y(n_3091)
);

NOR3xp33_ASAP7_75t_L g3092 ( 
.A(n_2624),
.B(n_47),
.C(n_46),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2392),
.B(n_45),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_SL g3094 ( 
.A(n_2647),
.B(n_47),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2610),
.Y(n_3095)
);

OR2x6_ASAP7_75t_L g3096 ( 
.A(n_2631),
.B(n_46),
.Y(n_3096)
);

AOI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_2395),
.A2(n_49),
.B1(n_46),
.B2(n_48),
.Y(n_3097)
);

OAI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2392),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2392),
.B(n_48),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2610),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2610),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2610),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2392),
.B(n_49),
.Y(n_3103)
);

AOI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2395),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_3104)
);

INVx2_ASAP7_75t_SL g3105 ( 
.A(n_2344),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2392),
.B(n_50),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2610),
.Y(n_3107)
);

OAI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_2332),
.A2(n_55),
.B1(n_52),
.B2(n_53),
.Y(n_3108)
);

AO221x1_ASAP7_75t_L g3109 ( 
.A1(n_2351),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.C(n_57),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2610),
.Y(n_3110)
);

NOR3xp33_ASAP7_75t_L g3111 ( 
.A(n_2624),
.B(n_56),
.C(n_55),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2647),
.B(n_56),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2610),
.Y(n_3113)
);

NOR2xp67_ASAP7_75t_SL g3114 ( 
.A(n_2631),
.B(n_53),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2392),
.B(n_58),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2392),
.B(n_59),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2610),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2392),
.B(n_59),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_2647),
.Y(n_3119)
);

NOR3xp33_ASAP7_75t_L g3120 ( 
.A(n_2624),
.B(n_61),
.C(n_60),
.Y(n_3120)
);

BUFx6f_ASAP7_75t_SL g3121 ( 
.A(n_2318),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2610),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2392),
.B(n_59),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2392),
.B(n_60),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_SL g3125 ( 
.A(n_2647),
.B(n_62),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2488),
.B(n_61),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2392),
.B(n_63),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2610),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2488),
.B(n_63),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_SL g3130 ( 
.A(n_2647),
.B(n_64),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2392),
.B(n_63),
.Y(n_3131)
);

INVx2_ASAP7_75t_SL g3132 ( 
.A(n_2344),
.Y(n_3132)
);

INVx2_ASAP7_75t_SL g3133 ( 
.A(n_2344),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2392),
.B(n_64),
.Y(n_3134)
);

INVxp67_ASAP7_75t_L g3135 ( 
.A(n_2647),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_L g3136 ( 
.A(n_2488),
.B(n_64),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2392),
.B(n_65),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_2647),
.B(n_66),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2381),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_3139)
);

BUFx8_ASAP7_75t_L g3140 ( 
.A(n_2318),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2610),
.Y(n_3141)
);

INVx2_ASAP7_75t_SL g3142 ( 
.A(n_2344),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_SL g3143 ( 
.A(n_2647),
.B(n_67),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2392),
.B(n_66),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2610),
.Y(n_3145)
);

NOR2xp33_ASAP7_75t_L g3146 ( 
.A(n_2488),
.B(n_67),
.Y(n_3146)
);

AND2x2_ASAP7_75t_SL g3147 ( 
.A(n_2538),
.B(n_68),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2392),
.B(n_68),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2392),
.B(n_68),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2610),
.Y(n_3150)
);

OAI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_2392),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2392),
.B(n_69),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2610),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2392),
.B(n_69),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2392),
.B(n_70),
.Y(n_3155)
);

OAI22xp5_ASAP7_75t_L g3156 ( 
.A1(n_2392),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_2395),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_3157)
);

NOR3xp33_ASAP7_75t_L g3158 ( 
.A(n_2624),
.B(n_75),
.C(n_74),
.Y(n_3158)
);

AOI22xp5_ASAP7_75t_L g3159 ( 
.A1(n_2395),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_3159)
);

NOR3xp33_ASAP7_75t_L g3160 ( 
.A(n_2624),
.B(n_77),
.C(n_76),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_SL g3161 ( 
.A(n_2647),
.B(n_76),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2392),
.B(n_75),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2610),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2610),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2392),
.B(n_76),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2392),
.B(n_77),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2392),
.B(n_78),
.Y(n_3167)
);

NOR2xp33_ASAP7_75t_L g3168 ( 
.A(n_2488),
.B(n_78),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2392),
.B(n_78),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2610),
.Y(n_3170)
);

INVxp67_ASAP7_75t_L g3171 ( 
.A(n_2647),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2392),
.B(n_79),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2392),
.B(n_79),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2610),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2610),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2610),
.Y(n_3176)
);

OR2x2_ASAP7_75t_L g3177 ( 
.A(n_2647),
.B(n_80),
.Y(n_3177)
);

OR2x6_ASAP7_75t_L g3178 ( 
.A(n_2631),
.B(n_80),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2392),
.B(n_80),
.Y(n_3179)
);

INVx1_ASAP7_75t_SL g3180 ( 
.A(n_2647),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_SL g3181 ( 
.A(n_2647),
.B(n_82),
.Y(n_3181)
);

OAI22xp5_ASAP7_75t_L g3182 ( 
.A1(n_2392),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3182)
);

INVx2_ASAP7_75t_SL g3183 ( 
.A(n_2344),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_2488),
.B(n_81),
.Y(n_3184)
);

OAI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_2392),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2610),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_2610),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2392),
.B(n_83),
.Y(n_3188)
);

OAI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2508),
.A2(n_84),
.B(n_85),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2392),
.B(n_84),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2610),
.Y(n_3191)
);

OAI22x1_ASAP7_75t_R g3192 ( 
.A1(n_2404),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_3192)
);

NAND3xp33_ASAP7_75t_L g3193 ( 
.A(n_2519),
.B(n_85),
.C(n_86),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_SL g3194 ( 
.A(n_2647),
.B(n_87),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_2647),
.B(n_86),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2610),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2392),
.B(n_87),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2392),
.B(n_88),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_SL g3199 ( 
.A(n_2647),
.B(n_89),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2392),
.B(n_88),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_SL g3201 ( 
.A(n_2647),
.B(n_90),
.Y(n_3201)
);

HB1xp67_ASAP7_75t_L g3202 ( 
.A(n_2647),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2392),
.B(n_89),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_SL g3204 ( 
.A(n_2647),
.B(n_91),
.Y(n_3204)
);

INVx1_ASAP7_75t_SL g3205 ( 
.A(n_2647),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2392),
.B(n_90),
.Y(n_3206)
);

NOR2xp67_ASAP7_75t_L g3207 ( 
.A(n_2623),
.B(n_90),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2610),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2392),
.B(n_91),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_2647),
.B(n_91),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2392),
.B(n_92),
.Y(n_3211)
);

INVxp67_ASAP7_75t_L g3212 ( 
.A(n_2647),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2392),
.B(n_92),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2392),
.B(n_92),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2610),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_SL g3216 ( 
.A(n_2647),
.B(n_94),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2392),
.B(n_93),
.Y(n_3217)
);

NOR2xp67_ASAP7_75t_L g3218 ( 
.A(n_2623),
.B(n_93),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2392),
.B(n_93),
.Y(n_3219)
);

AND2x2_ASAP7_75t_SL g3220 ( 
.A(n_2538),
.B(n_94),
.Y(n_3220)
);

INVx8_ASAP7_75t_L g3221 ( 
.A(n_2267),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2392),
.B(n_94),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2610),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_2488),
.B(n_95),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2610),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2392),
.B(n_95),
.Y(n_3226)
);

INVx2_ASAP7_75t_SL g3227 ( 
.A(n_2344),
.Y(n_3227)
);

INVx3_ASAP7_75t_L g3228 ( 
.A(n_2444),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2610),
.Y(n_3229)
);

AOI22xp33_ASAP7_75t_L g3230 ( 
.A1(n_2381),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_2647),
.B(n_97),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2610),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2392),
.B(n_96),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2610),
.Y(n_3234)
);

BUFx3_ASAP7_75t_L g3235 ( 
.A(n_2548),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_2647),
.B(n_96),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_2488),
.B(n_97),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2610),
.Y(n_3238)
);

NOR3xp33_ASAP7_75t_L g3239 ( 
.A(n_2624),
.B(n_100),
.C(n_99),
.Y(n_3239)
);

INVxp67_ASAP7_75t_L g3240 ( 
.A(n_2647),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2610),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2610),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2392),
.B(n_98),
.Y(n_3243)
);

BUFx6f_ASAP7_75t_L g3244 ( 
.A(n_2444),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2392),
.B(n_98),
.Y(n_3245)
);

AND2x4_ASAP7_75t_L g3246 ( 
.A(n_2392),
.B(n_98),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2392),
.B(n_99),
.Y(n_3247)
);

BUFx3_ASAP7_75t_L g3248 ( 
.A(n_2548),
.Y(n_3248)
);

AND2x4_ASAP7_75t_L g3249 ( 
.A(n_2392),
.B(n_99),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2610),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2392),
.B(n_100),
.Y(n_3251)
);

BUFx6f_ASAP7_75t_L g3252 ( 
.A(n_2444),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_L g3253 ( 
.A(n_2488),
.B(n_100),
.Y(n_3253)
);

AND2x4_ASAP7_75t_L g3254 ( 
.A(n_2392),
.B(n_101),
.Y(n_3254)
);

AND2x6_ASAP7_75t_L g3255 ( 
.A(n_2392),
.B(n_101),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2610),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_2610),
.Y(n_3257)
);

NOR3xp33_ASAP7_75t_L g3258 ( 
.A(n_2624),
.B(n_104),
.C(n_103),
.Y(n_3258)
);

NAND2x1_ASAP7_75t_L g3259 ( 
.A(n_2289),
.B(n_102),
.Y(n_3259)
);

OAI221xp5_ASAP7_75t_L g3260 ( 
.A1(n_2395),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.C(n_106),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2392),
.B(n_105),
.Y(n_3261)
);

HB1xp67_ASAP7_75t_L g3262 ( 
.A(n_2647),
.Y(n_3262)
);

INVx2_ASAP7_75t_SL g3263 ( 
.A(n_2344),
.Y(n_3263)
);

BUFx2_ASAP7_75t_L g3264 ( 
.A(n_2647),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_2392),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_3265)
);

NOR2xp33_ASAP7_75t_L g3266 ( 
.A(n_2488),
.B(n_106),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2647),
.B(n_108),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_SL g3268 ( 
.A(n_2647),
.B(n_108),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_2647),
.B(n_107),
.Y(n_3269)
);

O2A1O1Ixp33_ASAP7_75t_L g3270 ( 
.A1(n_2521),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_2392),
.B(n_109),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_SL g3272 ( 
.A(n_2647),
.B(n_110),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_2395),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2392),
.B(n_111),
.Y(n_3274)
);

O2A1O1Ixp33_ASAP7_75t_L g3275 ( 
.A1(n_2521),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2392),
.B(n_112),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2392),
.B(n_112),
.Y(n_3277)
);

INVx2_ASAP7_75t_SL g3278 ( 
.A(n_2344),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2610),
.Y(n_3279)
);

CKINVDCx5p33_ASAP7_75t_R g3280 ( 
.A(n_2623),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2392),
.B(n_113),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2392),
.B(n_113),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2610),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_2610),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2392),
.B(n_114),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2392),
.B(n_115),
.Y(n_3286)
);

INVx3_ASAP7_75t_L g3287 ( 
.A(n_2444),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2488),
.B(n_116),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2392),
.B(n_116),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2610),
.Y(n_3290)
);

NAND3xp33_ASAP7_75t_L g3291 ( 
.A(n_2519),
.B(n_116),
.C(n_117),
.Y(n_3291)
);

CKINVDCx5p33_ASAP7_75t_R g3292 ( 
.A(n_3062),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2650),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2657),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2878),
.B(n_117),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2736),
.B(n_117),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_SL g3297 ( 
.A(n_3053),
.B(n_3180),
.Y(n_3297)
);

BUFx6f_ASAP7_75t_L g3298 ( 
.A(n_2701),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2817),
.B(n_118),
.Y(n_3299)
);

CKINVDCx20_ASAP7_75t_R g3300 ( 
.A(n_3062),
.Y(n_3300)
);

NOR2xp33_ASAP7_75t_L g3301 ( 
.A(n_2722),
.B(n_2725),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3052),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_2817),
.B(n_118),
.Y(n_3303)
);

OAI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_3096),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_3304)
);

AND2x4_ASAP7_75t_L g3305 ( 
.A(n_3283),
.B(n_119),
.Y(n_3305)
);

AOI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3147),
.A2(n_3220),
.B1(n_2763),
.B2(n_2754),
.Y(n_3306)
);

NOR2xp33_ASAP7_75t_L g3307 ( 
.A(n_2742),
.B(n_120),
.Y(n_3307)
);

NOR3xp33_ASAP7_75t_L g3308 ( 
.A(n_3260),
.B(n_120),
.C(n_121),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3064),
.Y(n_3309)
);

NOR2x1_ASAP7_75t_L g3310 ( 
.A(n_3096),
.B(n_121),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3086),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2653),
.B(n_121),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3088),
.Y(n_3313)
);

NAND2xp33_ASAP7_75t_L g3314 ( 
.A(n_2924),
.B(n_122),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_2755),
.B(n_122),
.Y(n_3315)
);

BUFx3_ASAP7_75t_L g3316 ( 
.A(n_3140),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2655),
.B(n_122),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_L g3318 ( 
.A(n_2787),
.B(n_123),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3284),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_SL g3320 ( 
.A(n_3053),
.B(n_577),
.Y(n_3320)
);

HB1xp67_ASAP7_75t_L g3321 ( 
.A(n_3119),
.Y(n_3321)
);

INVx3_ASAP7_75t_L g3322 ( 
.A(n_3221),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2659),
.B(n_123),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3065),
.B(n_123),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3102),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_2926),
.A2(n_124),
.B(n_125),
.Y(n_3326)
);

INVx2_ASAP7_75t_SL g3327 ( 
.A(n_3221),
.Y(n_3327)
);

AOI22xp5_ASAP7_75t_L g3328 ( 
.A1(n_2763),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3070),
.B(n_126),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3107),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_3117),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_2686),
.B(n_126),
.Y(n_3332)
);

AND2x4_ASAP7_75t_L g3333 ( 
.A(n_3141),
.B(n_127),
.Y(n_3333)
);

NOR3xp33_ASAP7_75t_SL g3334 ( 
.A(n_2782),
.B(n_127),
.C(n_128),
.Y(n_3334)
);

AND2x4_ASAP7_75t_L g3335 ( 
.A(n_3153),
.B(n_127),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3175),
.Y(n_3336)
);

BUFx4f_ASAP7_75t_L g3337 ( 
.A(n_3096),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3071),
.B(n_128),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3186),
.Y(n_3339)
);

AND2x4_ASAP7_75t_L g3340 ( 
.A(n_3187),
.B(n_129),
.Y(n_3340)
);

OAI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_3077),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3196),
.Y(n_3342)
);

BUFx2_ASAP7_75t_L g3343 ( 
.A(n_3264),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_3180),
.B(n_3205),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3074),
.B(n_129),
.Y(n_3345)
);

BUFx3_ASAP7_75t_L g3346 ( 
.A(n_3140),
.Y(n_3346)
);

AND2x4_ASAP7_75t_L g3347 ( 
.A(n_3208),
.B(n_130),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3225),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3234),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_SL g3350 ( 
.A(n_3205),
.B(n_577),
.Y(n_3350)
);

INVx2_ASAP7_75t_SL g3351 ( 
.A(n_3221),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_2686),
.B(n_131),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3238),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3078),
.B(n_132),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3079),
.B(n_132),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3095),
.B(n_133),
.Y(n_3356)
);

NOR2x1p5_ASAP7_75t_L g3357 ( 
.A(n_2766),
.B(n_133),
.Y(n_3357)
);

CKINVDCx5p33_ASAP7_75t_R g3358 ( 
.A(n_3121),
.Y(n_3358)
);

AND2x4_ASAP7_75t_L g3359 ( 
.A(n_3242),
.B(n_133),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3250),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_3121),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3100),
.B(n_134),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3257),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_2668),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_R g3365 ( 
.A(n_2714),
.B(n_134),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_3135),
.B(n_3171),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_2933),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3101),
.B(n_135),
.Y(n_3368)
);

HB1xp67_ASAP7_75t_L g3369 ( 
.A(n_3202),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3110),
.B(n_136),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2670),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3113),
.B(n_136),
.Y(n_3372)
);

INVx1_ASAP7_75t_SL g3373 ( 
.A(n_3262),
.Y(n_3373)
);

NOR3xp33_ASAP7_75t_L g3374 ( 
.A(n_2999),
.B(n_137),
.C(n_138),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_2675),
.Y(n_3375)
);

CKINVDCx11_ASAP7_75t_R g3376 ( 
.A(n_2747),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_2933),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_3377)
);

NAND3xp33_ASAP7_75t_SL g3378 ( 
.A(n_2667),
.B(n_2674),
.C(n_2662),
.Y(n_3378)
);

BUFx6f_ASAP7_75t_L g3379 ( 
.A(n_2701),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3122),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3128),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3145),
.B(n_137),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3150),
.Y(n_3383)
);

BUFx4f_ASAP7_75t_L g3384 ( 
.A(n_3178),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_R g3385 ( 
.A(n_3280),
.B(n_2708),
.Y(n_3385)
);

AOI21xp33_ASAP7_75t_L g3386 ( 
.A1(n_2658),
.A2(n_138),
.B(n_139),
.Y(n_3386)
);

NOR2xp33_ASAP7_75t_L g3387 ( 
.A(n_2988),
.B(n_2938),
.Y(n_3387)
);

OR2x6_ASAP7_75t_L g3388 ( 
.A(n_3178),
.B(n_139),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3163),
.B(n_140),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3164),
.B(n_140),
.Y(n_3390)
);

INVx4_ASAP7_75t_L g3391 ( 
.A(n_3178),
.Y(n_3391)
);

CKINVDCx5p33_ASAP7_75t_R g3392 ( 
.A(n_2708),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3170),
.B(n_141),
.Y(n_3393)
);

BUFx6f_ASAP7_75t_L g3394 ( 
.A(n_2701),
.Y(n_3394)
);

AOI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_2682),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_2683),
.Y(n_3396)
);

NOR2x1p5_ASAP7_75t_L g3397 ( 
.A(n_3083),
.B(n_142),
.Y(n_3397)
);

O2A1O1Ixp33_ASAP7_75t_L g3398 ( 
.A1(n_2706),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_3398)
);

NOR3xp33_ASAP7_75t_SL g3399 ( 
.A(n_3108),
.B(n_143),
.C(n_144),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_2747),
.Y(n_3400)
);

BUFx6f_ASAP7_75t_L g3401 ( 
.A(n_2769),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3174),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_2709),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_2666),
.B(n_145),
.Y(n_3404)
);

NOR2xp33_ASAP7_75t_L g3405 ( 
.A(n_2896),
.B(n_146),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_2739),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3176),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3191),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3215),
.Y(n_3409)
);

INVxp67_ASAP7_75t_L g3410 ( 
.A(n_2680),
.Y(n_3410)
);

HB1xp67_ASAP7_75t_L g3411 ( 
.A(n_3212),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_2678),
.B(n_3240),
.Y(n_3412)
);

BUFx6f_ASAP7_75t_L g3413 ( 
.A(n_2769),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3223),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3229),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3232),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_2667),
.B(n_2769),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_2698),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2702),
.Y(n_3419)
);

OR2x6_ASAP7_75t_L g3420 ( 
.A(n_2843),
.B(n_146),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3241),
.B(n_147),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3256),
.Y(n_3422)
);

INVx6_ASAP7_75t_L g3423 ( 
.A(n_2794),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3091),
.B(n_578),
.Y(n_3424)
);

NOR3xp33_ASAP7_75t_SL g3425 ( 
.A(n_2690),
.B(n_147),
.C(n_148),
.Y(n_3425)
);

INVx5_ASAP7_75t_L g3426 ( 
.A(n_3091),
.Y(n_3426)
);

INVx2_ASAP7_75t_SL g3427 ( 
.A(n_2811),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3279),
.B(n_147),
.Y(n_3428)
);

OR2x4_ASAP7_75t_L g3429 ( 
.A(n_2875),
.B(n_148),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_SL g3430 ( 
.A1(n_3255),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_2756),
.Y(n_3431)
);

NAND2xp33_ASAP7_75t_SL g3432 ( 
.A(n_3114),
.B(n_3077),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2786),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_2821),
.Y(n_3434)
);

NAND2x1p5_ASAP7_75t_L g3435 ( 
.A(n_2812),
.B(n_149),
.Y(n_3435)
);

NOR2x2_ASAP7_75t_L g3436 ( 
.A(n_2843),
.B(n_150),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_3091),
.B(n_578),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2844),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3290),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_3244),
.B(n_579),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_2815),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_2848),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2672),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2684),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3235),
.Y(n_3445)
);

AOI22xp5_ASAP7_75t_L g3446 ( 
.A1(n_3106),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_2707),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_2851),
.Y(n_3448)
);

NOR2x1p5_ASAP7_75t_L g3449 ( 
.A(n_3248),
.B(n_151),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3244),
.B(n_579),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_2860),
.B(n_152),
.Y(n_3451)
);

BUFx3_ASAP7_75t_L g3452 ( 
.A(n_2721),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_2693),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_2879),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_2836),
.B(n_152),
.Y(n_3455)
);

INVx1_ASAP7_75t_SL g3456 ( 
.A(n_2773),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_2717),
.B(n_153),
.Y(n_3457)
);

BUFx3_ASAP7_75t_L g3458 ( 
.A(n_2726),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_2732),
.B(n_153),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_2729),
.B(n_154),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_2710),
.B(n_154),
.Y(n_3461)
);

AOI22xp5_ASAP7_75t_L g3462 ( 
.A1(n_3106),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_2734),
.Y(n_3463)
);

INVxp67_ASAP7_75t_L g3464 ( 
.A(n_2685),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_2735),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2741),
.Y(n_3466)
);

INVx3_ASAP7_75t_L g3467 ( 
.A(n_2707),
.Y(n_3467)
);

INVx3_ASAP7_75t_L g3468 ( 
.A(n_3008),
.Y(n_3468)
);

AOI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_3246),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_2843),
.Y(n_3470)
);

NAND3xp33_ASAP7_75t_SL g3471 ( 
.A(n_2674),
.B(n_155),
.C(n_157),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2760),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_SL g3473 ( 
.A(n_3244),
.B(n_580),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_2715),
.B(n_158),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_3252),
.B(n_580),
.Y(n_3475)
);

AND2x2_ASAP7_75t_L g3476 ( 
.A(n_3246),
.B(n_159),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_2765),
.Y(n_3477)
);

AND2x4_ASAP7_75t_L g3478 ( 
.A(n_2983),
.B(n_159),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_2768),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_2774),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_2776),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2718),
.B(n_160),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_2987),
.A2(n_161),
.B(n_162),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_2777),
.Y(n_3484)
);

INVx4_ASAP7_75t_L g3485 ( 
.A(n_3252),
.Y(n_3485)
);

INVx3_ASAP7_75t_L g3486 ( 
.A(n_3008),
.Y(n_3486)
);

INVx8_ASAP7_75t_L g3487 ( 
.A(n_2802),
.Y(n_3487)
);

AND2x4_ASAP7_75t_L g3488 ( 
.A(n_3249),
.B(n_3254),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_2797),
.B(n_161),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_2781),
.Y(n_3490)
);

INVx1_ASAP7_75t_SL g3491 ( 
.A(n_2792),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_2941),
.B(n_161),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_2788),
.Y(n_3493)
);

AND2x2_ASAP7_75t_L g3494 ( 
.A(n_3249),
.B(n_162),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_L g3495 ( 
.A(n_2908),
.B(n_2958),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_2791),
.Y(n_3496)
);

OR2x2_ASAP7_75t_SL g3497 ( 
.A(n_3192),
.B(n_162),
.Y(n_3497)
);

BUFx3_ASAP7_75t_L g3498 ( 
.A(n_3063),
.Y(n_3498)
);

INVx1_ASAP7_75t_SL g3499 ( 
.A(n_2906),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_3252),
.B(n_581),
.Y(n_3500)
);

BUFx2_ASAP7_75t_L g3501 ( 
.A(n_2802),
.Y(n_3501)
);

INVx2_ASAP7_75t_SL g3502 ( 
.A(n_3105),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_2887),
.B(n_163),
.Y(n_3503)
);

BUFx3_ASAP7_75t_L g3504 ( 
.A(n_3132),
.Y(n_3504)
);

INVx1_ASAP7_75t_SL g3505 ( 
.A(n_3133),
.Y(n_3505)
);

INVx1_ASAP7_75t_SL g3506 ( 
.A(n_3142),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_2888),
.B(n_163),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_2800),
.B(n_163),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_2838),
.B(n_164),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2852),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_2873),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_2871),
.Y(n_3512)
);

INVx3_ASAP7_75t_L g3513 ( 
.A(n_2835),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_2959),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_2872),
.B(n_164),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3060),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3061),
.Y(n_3517)
);

INVx3_ASAP7_75t_L g3518 ( 
.A(n_2841),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_2968),
.Y(n_3519)
);

AND2x4_ASAP7_75t_L g3520 ( 
.A(n_3254),
.B(n_165),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_2886),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_2890),
.Y(n_3522)
);

AO22x1_ASAP7_75t_L g3523 ( 
.A1(n_3255),
.A2(n_2802),
.B1(n_3092),
.B2(n_3058),
.Y(n_3523)
);

HB1xp67_ASAP7_75t_L g3524 ( 
.A(n_2832),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_2733),
.B(n_165),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3066),
.Y(n_3526)
);

INVx1_ASAP7_75t_SL g3527 ( 
.A(n_3183),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3067),
.Y(n_3528)
);

BUFx3_ASAP7_75t_L g3529 ( 
.A(n_3227),
.Y(n_3529)
);

O2A1O1Ixp33_ASAP7_75t_L g3530 ( 
.A1(n_2952),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_2874),
.B(n_166),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_2891),
.Y(n_3532)
);

AND2x4_ASAP7_75t_L g3533 ( 
.A(n_2925),
.B(n_166),
.Y(n_3533)
);

OR2x6_ASAP7_75t_L g3534 ( 
.A(n_2924),
.B(n_167),
.Y(n_3534)
);

INVx2_ASAP7_75t_SL g3535 ( 
.A(n_3263),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_2934),
.B(n_167),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_2826),
.B(n_168),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_2892),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_2688),
.B(n_168),
.Y(n_3539)
);

AND2x6_ASAP7_75t_L g3540 ( 
.A(n_3046),
.B(n_169),
.Y(n_3540)
);

BUFx6f_ASAP7_75t_L g3541 ( 
.A(n_2892),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3073),
.Y(n_3542)
);

AOI22xp33_ASAP7_75t_L g3543 ( 
.A1(n_3057),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_2882),
.B(n_169),
.Y(n_3544)
);

AOI211xp5_ASAP7_75t_L g3545 ( 
.A1(n_3017),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_3545)
);

BUFx6f_ASAP7_75t_L g3546 ( 
.A(n_2892),
.Y(n_3546)
);

INVx2_ASAP7_75t_SL g3547 ( 
.A(n_3278),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_2921),
.Y(n_3548)
);

INVx4_ASAP7_75t_L g3549 ( 
.A(n_2833),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3075),
.Y(n_3550)
);

BUFx6f_ASAP7_75t_L g3551 ( 
.A(n_2924),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3080),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_2840),
.B(n_170),
.Y(n_3553)
);

AND2x6_ASAP7_75t_L g3554 ( 
.A(n_3032),
.B(n_3040),
.Y(n_3554)
);

AOI22xp33_ASAP7_75t_L g3555 ( 
.A1(n_3255),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_3555)
);

HB1xp67_ASAP7_75t_L g3556 ( 
.A(n_3255),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_3084),
.B(n_172),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3089),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_2737),
.B(n_173),
.Y(n_3559)
);

INVx2_ASAP7_75t_SL g3560 ( 
.A(n_2778),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_2673),
.B(n_173),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_2922),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3090),
.Y(n_3563)
);

INVx4_ASAP7_75t_L g3564 ( 
.A(n_2833),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_2928),
.Y(n_3565)
);

BUFx2_ASAP7_75t_L g3566 ( 
.A(n_2802),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3093),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_SL g3568 ( 
.A(n_2796),
.B(n_581),
.Y(n_3568)
);

INVxp67_ASAP7_75t_L g3569 ( 
.A(n_2764),
.Y(n_3569)
);

BUFx8_ASAP7_75t_L g3570 ( 
.A(n_3024),
.Y(n_3570)
);

AND2x4_ASAP7_75t_L g3571 ( 
.A(n_2925),
.B(n_174),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_2679),
.B(n_175),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_R g3573 ( 
.A(n_2772),
.B(n_2730),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3109),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3574)
);

CKINVDCx20_ASAP7_75t_R g3575 ( 
.A(n_2939),
.Y(n_3575)
);

INVx2_ASAP7_75t_SL g3576 ( 
.A(n_2779),
.Y(n_3576)
);

AOI22xp33_ASAP7_75t_L g3577 ( 
.A1(n_2761),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3577)
);

AOI22xp33_ASAP7_75t_L g3578 ( 
.A1(n_2902),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3195),
.B(n_179),
.Y(n_3579)
);

CKINVDCx16_ASAP7_75t_R g3580 ( 
.A(n_2796),
.Y(n_3580)
);

INVx2_ASAP7_75t_SL g3581 ( 
.A(n_2943),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3099),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_SL g3583 ( 
.A(n_2808),
.B(n_582),
.Y(n_3583)
);

NAND2xp33_ASAP7_75t_SL g3584 ( 
.A(n_3032),
.B(n_179),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3103),
.B(n_179),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3115),
.B(n_180),
.Y(n_3586)
);

AND2x4_ASAP7_75t_L g3587 ( 
.A(n_2978),
.B(n_180),
.Y(n_3587)
);

NAND3xp33_ASAP7_75t_L g3588 ( 
.A(n_3111),
.B(n_180),
.C(n_181),
.Y(n_3588)
);

NOR2xp67_ASAP7_75t_L g3589 ( 
.A(n_2895),
.B(n_182),
.Y(n_3589)
);

BUFx3_ASAP7_75t_L g3590 ( 
.A(n_3002),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_SL g3591 ( 
.A(n_2808),
.B(n_583),
.Y(n_3591)
);

INVx4_ASAP7_75t_L g3592 ( 
.A(n_3004),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3116),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3118),
.Y(n_3594)
);

HB1xp67_ASAP7_75t_L g3595 ( 
.A(n_2953),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_2931),
.Y(n_3596)
);

BUFx6f_ASAP7_75t_L g3597 ( 
.A(n_2937),
.Y(n_3597)
);

INVx1_ASAP7_75t_SL g3598 ( 
.A(n_2981),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3123),
.B(n_182),
.Y(n_3599)
);

NAND2xp33_ASAP7_75t_SL g3600 ( 
.A(n_3032),
.B(n_183),
.Y(n_3600)
);

INVx3_ASAP7_75t_L g3601 ( 
.A(n_2898),
.Y(n_3601)
);

INVx2_ASAP7_75t_SL g3602 ( 
.A(n_2713),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_2951),
.Y(n_3603)
);

AND2x4_ASAP7_75t_L g3604 ( 
.A(n_2842),
.B(n_183),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_2963),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3124),
.B(n_183),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3127),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3131),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3134),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_2976),
.Y(n_3610)
);

CKINVDCx5p33_ASAP7_75t_R g3611 ( 
.A(n_3004),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_2977),
.Y(n_3612)
);

BUFx4f_ASAP7_75t_L g3613 ( 
.A(n_3081),
.Y(n_3613)
);

AND2x4_ASAP7_75t_L g3614 ( 
.A(n_2656),
.B(n_184),
.Y(n_3614)
);

INVx4_ASAP7_75t_L g3615 ( 
.A(n_3081),
.Y(n_3615)
);

AND2x2_ASAP7_75t_SL g3616 ( 
.A(n_2979),
.B(n_184),
.Y(n_3616)
);

HB1xp67_ASAP7_75t_L g3617 ( 
.A(n_2986),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3137),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3144),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3148),
.Y(n_3620)
);

OR2x6_ASAP7_75t_L g3621 ( 
.A(n_2937),
.B(n_2969),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_2889),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3149),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3152),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_2897),
.Y(n_3625)
);

A2O1A1Ixp33_ASAP7_75t_L g3626 ( 
.A1(n_3054),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_3626)
);

INVx4_ASAP7_75t_L g3627 ( 
.A(n_2898),
.Y(n_3627)
);

AOI22xp33_ASAP7_75t_L g3628 ( 
.A1(n_3056),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_3628)
);

INVx4_ASAP7_75t_L g3629 ( 
.A(n_2937),
.Y(n_3629)
);

INVx2_ASAP7_75t_SL g3630 ( 
.A(n_3006),
.Y(n_3630)
);

AND2x2_ASAP7_75t_SL g3631 ( 
.A(n_3009),
.B(n_186),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3154),
.B(n_187),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3155),
.Y(n_3633)
);

INVx4_ASAP7_75t_L g3634 ( 
.A(n_2927),
.Y(n_3634)
);

INVx4_ASAP7_75t_L g3635 ( 
.A(n_2927),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3162),
.B(n_3276),
.Y(n_3636)
);

INVx2_ASAP7_75t_L g3637 ( 
.A(n_2900),
.Y(n_3637)
);

INVxp67_ASAP7_75t_L g3638 ( 
.A(n_3177),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3165),
.B(n_187),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_R g3640 ( 
.A(n_2969),
.B(n_188),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3166),
.Y(n_3641)
);

INVx2_ASAP7_75t_SL g3642 ( 
.A(n_3006),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3167),
.Y(n_3643)
);

INVx1_ASAP7_75t_SL g3644 ( 
.A(n_3023),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3169),
.Y(n_3645)
);

INVx5_ASAP7_75t_L g3646 ( 
.A(n_2969),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_2663),
.B(n_584),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3172),
.B(n_189),
.Y(n_3648)
);

CKINVDCx11_ASAP7_75t_R g3649 ( 
.A(n_2827),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3173),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_R g3651 ( 
.A(n_2916),
.B(n_189),
.Y(n_3651)
);

INVx3_ASAP7_75t_L g3652 ( 
.A(n_2935),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_2691),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3179),
.Y(n_3654)
);

AOI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_2687),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_2656),
.B(n_190),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3210),
.B(n_3236),
.Y(n_3657)
);

INVx2_ASAP7_75t_SL g3658 ( 
.A(n_3027),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3188),
.B(n_3190),
.Y(n_3659)
);

AND3x2_ASAP7_75t_SL g3660 ( 
.A(n_2703),
.B(n_191),
.C(n_193),
.Y(n_3660)
);

AOI22xp5_ASAP7_75t_L g3661 ( 
.A1(n_2705),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_3661)
);

AOI22xp5_ASAP7_75t_L g3662 ( 
.A1(n_2762),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_3662)
);

BUFx6f_ASAP7_75t_L g3663 ( 
.A(n_2689),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3197),
.B(n_194),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3198),
.B(n_196),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_2903),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_2910),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_SL g3668 ( 
.A(n_2916),
.B(n_584),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_SL g3669 ( 
.A(n_2918),
.B(n_586),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_2913),
.Y(n_3670)
);

AOI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_2801),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_3671)
);

NOR2xp33_ASAP7_75t_L g3672 ( 
.A(n_2917),
.B(n_196),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3200),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_2813),
.B(n_198),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3203),
.B(n_198),
.Y(n_3675)
);

OR2x6_ASAP7_75t_L g3676 ( 
.A(n_2789),
.B(n_199),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3206),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3209),
.B(n_199),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3211),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3213),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_L g3681 ( 
.A(n_2738),
.B(n_200),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_2915),
.Y(n_3682)
);

NOR2xp33_ASAP7_75t_L g3683 ( 
.A(n_2744),
.B(n_200),
.Y(n_3683)
);

AOI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3059),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_3684)
);

AND2x4_ASAP7_75t_L g3685 ( 
.A(n_2751),
.B(n_201),
.Y(n_3685)
);

AOI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_2984),
.A2(n_2885),
.B(n_2946),
.Y(n_3686)
);

NOR3xp33_ASAP7_75t_SL g3687 ( 
.A(n_3019),
.B(n_201),
.C(n_202),
.Y(n_3687)
);

INVx3_ASAP7_75t_L g3688 ( 
.A(n_2935),
.Y(n_3688)
);

NOR3xp33_ASAP7_75t_SL g3689 ( 
.A(n_3068),
.B(n_203),
.C(n_204),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3214),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3018),
.Y(n_3691)
);

OAI22xp5_ASAP7_75t_SL g3692 ( 
.A1(n_3037),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_3692)
);

CKINVDCx5p33_ASAP7_75t_R g3693 ( 
.A(n_3021),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3217),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3219),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3020),
.Y(n_3696)
);

INVx5_ASAP7_75t_L g3697 ( 
.A(n_2751),
.Y(n_3697)
);

INVx3_ASAP7_75t_L g3698 ( 
.A(n_2696),
.Y(n_3698)
);

NOR2x2_ASAP7_75t_L g3699 ( 
.A(n_3012),
.B(n_3026),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3222),
.Y(n_3700)
);

AOI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_2803),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3035),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_2918),
.B(n_586),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_SL g3704 ( 
.A(n_2942),
.B(n_587),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3226),
.B(n_205),
.Y(n_3705)
);

INVx3_ASAP7_75t_L g3706 ( 
.A(n_2696),
.Y(n_3706)
);

AOI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_2671),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3233),
.B(n_207),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3243),
.B(n_207),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_SL g3710 ( 
.A(n_2942),
.B(n_588),
.Y(n_3710)
);

BUFx2_ASAP7_75t_SL g3711 ( 
.A(n_2716),
.Y(n_3711)
);

A2O1A1Ixp33_ASAP7_75t_L g3712 ( 
.A1(n_3270),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3245),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3247),
.Y(n_3714)
);

OR2x2_ASAP7_75t_L g3715 ( 
.A(n_2692),
.B(n_209),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3251),
.Y(n_3716)
);

INVx2_ASAP7_75t_SL g3717 ( 
.A(n_2966),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_2669),
.B(n_209),
.Y(n_3718)
);

NOR2xp33_ASAP7_75t_L g3719 ( 
.A(n_2759),
.B(n_210),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3261),
.B(n_3271),
.Y(n_3720)
);

AOI22xp5_ASAP7_75t_L g3721 ( 
.A1(n_2660),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_3721)
);

INVx5_ASAP7_75t_L g3722 ( 
.A(n_2810),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3274),
.B(n_211),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3277),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3281),
.B(n_3282),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_SL g3726 ( 
.A(n_2719),
.B(n_589),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3042),
.Y(n_3727)
);

BUFx4f_ASAP7_75t_L g3728 ( 
.A(n_2829),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3285),
.B(n_212),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_SL g3730 ( 
.A(n_2719),
.B(n_2828),
.Y(n_3730)
);

BUFx2_ASAP7_75t_L g3731 ( 
.A(n_2689),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3286),
.Y(n_3732)
);

NOR2xp33_ASAP7_75t_L g3733 ( 
.A(n_2704),
.B(n_213),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_2992),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_3001),
.Y(n_3735)
);

AND2x4_ASAP7_75t_L g3736 ( 
.A(n_2810),
.B(n_213),
.Y(n_3736)
);

AND2x2_ASAP7_75t_SL g3737 ( 
.A(n_3097),
.B(n_214),
.Y(n_3737)
);

NOR2xp33_ASAP7_75t_L g3738 ( 
.A(n_2731),
.B(n_214),
.Y(n_3738)
);

NAND3xp33_ASAP7_75t_SL g3739 ( 
.A(n_3097),
.B(n_3157),
.C(n_3104),
.Y(n_3739)
);

AO22x1_ASAP7_75t_L g3740 ( 
.A1(n_3120),
.A2(n_3160),
.B1(n_3239),
.B2(n_3158),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3289),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_2901),
.B(n_215),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_2824),
.B(n_215),
.Y(n_3743)
);

NOR2xp33_ASAP7_75t_L g3744 ( 
.A(n_2695),
.B(n_216),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3044),
.Y(n_3745)
);

AND2x4_ASAP7_75t_L g3746 ( 
.A(n_3076),
.B(n_216),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_2830),
.B(n_216),
.Y(n_3747)
);

INVx3_ASAP7_75t_L g3748 ( 
.A(n_3076),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3003),
.Y(n_3749)
);

AND2x4_ASAP7_75t_L g3750 ( 
.A(n_3087),
.B(n_217),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3043),
.Y(n_3751)
);

OAI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3104),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3036),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_2991),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_2831),
.B(n_217),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_2652),
.B(n_218),
.Y(n_3756)
);

INVx5_ASAP7_75t_L g3757 ( 
.A(n_3087),
.Y(n_3757)
);

INVx5_ASAP7_75t_L g3758 ( 
.A(n_3228),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3228),
.Y(n_3759)
);

AND2x6_ASAP7_75t_L g3760 ( 
.A(n_3040),
.B(n_218),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_2985),
.Y(n_3761)
);

A2O1A1Ixp33_ASAP7_75t_L g3762 ( 
.A1(n_3275),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3085),
.B(n_219),
.Y(n_3763)
);

BUFx6f_ASAP7_75t_L g3764 ( 
.A(n_3048),
.Y(n_3764)
);

CKINVDCx5p33_ASAP7_75t_R g3765 ( 
.A(n_3269),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3041),
.Y(n_3766)
);

O2A1O1Ixp5_ASAP7_75t_L g3767 ( 
.A1(n_2911),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3287),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_SL g3769 ( 
.A1(n_3055),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_3769)
);

BUFx6f_ASAP7_75t_L g3770 ( 
.A(n_3048),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3055),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3126),
.B(n_3129),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3098),
.Y(n_3773)
);

OR2x6_ASAP7_75t_L g3774 ( 
.A(n_3259),
.B(n_2694),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3287),
.Y(n_3775)
);

NOR2x1_ASAP7_75t_L g3776 ( 
.A(n_3207),
.B(n_222),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3151),
.Y(n_3777)
);

BUFx3_ASAP7_75t_L g3778 ( 
.A(n_2863),
.Y(n_3778)
);

INVxp67_ASAP7_75t_SL g3779 ( 
.A(n_2876),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3016),
.Y(n_3780)
);

NOR2xp33_ASAP7_75t_L g3781 ( 
.A(n_2807),
.B(n_223),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3136),
.B(n_224),
.Y(n_3782)
);

NOR2x2_ASAP7_75t_L g3783 ( 
.A(n_3218),
.B(n_225),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3156),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_3022),
.Y(n_3785)
);

AND2x4_ASAP7_75t_L g3786 ( 
.A(n_3028),
.B(n_224),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_SL g3787 ( 
.A(n_3039),
.B(n_589),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3030),
.Y(n_3788)
);

AND2x4_ASAP7_75t_L g3789 ( 
.A(n_3033),
.B(n_224),
.Y(n_3789)
);

CKINVDCx5p33_ASAP7_75t_R g3790 ( 
.A(n_2881),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_SL g3791 ( 
.A(n_2936),
.B(n_590),
.Y(n_3791)
);

BUFx3_ASAP7_75t_L g3792 ( 
.A(n_2866),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_2957),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_2818),
.B(n_2767),
.Y(n_3794)
);

INVx2_ASAP7_75t_SL g3795 ( 
.A(n_2711),
.Y(n_3795)
);

OAI22xp5_ASAP7_75t_SL g3796 ( 
.A1(n_3157),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_3796)
);

A2O1A1Ixp33_ASAP7_75t_L g3797 ( 
.A1(n_3014),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_3797)
);

OAI22xp5_ASAP7_75t_SL g3798 ( 
.A1(n_3159),
.A2(n_229),
.B1(n_226),
.B2(n_228),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3182),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3185),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3146),
.B(n_3168),
.Y(n_3801)
);

AND2x4_ASAP7_75t_L g3802 ( 
.A(n_3034),
.B(n_228),
.Y(n_3802)
);

AND2x4_ASAP7_75t_L g3803 ( 
.A(n_3034),
.B(n_229),
.Y(n_3803)
);

BUFx2_ASAP7_75t_L g3804 ( 
.A(n_2972),
.Y(n_3804)
);

BUFx2_ASAP7_75t_L g3805 ( 
.A(n_2980),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3184),
.B(n_229),
.Y(n_3806)
);

BUFx3_ASAP7_75t_L g3807 ( 
.A(n_2974),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3265),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_2973),
.Y(n_3809)
);

AND2x4_ASAP7_75t_L g3810 ( 
.A(n_2989),
.B(n_230),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_2954),
.Y(n_3811)
);

AOI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_2651),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_3812)
);

INVxp67_ASAP7_75t_L g3813 ( 
.A(n_3224),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_L g3814 ( 
.A(n_2767),
.B(n_230),
.Y(n_3814)
);

AOI22x1_ASAP7_75t_L g3815 ( 
.A1(n_2814),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3815)
);

BUFx2_ASAP7_75t_L g3816 ( 
.A(n_2814),
.Y(n_3816)
);

NOR3xp33_ASAP7_75t_SL g3817 ( 
.A(n_3069),
.B(n_231),
.C(n_233),
.Y(n_3817)
);

INVx2_ASAP7_75t_SL g3818 ( 
.A(n_2827),
.Y(n_3818)
);

INVx3_ASAP7_75t_L g3819 ( 
.A(n_2839),
.Y(n_3819)
);

AOI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3237),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_3820)
);

AOI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_2905),
.A2(n_234),
.B(n_235),
.Y(n_3821)
);

BUFx3_ASAP7_75t_L g3822 ( 
.A(n_2839),
.Y(n_3822)
);

INVx2_ASAP7_75t_SL g3823 ( 
.A(n_2724),
.Y(n_3823)
);

O2A1O1Ixp33_ASAP7_75t_L g3824 ( 
.A1(n_3072),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_3824)
);

BUFx6f_ASAP7_75t_L g3825 ( 
.A(n_3048),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_2954),
.Y(n_3826)
);

BUFx6f_ASAP7_75t_L g3827 ( 
.A(n_2920),
.Y(n_3827)
);

INVx2_ASAP7_75t_SL g3828 ( 
.A(n_2785),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3253),
.B(n_236),
.Y(n_3829)
);

NOR2xp33_ASAP7_75t_L g3830 ( 
.A(n_2798),
.B(n_236),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_SL g3831 ( 
.A(n_2865),
.B(n_590),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_2960),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3266),
.B(n_237),
.Y(n_3833)
);

AOI22xp5_ASAP7_75t_L g3834 ( 
.A1(n_3288),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_2798),
.B(n_237),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_2865),
.B(n_238),
.Y(n_3836)
);

BUFx3_ASAP7_75t_L g3837 ( 
.A(n_3015),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_SL g3838 ( 
.A(n_3189),
.B(n_592),
.Y(n_3838)
);

OAI22xp5_ASAP7_75t_L g3839 ( 
.A1(n_3159),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_2846),
.B(n_241),
.Y(n_3840)
);

NOR2xp33_ASAP7_75t_R g3841 ( 
.A(n_2893),
.B(n_242),
.Y(n_3841)
);

AND2x2_ASAP7_75t_SL g3842 ( 
.A(n_3273),
.B(n_243),
.Y(n_3842)
);

BUFx3_ASAP7_75t_L g3843 ( 
.A(n_2949),
.Y(n_3843)
);

BUFx6f_ASAP7_75t_L g3844 ( 
.A(n_2930),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_2960),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_2909),
.Y(n_3846)
);

BUFx6f_ASAP7_75t_L g3847 ( 
.A(n_2961),
.Y(n_3847)
);

NAND2x1p5_ASAP7_75t_L g3848 ( 
.A(n_2853),
.B(n_243),
.Y(n_3848)
);

NOR2x2_ASAP7_75t_L g3849 ( 
.A(n_2825),
.B(n_244),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_2799),
.B(n_243),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3337),
.B(n_3193),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3811),
.B(n_3273),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_SL g3853 ( 
.A(n_3384),
.B(n_3580),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3651),
.B(n_3193),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3613),
.B(n_3291),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_SL g3856 ( 
.A(n_3391),
.B(n_3291),
.Y(n_3856)
);

NAND2xp33_ASAP7_75t_SL g3857 ( 
.A(n_3640),
.B(n_2970),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3391),
.B(n_3029),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3476),
.B(n_2664),
.Y(n_3859)
);

AND2x4_ASAP7_75t_L g3860 ( 
.A(n_3615),
.B(n_2837),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_SL g3861 ( 
.A(n_3737),
.B(n_3031),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3826),
.B(n_3139),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_SL g3863 ( 
.A(n_3842),
.B(n_2805),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_SL g3864 ( 
.A(n_3616),
.B(n_2805),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3790),
.B(n_3230),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_3631),
.B(n_3258),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3432),
.B(n_3488),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_SL g3868 ( 
.A(n_3488),
.B(n_2745),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3494),
.B(n_2799),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3556),
.B(n_2975),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3301),
.B(n_2806),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_SL g3872 ( 
.A(n_3306),
.B(n_3000),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_SL g3873 ( 
.A(n_3663),
.B(n_3000),
.Y(n_3873)
);

NOR2xp33_ASAP7_75t_SL g3874 ( 
.A(n_3300),
.B(n_3388),
.Y(n_3874)
);

AND2x4_ASAP7_75t_L g3875 ( 
.A(n_3621),
.B(n_2962),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_SL g3876 ( 
.A(n_3663),
.B(n_2971),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_SL g3877 ( 
.A(n_3663),
.B(n_3049),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_3728),
.B(n_3272),
.Y(n_3878)
);

NAND2xp33_ASAP7_75t_SL g3879 ( 
.A(n_3573),
.B(n_2990),
.Y(n_3879)
);

NAND2xp33_ASAP7_75t_SL g3880 ( 
.A(n_3841),
.B(n_2967),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_SL g3881 ( 
.A(n_3731),
.B(n_3426),
.Y(n_3881)
);

NAND2xp33_ASAP7_75t_SL g3882 ( 
.A(n_3699),
.B(n_3082),
.Y(n_3882)
);

NAND2xp33_ASAP7_75t_SL g3883 ( 
.A(n_3687),
.B(n_3399),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_SL g3884 ( 
.A(n_3426),
.B(n_3130),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_3426),
.B(n_3138),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_SL g3886 ( 
.A(n_3816),
.B(n_3143),
.Y(n_3886)
);

NAND2xp33_ASAP7_75t_SL g3887 ( 
.A(n_3689),
.B(n_3094),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_SL g3888 ( 
.A(n_3310),
.B(n_3181),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3794),
.B(n_2806),
.Y(n_3889)
);

NAND2xp33_ASAP7_75t_SL g3890 ( 
.A(n_3817),
.B(n_3112),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3478),
.B(n_3201),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3478),
.B(n_3204),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3501),
.B(n_3216),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_SL g3894 ( 
.A(n_3566),
.B(n_3231),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_SL g3895 ( 
.A(n_3417),
.B(n_3267),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_SL g3896 ( 
.A(n_3305),
.B(n_3268),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_SL g3897 ( 
.A(n_3305),
.B(n_3125),
.Y(n_3897)
);

XNOR2x2_ASAP7_75t_L g3898 ( 
.A(n_3378),
.B(n_3161),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3832),
.B(n_2816),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_SL g3900 ( 
.A(n_3333),
.B(n_3194),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_SL g3901 ( 
.A(n_3333),
.B(n_3199),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_3335),
.B(n_3051),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_SL g3903 ( 
.A(n_3335),
.B(n_3047),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_3340),
.B(n_2997),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_3340),
.B(n_3007),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_SL g3906 ( 
.A(n_3347),
.B(n_2982),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3845),
.B(n_3387),
.Y(n_3907)
);

NAND2xp33_ASAP7_75t_SL g3908 ( 
.A(n_3365),
.B(n_3796),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_3347),
.B(n_2856),
.Y(n_3909)
);

NAND2xp33_ASAP7_75t_SL g3910 ( 
.A(n_3798),
.B(n_3038),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_SL g3911 ( 
.A(n_3359),
.B(n_2816),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_SL g3912 ( 
.A(n_3359),
.B(n_2855),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_SL g3913 ( 
.A(n_3589),
.B(n_3045),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_SL g3914 ( 
.A(n_3470),
.B(n_2909),
.Y(n_3914)
);

AND2x4_ASAP7_75t_L g3915 ( 
.A(n_3621),
.B(n_3005),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_SL g3916 ( 
.A(n_3520),
.B(n_3050),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3520),
.B(n_2758),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_SL g3918 ( 
.A(n_3430),
.B(n_2758),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_SL g3919 ( 
.A(n_3304),
.B(n_2965),
.Y(n_3919)
);

NAND2xp33_ASAP7_75t_SL g3920 ( 
.A(n_3385),
.B(n_3013),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_SL g3921 ( 
.A(n_3769),
.B(n_3298),
.Y(n_3921)
);

NAND2xp33_ASAP7_75t_SL g3922 ( 
.A(n_3357),
.B(n_3011),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_SL g3923 ( 
.A(n_3298),
.B(n_2854),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3298),
.B(n_2864),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3405),
.B(n_2858),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_SL g3926 ( 
.A(n_3379),
.B(n_2743),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3388),
.B(n_3420),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_SL g3928 ( 
.A(n_3379),
.B(n_2746),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_SL g3929 ( 
.A(n_3379),
.B(n_2752),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_3394),
.B(n_2993),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_SL g3931 ( 
.A(n_3394),
.B(n_2771),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_3394),
.B(n_2780),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_SL g3933 ( 
.A(n_3401),
.B(n_2720),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_SL g3934 ( 
.A(n_3401),
.B(n_2859),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_SL g3935 ( 
.A(n_3401),
.B(n_2861),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_SL g3936 ( 
.A(n_3413),
.B(n_3538),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3489),
.B(n_2870),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3420),
.B(n_2793),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3413),
.B(n_2868),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_SL g3940 ( 
.A(n_3413),
.B(n_2857),
.Y(n_3940)
);

NAND2xp33_ASAP7_75t_SL g3941 ( 
.A(n_3397),
.B(n_3025),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3657),
.B(n_2894),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_SL g3943 ( 
.A(n_3538),
.B(n_2857),
.Y(n_3943)
);

NAND2xp33_ASAP7_75t_SL g3944 ( 
.A(n_3449),
.B(n_2862),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_SL g3945 ( 
.A(n_3538),
.B(n_2955),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3850),
.B(n_2795),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3541),
.B(n_2950),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3598),
.B(n_2654),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_SL g3949 ( 
.A(n_3541),
.B(n_3546),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_SL g3950 ( 
.A(n_3541),
.B(n_2994),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3546),
.B(n_3587),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3569),
.B(n_2845),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_SL g3953 ( 
.A(n_3546),
.B(n_2996),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3380),
.B(n_2877),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_SL g3955 ( 
.A(n_3587),
.B(n_2998),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3381),
.B(n_2880),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3315),
.B(n_2995),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_SL g3958 ( 
.A(n_3604),
.B(n_2940),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3383),
.B(n_2834),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_3604),
.B(n_2914),
.Y(n_3960)
);

NAND2xp33_ASAP7_75t_SL g3961 ( 
.A(n_3629),
.B(n_3551),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3810),
.B(n_2740),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3810),
.B(n_2883),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_SL g3964 ( 
.A(n_3802),
.B(n_2749),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3802),
.B(n_2649),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_SL g3966 ( 
.A(n_3803),
.B(n_2757),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_SL g3967 ( 
.A(n_3803),
.B(n_3646),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3646),
.B(n_2770),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3646),
.B(n_2783),
.Y(n_3969)
);

NAND2xp33_ASAP7_75t_SL g3970 ( 
.A(n_3629),
.B(n_2964),
.Y(n_3970)
);

NAND2xp33_ASAP7_75t_SL g3971 ( 
.A(n_3551),
.B(n_2956),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_SL g3972 ( 
.A(n_3533),
.B(n_3571),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_SL g3973 ( 
.A(n_3533),
.B(n_3571),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_SL g3974 ( 
.A(n_3730),
.B(n_2823),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3402),
.B(n_2847),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3460),
.B(n_3461),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3485),
.B(n_2790),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_SL g3978 ( 
.A(n_3485),
.B(n_2819),
.Y(n_3978)
);

NAND2xp33_ASAP7_75t_SL g3979 ( 
.A(n_3551),
.B(n_2723),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3456),
.B(n_2820),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_SL g3981 ( 
.A(n_3549),
.B(n_2822),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_SL g3982 ( 
.A(n_3564),
.B(n_2753),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_SL g3983 ( 
.A(n_3807),
.B(n_2849),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_SL g3984 ( 
.A(n_3491),
.B(n_2850),
.Y(n_3984)
);

XNOR2x2_ASAP7_75t_L g3985 ( 
.A(n_3739),
.B(n_2748),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3407),
.B(n_2869),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_SL g3987 ( 
.A(n_3837),
.B(n_2661),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3408),
.B(n_3409),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_SL g3989 ( 
.A(n_3373),
.B(n_2665),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_SL g3990 ( 
.A(n_3614),
.B(n_2676),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_3614),
.B(n_2677),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_3656),
.B(n_2681),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_3656),
.B(n_2697),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3414),
.B(n_2884),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_SL g3995 ( 
.A(n_3685),
.B(n_2699),
.Y(n_3995)
);

NAND2xp33_ASAP7_75t_L g3996 ( 
.A(n_3487),
.B(n_2700),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_SL g3997 ( 
.A(n_3685),
.B(n_2712),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_SL g3998 ( 
.A(n_3736),
.B(n_2727),
.Y(n_3998)
);

AND2x4_ASAP7_75t_L g3999 ( 
.A(n_3465),
.B(n_3010),
.Y(n_3999)
);

NAND2xp33_ASAP7_75t_SL g4000 ( 
.A(n_3597),
.B(n_2804),
.Y(n_4000)
);

NAND2xp33_ASAP7_75t_SL g4001 ( 
.A(n_3597),
.B(n_2750),
.Y(n_4001)
);

NAND2xp33_ASAP7_75t_SL g4002 ( 
.A(n_3597),
.B(n_2775),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3736),
.B(n_2728),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_SL g4004 ( 
.A(n_3746),
.B(n_2948),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3746),
.B(n_2923),
.Y(n_4005)
);

NOR2xp33_ASAP7_75t_L g4006 ( 
.A(n_3813),
.B(n_2945),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_SL g4007 ( 
.A(n_3750),
.B(n_2907),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3750),
.B(n_3822),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_SL g4009 ( 
.A(n_3447),
.B(n_2784),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3557),
.B(n_2912),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_SL g4011 ( 
.A(n_3467),
.B(n_2867),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_SL g4012 ( 
.A(n_3819),
.B(n_2899),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_SL g4013 ( 
.A(n_3343),
.B(n_2904),
.Y(n_4013)
);

NAND2xp33_ASAP7_75t_SL g4014 ( 
.A(n_3427),
.B(n_3425),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_SL g4015 ( 
.A(n_3698),
.B(n_2947),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_SL g4016 ( 
.A(n_3706),
.B(n_2919),
.Y(n_4016)
);

NAND2xp33_ASAP7_75t_SL g4017 ( 
.A(n_3555),
.B(n_2809),
.Y(n_4017)
);

NAND2xp33_ASAP7_75t_SL g4018 ( 
.A(n_3334),
.B(n_2929),
.Y(n_4018)
);

NAND2xp33_ASAP7_75t_SL g4019 ( 
.A(n_3752),
.B(n_2932),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3415),
.B(n_2944),
.Y(n_4020)
);

NAND2xp33_ASAP7_75t_SL g4021 ( 
.A(n_3839),
.B(n_244),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_3584),
.B(n_245),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3416),
.B(n_245),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_SL g4024 ( 
.A(n_3600),
.B(n_245),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3422),
.B(n_246),
.Y(n_4025)
);

NAND2xp33_ASAP7_75t_SL g4026 ( 
.A(n_3392),
.B(n_246),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_SL g4027 ( 
.A(n_3818),
.B(n_246),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_SL g4028 ( 
.A(n_3693),
.B(n_247),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3579),
.B(n_247),
.Y(n_4029)
);

AND2x2_ASAP7_75t_SL g4030 ( 
.A(n_3314),
.B(n_247),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_SL g4031 ( 
.A(n_3344),
.B(n_248),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_SL g4032 ( 
.A(n_3468),
.B(n_248),
.Y(n_4032)
);

NAND2xp33_ASAP7_75t_SL g4033 ( 
.A(n_3341),
.B(n_249),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_SL g4034 ( 
.A(n_3486),
.B(n_249),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_SL g4035 ( 
.A(n_3745),
.B(n_249),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_SL g4036 ( 
.A(n_3499),
.B(n_3717),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_3827),
.B(n_250),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3439),
.B(n_250),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3827),
.B(n_251),
.Y(n_4039)
);

NAND2xp33_ASAP7_75t_SL g4040 ( 
.A(n_3299),
.B(n_251),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3827),
.B(n_251),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3443),
.B(n_252),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_SL g4043 ( 
.A(n_3844),
.B(n_252),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_3844),
.B(n_252),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3444),
.B(n_254),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_SL g4046 ( 
.A(n_3844),
.B(n_254),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_SL g4047 ( 
.A(n_3847),
.B(n_254),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_SL g4048 ( 
.A(n_3847),
.B(n_255),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_SL g4049 ( 
.A(n_3847),
.B(n_255),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_SL g4050 ( 
.A(n_3545),
.B(n_256),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_SL g4051 ( 
.A(n_3776),
.B(n_257),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_SL g4052 ( 
.A(n_3765),
.B(n_257),
.Y(n_4052)
);

NAND2xp33_ASAP7_75t_SL g4053 ( 
.A(n_3303),
.B(n_3692),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_SL g4054 ( 
.A(n_3697),
.B(n_257),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3453),
.B(n_258),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3697),
.B(n_259),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_SL g4057 ( 
.A(n_3697),
.B(n_259),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3463),
.B(n_259),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_3722),
.B(n_260),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3466),
.B(n_3472),
.Y(n_4060)
);

AND2x2_ASAP7_75t_SL g4061 ( 
.A(n_3771),
.B(n_260),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_SL g4062 ( 
.A(n_3722),
.B(n_261),
.Y(n_4062)
);

NAND2xp33_ASAP7_75t_SL g4063 ( 
.A(n_3543),
.B(n_261),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_SL g4064 ( 
.A(n_3722),
.B(n_261),
.Y(n_4064)
);

NAND2xp33_ASAP7_75t_SL g4065 ( 
.A(n_3575),
.B(n_262),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_SL g4066 ( 
.A(n_3757),
.B(n_262),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_SL g4067 ( 
.A(n_3757),
.B(n_262),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_SL g4068 ( 
.A(n_3757),
.B(n_263),
.Y(n_4068)
);

NAND2xp33_ASAP7_75t_SL g4069 ( 
.A(n_3327),
.B(n_263),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_SL g4070 ( 
.A(n_3758),
.B(n_3374),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_3758),
.B(n_263),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3479),
.B(n_264),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_SL g4073 ( 
.A(n_3758),
.B(n_264),
.Y(n_4073)
);

NAND2xp33_ASAP7_75t_SL g4074 ( 
.A(n_3351),
.B(n_264),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_SL g4075 ( 
.A(n_3297),
.B(n_265),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_SL g4076 ( 
.A(n_3644),
.B(n_265),
.Y(n_4076)
);

NAND2xp33_ASAP7_75t_SL g4077 ( 
.A(n_3487),
.B(n_266),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_SL g4078 ( 
.A(n_3741),
.B(n_3786),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_SL g4079 ( 
.A(n_3786),
.B(n_266),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_3789),
.B(n_3595),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3480),
.B(n_267),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_SL g4082 ( 
.A(n_3789),
.B(n_267),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_3617),
.B(n_267),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_SL g4084 ( 
.A(n_3464),
.B(n_268),
.Y(n_4084)
);

NAND2xp33_ASAP7_75t_SL g4085 ( 
.A(n_3574),
.B(n_268),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_SL g4086 ( 
.A(n_3764),
.B(n_269),
.Y(n_4086)
);

NAND2xp33_ASAP7_75t_SL g4087 ( 
.A(n_3358),
.B(n_3361),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_SL g4088 ( 
.A(n_3764),
.B(n_269),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_SL g4089 ( 
.A(n_3764),
.B(n_3770),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3490),
.B(n_269),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_SL g4091 ( 
.A(n_3770),
.B(n_270),
.Y(n_4091)
);

NAND2xp33_ASAP7_75t_SL g4092 ( 
.A(n_3292),
.B(n_270),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_SL g4093 ( 
.A(n_3770),
.B(n_270),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_SL g4094 ( 
.A(n_3825),
.B(n_271),
.Y(n_4094)
);

NAND2xp33_ASAP7_75t_SL g4095 ( 
.A(n_3367),
.B(n_271),
.Y(n_4095)
);

NAND2xp33_ASAP7_75t_SL g4096 ( 
.A(n_3377),
.B(n_271),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_SL g4097 ( 
.A(n_3825),
.B(n_3753),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_SL g4098 ( 
.A(n_3825),
.B(n_3410),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_SL g4099 ( 
.A(n_3446),
.B(n_272),
.Y(n_4099)
);

NAND2xp33_ASAP7_75t_SL g4100 ( 
.A(n_3602),
.B(n_273),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_SL g4101 ( 
.A(n_3462),
.B(n_3469),
.Y(n_4101)
);

NAND2xp33_ASAP7_75t_SL g4102 ( 
.A(n_3592),
.B(n_273),
.Y(n_4102)
);

NAND2xp33_ASAP7_75t_SL g4103 ( 
.A(n_3831),
.B(n_3836),
.Y(n_4103)
);

NAND2xp33_ASAP7_75t_SL g4104 ( 
.A(n_3726),
.B(n_274),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_SL g4105 ( 
.A(n_3369),
.B(n_3505),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_SL g4106 ( 
.A(n_3506),
.B(n_274),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_SL g4107 ( 
.A(n_3527),
.B(n_274),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_SL g4108 ( 
.A(n_3321),
.B(n_275),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_SL g4109 ( 
.A(n_3779),
.B(n_276),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_SL g4110 ( 
.A(n_3848),
.B(n_276),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_3411),
.B(n_277),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_SL g4112 ( 
.A(n_3668),
.B(n_278),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_SL g4113 ( 
.A(n_3669),
.B(n_278),
.Y(n_4113)
);

NAND2xp33_ASAP7_75t_L g4114 ( 
.A(n_3540),
.B(n_278),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_SL g4115 ( 
.A(n_3703),
.B(n_279),
.Y(n_4115)
);

NAND2xp33_ASAP7_75t_SL g4116 ( 
.A(n_3322),
.B(n_279),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_3704),
.B(n_3710),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_SL g4118 ( 
.A(n_3686),
.B(n_280),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_3581),
.B(n_280),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3630),
.B(n_280),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_SL g4121 ( 
.A(n_3642),
.B(n_281),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3496),
.B(n_281),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3510),
.B(n_282),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_3511),
.B(n_3749),
.Y(n_4124)
);

NAND2xp33_ASAP7_75t_SL g4125 ( 
.A(n_3611),
.B(n_282),
.Y(n_4125)
);

NAND2xp33_ASAP7_75t_SL g4126 ( 
.A(n_3838),
.B(n_283),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_SL g4127 ( 
.A(n_3809),
.B(n_283),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_SL g4128 ( 
.A(n_3452),
.B(n_283),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_SL g4129 ( 
.A(n_3458),
.B(n_284),
.Y(n_4129)
);

AND2x4_ASAP7_75t_L g4130 ( 
.A(n_3477),
.B(n_3481),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_SL g4131 ( 
.A(n_3498),
.B(n_284),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_SL g4132 ( 
.A(n_3504),
.B(n_3529),
.Y(n_4132)
);

NAND2xp33_ASAP7_75t_SL g4133 ( 
.A(n_3568),
.B(n_285),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_3386),
.B(n_285),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_SL g4135 ( 
.A(n_3846),
.B(n_285),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_SL g4136 ( 
.A(n_3560),
.B(n_286),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3516),
.B(n_3517),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_SL g4138 ( 
.A(n_3576),
.B(n_286),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_SL g4139 ( 
.A(n_3332),
.B(n_286),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_SL g4140 ( 
.A(n_3352),
.B(n_287),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_SL g4141 ( 
.A(n_3804),
.B(n_287),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_SL g4142 ( 
.A(n_3805),
.B(n_287),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_SL g4143 ( 
.A(n_3815),
.B(n_288),
.Y(n_4143)
);

AND2x2_ASAP7_75t_L g4144 ( 
.A(n_3404),
.B(n_288),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_SL g4145 ( 
.A(n_3502),
.B(n_288),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3526),
.B(n_289),
.Y(n_4146)
);

NAND2xp33_ASAP7_75t_SL g4147 ( 
.A(n_3583),
.B(n_289),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_SL g4148 ( 
.A(n_3535),
.B(n_290),
.Y(n_4148)
);

NAND2xp33_ASAP7_75t_SL g4149 ( 
.A(n_3591),
.B(n_3715),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_SL g4150 ( 
.A(n_3547),
.B(n_291),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3773),
.B(n_291),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_SL g4152 ( 
.A(n_3777),
.B(n_292),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_SL g4153 ( 
.A(n_3784),
.B(n_292),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_SL g4154 ( 
.A(n_3799),
.B(n_292),
.Y(n_4154)
);

NAND2xp33_ASAP7_75t_SL g4155 ( 
.A(n_3787),
.B(n_293),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_SL g4156 ( 
.A(n_3800),
.B(n_293),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_SL g4157 ( 
.A(n_3808),
.B(n_3435),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_SL g4158 ( 
.A(n_3590),
.B(n_293),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_SL g4159 ( 
.A(n_3636),
.B(n_294),
.Y(n_4159)
);

NAND2xp33_ASAP7_75t_SL g4160 ( 
.A(n_3627),
.B(n_294),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_3659),
.B(n_294),
.Y(n_4161)
);

NAND2xp33_ASAP7_75t_SL g4162 ( 
.A(n_3634),
.B(n_295),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_SL g4163 ( 
.A(n_3720),
.B(n_295),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_SL g4164 ( 
.A(n_3725),
.B(n_295),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_SL g4165 ( 
.A(n_3672),
.B(n_296),
.Y(n_4165)
);

NAND2xp33_ASAP7_75t_SL g4166 ( 
.A(n_3635),
.B(n_296),
.Y(n_4166)
);

NAND2xp33_ASAP7_75t_SL g4167 ( 
.A(n_3524),
.B(n_297),
.Y(n_4167)
);

NAND2xp33_ASAP7_75t_SL g4168 ( 
.A(n_3791),
.B(n_298),
.Y(n_4168)
);

NAND2xp33_ASAP7_75t_SL g4169 ( 
.A(n_3320),
.B(n_298),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3528),
.B(n_298),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_SL g4171 ( 
.A(n_3530),
.B(n_299),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_3542),
.B(n_299),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3550),
.B(n_299),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_SL g4174 ( 
.A(n_3552),
.B(n_300),
.Y(n_4174)
);

NAND2xp33_ASAP7_75t_SL g4175 ( 
.A(n_3350),
.B(n_300),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_SL g4176 ( 
.A(n_3558),
.B(n_301),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_SL g4177 ( 
.A(n_3563),
.B(n_3567),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3582),
.B(n_301),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_3302),
.B(n_302),
.Y(n_4179)
);

NAND2xp33_ASAP7_75t_SL g4180 ( 
.A(n_3436),
.B(n_302),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_SL g4181 ( 
.A(n_3593),
.B(n_302),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_SL g4182 ( 
.A(n_3594),
.B(n_303),
.Y(n_4182)
);

NAND2xp33_ASAP7_75t_SL g4183 ( 
.A(n_3534),
.B(n_303),
.Y(n_4183)
);

NAND2xp33_ASAP7_75t_SL g4184 ( 
.A(n_3534),
.B(n_303),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_SL g4185 ( 
.A(n_3607),
.B(n_304),
.Y(n_4185)
);

NAND2xp33_ASAP7_75t_SL g4186 ( 
.A(n_3577),
.B(n_304),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_SL g4187 ( 
.A(n_3608),
.B(n_304),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_SL g4188 ( 
.A(n_3609),
.B(n_305),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_3618),
.B(n_305),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_SL g4190 ( 
.A(n_3619),
.B(n_305),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_3620),
.B(n_3623),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_SL g4192 ( 
.A(n_3624),
.B(n_3633),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_SL g4193 ( 
.A(n_3641),
.B(n_306),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_SL g4194 ( 
.A(n_3643),
.B(n_306),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_SL g4195 ( 
.A(n_3645),
.B(n_3650),
.Y(n_4195)
);

NAND2xp33_ASAP7_75t_SL g4196 ( 
.A(n_3441),
.B(n_306),
.Y(n_4196)
);

NAND2xp33_ASAP7_75t_SL g4197 ( 
.A(n_3539),
.B(n_307),
.Y(n_4197)
);

AND2x4_ASAP7_75t_L g4198 ( 
.A(n_3403),
.B(n_3406),
.Y(n_4198)
);

NAND2xp33_ASAP7_75t_SL g4199 ( 
.A(n_3578),
.B(n_307),
.Y(n_4199)
);

NAND2xp33_ASAP7_75t_SL g4200 ( 
.A(n_3455),
.B(n_307),
.Y(n_4200)
);

XNOR2xp5_ASAP7_75t_L g4201 ( 
.A(n_3497),
.B(n_308),
.Y(n_4201)
);

NAND2xp33_ASAP7_75t_SL g4202 ( 
.A(n_3474),
.B(n_308),
.Y(n_4202)
);

NAND2xp33_ASAP7_75t_SL g4203 ( 
.A(n_3482),
.B(n_309),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3654),
.B(n_309),
.Y(n_4204)
);

NAND2xp33_ASAP7_75t_SL g4205 ( 
.A(n_3531),
.B(n_309),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_SL g4206 ( 
.A(n_3673),
.B(n_310),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3677),
.B(n_3679),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_SL g4208 ( 
.A(n_3680),
.B(n_310),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_SL g4209 ( 
.A(n_3690),
.B(n_310),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_SL g4210 ( 
.A(n_3694),
.B(n_311),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_SL g4211 ( 
.A(n_3695),
.B(n_311),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_SL g4212 ( 
.A(n_3700),
.B(n_312),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_3713),
.B(n_312),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_SL g4214 ( 
.A(n_3714),
.B(n_313),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_SL g4215 ( 
.A(n_3716),
.B(n_313),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_SL g4216 ( 
.A(n_3724),
.B(n_314),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_3325),
.B(n_314),
.Y(n_4217)
);

NAND2xp33_ASAP7_75t_SL g4218 ( 
.A(n_3628),
.B(n_314),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_3732),
.B(n_315),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_SL g4220 ( 
.A(n_3754),
.B(n_315),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_3814),
.B(n_316),
.Y(n_4221)
);

AND2x4_ASAP7_75t_L g4222 ( 
.A(n_3484),
.B(n_316),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_3780),
.B(n_316),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_SL g4224 ( 
.A(n_3785),
.B(n_317),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_SL g4225 ( 
.A(n_3788),
.B(n_317),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_3308),
.B(n_317),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_SL g4227 ( 
.A(n_3681),
.B(n_318),
.Y(n_4227)
);

NAND2xp33_ASAP7_75t_SL g4228 ( 
.A(n_3684),
.B(n_318),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_SL g4229 ( 
.A(n_3830),
.B(n_3835),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_3766),
.B(n_319),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_SL g4231 ( 
.A(n_3781),
.B(n_319),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_3601),
.B(n_319),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_SL g4233 ( 
.A(n_3655),
.B(n_320),
.Y(n_4233)
);

AND2x4_ASAP7_75t_L g4234 ( 
.A(n_3493),
.B(n_320),
.Y(n_4234)
);

NAND2xp33_ASAP7_75t_SL g4235 ( 
.A(n_3647),
.B(n_320),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_SL g4236 ( 
.A(n_3721),
.B(n_321),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_SL g4237 ( 
.A(n_3395),
.B(n_321),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_SL g4238 ( 
.A(n_3328),
.B(n_321),
.Y(n_4238)
);

NAND2xp33_ASAP7_75t_SL g4239 ( 
.A(n_3424),
.B(n_322),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_SL g4240 ( 
.A(n_3738),
.B(n_322),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_SL g4241 ( 
.A(n_3658),
.B(n_323),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_SL g4242 ( 
.A(n_3661),
.B(n_323),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_SL g4243 ( 
.A(n_3653),
.B(n_323),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_3719),
.B(n_324),
.Y(n_4244)
);

AND2x4_ASAP7_75t_L g4245 ( 
.A(n_3605),
.B(n_324),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_SL g4246 ( 
.A(n_3707),
.B(n_325),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_3610),
.B(n_325),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_SL g4248 ( 
.A(n_3638),
.B(n_326),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_3612),
.B(n_3296),
.Y(n_4249)
);

NAND2xp33_ASAP7_75t_SL g4250 ( 
.A(n_3437),
.B(n_326),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_SL g4251 ( 
.A(n_3652),
.B(n_327),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_3688),
.B(n_327),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_SL g4253 ( 
.A(n_3366),
.B(n_328),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_SL g4254 ( 
.A(n_3326),
.B(n_328),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_SL g4255 ( 
.A(n_3772),
.B(n_328),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_SL g4256 ( 
.A(n_3801),
.B(n_329),
.Y(n_4256)
);

AND2x4_ASAP7_75t_L g4257 ( 
.A(n_3364),
.B(n_329),
.Y(n_4257)
);

NAND2xp33_ASAP7_75t_SL g4258 ( 
.A(n_3440),
.B(n_330),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_3330),
.B(n_330),
.Y(n_4259)
);

AND2x4_ASAP7_75t_L g4260 ( 
.A(n_3371),
.B(n_331),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_SL g4261 ( 
.A(n_3537),
.B(n_331),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_SL g4262 ( 
.A(n_3820),
.B(n_332),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_SL g4263 ( 
.A(n_3834),
.B(n_332),
.Y(n_4263)
);

NAND2xp33_ASAP7_75t_SL g4264 ( 
.A(n_3450),
.B(n_332),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_3331),
.B(n_333),
.Y(n_4265)
);

NAND2xp33_ASAP7_75t_SL g4266 ( 
.A(n_3473),
.B(n_333),
.Y(n_4266)
);

NAND2xp33_ASAP7_75t_SL g4267 ( 
.A(n_3475),
.B(n_333),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_SL g4268 ( 
.A(n_3588),
.B(n_334),
.Y(n_4268)
);

NAND2xp33_ASAP7_75t_SL g4269 ( 
.A(n_3500),
.B(n_334),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_SL g4270 ( 
.A(n_3797),
.B(n_334),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_SL g4271 ( 
.A(n_3824),
.B(n_3793),
.Y(n_4271)
);

AND2x4_ASAP7_75t_L g4272 ( 
.A(n_3293),
.B(n_335),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_SL g4273 ( 
.A(n_3348),
.B(n_335),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_3691),
.B(n_335),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_SL g4275 ( 
.A(n_3349),
.B(n_336),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_3353),
.B(n_336),
.Y(n_4276)
);

XNOR2xp5_ASAP7_75t_L g4277 ( 
.A(n_3316),
.B(n_337),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_3514),
.B(n_337),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_SL g4279 ( 
.A(n_3519),
.B(n_338),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_SL g4280 ( 
.A(n_3626),
.B(n_3712),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_SL g4281 ( 
.A(n_3762),
.B(n_338),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_3696),
.B(n_338),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_SL g4283 ( 
.A(n_3702),
.B(n_339),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_SL g4284 ( 
.A(n_3812),
.B(n_339),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_SL g4285 ( 
.A(n_3512),
.B(n_339),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_SL g4286 ( 
.A(n_3761),
.B(n_340),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_3751),
.B(n_340),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_3294),
.B(n_340),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_SL g4289 ( 
.A(n_3309),
.B(n_341),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_3311),
.B(n_341),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_SL g4291 ( 
.A(n_3313),
.B(n_342),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_SL g4292 ( 
.A(n_3319),
.B(n_342),
.Y(n_4292)
);

NAND2xp33_ASAP7_75t_SL g4293 ( 
.A(n_3445),
.B(n_3823),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_SL g4294 ( 
.A(n_3336),
.B(n_342),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_SL g4295 ( 
.A(n_3339),
.B(n_343),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_SL g4296 ( 
.A(n_3342),
.B(n_343),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_3907),
.B(n_3360),
.Y(n_4297)
);

INVx3_ASAP7_75t_L g4298 ( 
.A(n_3860),
.Y(n_4298)
);

NOR2xp67_ASAP7_75t_L g4299 ( 
.A(n_3927),
.B(n_3471),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4137),
.B(n_3363),
.Y(n_4300)
);

AOI22xp33_ASAP7_75t_L g4301 ( 
.A1(n_3910),
.A2(n_3676),
.B1(n_3540),
.B2(n_3318),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_3867),
.B(n_3760),
.Y(n_4302)
);

INVx3_ASAP7_75t_SL g4303 ( 
.A(n_4132),
.Y(n_4303)
);

OAI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_4226),
.A2(n_3866),
.B(n_3767),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4124),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_3976),
.B(n_3727),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_SL g4307 ( 
.A(n_3874),
.B(n_3570),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4198),
.Y(n_4308)
);

A2O1A1Ixp33_ASAP7_75t_L g4309 ( 
.A1(n_4183),
.A2(n_3398),
.B(n_3671),
.C(n_3662),
.Y(n_4309)
);

AOI22xp33_ASAP7_75t_L g4310 ( 
.A1(n_3883),
.A2(n_3676),
.B1(n_3540),
.B2(n_3760),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_SL g4311 ( 
.A(n_4030),
.B(n_3570),
.Y(n_4311)
);

CKINVDCx20_ASAP7_75t_R g4312 ( 
.A(n_4087),
.Y(n_4312)
);

BUFx8_ASAP7_75t_L g4313 ( 
.A(n_3938),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4198),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4198),
.Y(n_4315)
);

XOR2xp5_ASAP7_75t_L g4316 ( 
.A(n_4201),
.B(n_3346),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4207),
.B(n_3492),
.Y(n_4317)
);

CKINVDCx20_ASAP7_75t_R g4318 ( 
.A(n_4277),
.Y(n_4318)
);

INVx6_ASAP7_75t_L g4319 ( 
.A(n_3860),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4130),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3988),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4060),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4029),
.B(n_3622),
.Y(n_4323)
);

NOR2xp33_ASAP7_75t_L g4324 ( 
.A(n_3908),
.B(n_3429),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3899),
.B(n_3625),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4144),
.B(n_3637),
.Y(n_4326)
);

INVxp33_ASAP7_75t_L g4327 ( 
.A(n_3853),
.Y(n_4327)
);

AO22x1_ASAP7_75t_L g4328 ( 
.A1(n_4222),
.A2(n_3760),
.B1(n_3554),
.B2(n_3783),
.Y(n_4328)
);

INVxp67_ASAP7_75t_L g4329 ( 
.A(n_4036),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_3889),
.B(n_3666),
.Y(n_4330)
);

NOR2xp33_ASAP7_75t_L g4331 ( 
.A(n_4014),
.B(n_3649),
.Y(n_4331)
);

OR2x2_ASAP7_75t_L g4332 ( 
.A(n_4130),
.B(n_3843),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4222),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4177),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4222),
.Y(n_4335)
);

OAI21x1_ASAP7_75t_L g4336 ( 
.A1(n_4089),
.A2(n_3483),
.B(n_3821),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_4234),
.Y(n_4337)
);

OAI22xp5_ASAP7_75t_L g4338 ( 
.A1(n_4030),
.A2(n_3701),
.B1(n_3774),
.B2(n_3711),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4191),
.Y(n_4339)
);

OR2x2_ASAP7_75t_L g4340 ( 
.A(n_3942),
.B(n_3667),
.Y(n_4340)
);

BUFx6f_ASAP7_75t_L g4341 ( 
.A(n_3915),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_3869),
.B(n_3670),
.Y(n_4342)
);

AND2x2_ASAP7_75t_L g4343 ( 
.A(n_3957),
.B(n_3682),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_3859),
.B(n_3375),
.Y(n_4344)
);

BUFx2_ASAP7_75t_L g4345 ( 
.A(n_3970),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_4234),
.Y(n_4346)
);

OAI22xp5_ASAP7_75t_SL g4347 ( 
.A1(n_4061),
.A2(n_3774),
.B1(n_3660),
.B2(n_3849),
.Y(n_4347)
);

AOI22xp33_ASAP7_75t_L g4348 ( 
.A1(n_4053),
.A2(n_3733),
.B1(n_3572),
.B2(n_3718),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_3852),
.B(n_3312),
.Y(n_4349)
);

CKINVDCx5p33_ASAP7_75t_R g4350 ( 
.A(n_4180),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4010),
.B(n_3396),
.Y(n_4351)
);

BUFx3_ASAP7_75t_L g4352 ( 
.A(n_4272),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4192),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4234),
.Y(n_4354)
);

AND3x1_ASAP7_75t_SL g4355 ( 
.A(n_4184),
.B(n_3376),
.C(n_343),
.Y(n_4355)
);

OAI22xp5_ASAP7_75t_SL g4356 ( 
.A1(n_4061),
.A2(n_3423),
.B1(n_3307),
.B2(n_3412),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_3872),
.B(n_3317),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4195),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4272),
.B(n_3418),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_4249),
.B(n_3323),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_SL g4361 ( 
.A(n_3882),
.B(n_3400),
.Y(n_4361)
);

NAND2x1p5_ASAP7_75t_L g4362 ( 
.A(n_3967),
.B(n_3513),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4245),
.Y(n_4363)
);

BUFx6f_ASAP7_75t_L g4364 ( 
.A(n_3915),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4245),
.Y(n_4365)
);

CKINVDCx5p33_ASAP7_75t_R g4366 ( 
.A(n_4065),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_SL g4367 ( 
.A(n_4167),
.B(n_3795),
.Y(n_4367)
);

CKINVDCx5p33_ASAP7_75t_R g4368 ( 
.A(n_3920),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_3946),
.B(n_3324),
.Y(n_4369)
);

OAI22xp5_ASAP7_75t_L g4370 ( 
.A1(n_3861),
.A2(n_3747),
.B1(n_3755),
.B2(n_3743),
.Y(n_4370)
);

AOI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_4114),
.A2(n_3744),
.B1(n_3674),
.B2(n_3525),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_3862),
.B(n_3329),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4245),
.Y(n_4373)
);

INVx3_ASAP7_75t_L g4374 ( 
.A(n_3875),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4257),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4288),
.B(n_3419),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4290),
.B(n_3431),
.Y(n_4377)
);

BUFx3_ASAP7_75t_L g4378 ( 
.A(n_4257),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4257),
.Y(n_4379)
);

INVx2_ASAP7_75t_L g4380 ( 
.A(n_4260),
.Y(n_4380)
);

CKINVDCx20_ASAP7_75t_R g4381 ( 
.A(n_4293),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4179),
.Y(n_4382)
);

NOR2xp67_ASAP7_75t_L g4383 ( 
.A(n_3854),
.B(n_3828),
.Y(n_4383)
);

NOR2xp33_ASAP7_75t_SL g4384 ( 
.A(n_3875),
.B(n_3423),
.Y(n_4384)
);

BUFx6f_ASAP7_75t_L g4385 ( 
.A(n_3881),
.Y(n_4385)
);

HB1xp67_ASAP7_75t_L g4386 ( 
.A(n_4260),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_3871),
.B(n_3338),
.Y(n_4387)
);

NOR2xp67_ASAP7_75t_L g4388 ( 
.A(n_4157),
.B(n_3495),
.Y(n_4388)
);

BUFx3_ASAP7_75t_L g4389 ( 
.A(n_4260),
.Y(n_4389)
);

OR2x2_ASAP7_75t_L g4390 ( 
.A(n_4105),
.B(n_3433),
.Y(n_4390)
);

INVx2_ASAP7_75t_SL g4391 ( 
.A(n_4008),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4217),
.Y(n_4392)
);

CKINVDCx5p33_ASAP7_75t_R g4393 ( 
.A(n_4092),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_3922),
.Y(n_4394)
);

BUFx6f_ASAP7_75t_L g4395 ( 
.A(n_3951),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4259),
.Y(n_4396)
);

A2O1A1Ixp33_ASAP7_75t_L g4397 ( 
.A1(n_4160),
.A2(n_3683),
.B(n_3559),
.C(n_3544),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_3999),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4265),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_3954),
.B(n_3956),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4006),
.B(n_3434),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4006),
.B(n_3438),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_3959),
.B(n_3345),
.Y(n_4403)
);

BUFx4f_ASAP7_75t_L g4404 ( 
.A(n_3999),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_3972),
.B(n_3442),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4023),
.Y(n_4406)
);

AOI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_3880),
.A2(n_3740),
.B1(n_3515),
.B2(n_3561),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_SL g4408 ( 
.A(n_4149),
.B(n_3763),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_4020),
.Y(n_4409)
);

OAI22xp5_ASAP7_75t_SL g4410 ( 
.A1(n_4221),
.A2(n_3792),
.B1(n_3778),
.B2(n_3553),
.Y(n_4410)
);

BUFx3_ASAP7_75t_L g4411 ( 
.A(n_3948),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4247),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_3973),
.B(n_3983),
.Y(n_4413)
);

AND3x1_ASAP7_75t_SL g4414 ( 
.A(n_3941),
.B(n_344),
.C(n_345),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_3984),
.B(n_3448),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4274),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4025),
.Y(n_4417)
);

NAND2x1p5_ASAP7_75t_L g4418 ( 
.A(n_3855),
.B(n_3878),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_3975),
.B(n_3354),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_3987),
.B(n_3454),
.Y(n_4420)
);

OAI21x1_ASAP7_75t_L g4421 ( 
.A1(n_3936),
.A2(n_3768),
.B(n_3759),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4038),
.Y(n_4422)
);

INVx3_ASAP7_75t_L g4423 ( 
.A(n_3898),
.Y(n_4423)
);

AND3x1_ASAP7_75t_SL g4424 ( 
.A(n_3857),
.B(n_344),
.C(n_345),
.Y(n_4424)
);

INVx3_ASAP7_75t_L g4425 ( 
.A(n_3985),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_3986),
.B(n_3355),
.Y(n_4426)
);

BUFx3_ASAP7_75t_L g4427 ( 
.A(n_3952),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_3994),
.B(n_3356),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4080),
.B(n_3734),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_4229),
.B(n_3362),
.Y(n_4430)
);

CKINVDCx5p33_ASAP7_75t_R g4431 ( 
.A(n_3961),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_SL g4432 ( 
.A(n_4162),
.B(n_3782),
.Y(n_4432)
);

INVx3_ASAP7_75t_L g4433 ( 
.A(n_4282),
.Y(n_4433)
);

NAND2x1p5_ASAP7_75t_L g4434 ( 
.A(n_3968),
.B(n_3518),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_3865),
.B(n_3368),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4042),
.Y(n_4436)
);

AOI221x1_ASAP7_75t_L g4437 ( 
.A1(n_4017),
.A2(n_3833),
.B1(n_3829),
.B2(n_3806),
.C(n_3585),
.Y(n_4437)
);

NOR2xp33_ASAP7_75t_L g4438 ( 
.A(n_4028),
.B(n_4052),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4101),
.B(n_3370),
.Y(n_4439)
);

BUFx3_ASAP7_75t_L g4440 ( 
.A(n_4287),
.Y(n_4440)
);

AND2x4_ASAP7_75t_L g4441 ( 
.A(n_4078),
.B(n_3554),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4045),
.Y(n_4442)
);

BUFx8_ASAP7_75t_L g4443 ( 
.A(n_4125),
.Y(n_4443)
);

A2O1A1Ixp33_ASAP7_75t_L g4444 ( 
.A1(n_4166),
.A2(n_3756),
.B(n_3295),
.C(n_3507),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4055),
.Y(n_4445)
);

AOI22xp33_ASAP7_75t_L g4446 ( 
.A1(n_4021),
.A2(n_3840),
.B1(n_3536),
.B2(n_3742),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_SL g4447 ( 
.A(n_3851),
.B(n_3748),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_3925),
.B(n_3372),
.Y(n_4448)
);

AOI221xp5_ASAP7_75t_L g4449 ( 
.A1(n_3937),
.A2(n_3586),
.B1(n_3632),
.B2(n_3606),
.C(n_3599),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4139),
.B(n_3382),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4097),
.Y(n_4451)
);

OAI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_3863),
.A2(n_3911),
.B1(n_3864),
.B2(n_3905),
.Y(n_4452)
);

CKINVDCx5p33_ASAP7_75t_R g4453 ( 
.A(n_4026),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4140),
.B(n_4058),
.Y(n_4454)
);

AOI22xp5_ASAP7_75t_L g4455 ( 
.A1(n_4095),
.A2(n_3523),
.B1(n_3503),
.B2(n_3451),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_3989),
.B(n_3521),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4146),
.B(n_3522),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4072),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4170),
.B(n_3596),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4081),
.Y(n_4460)
);

CKINVDCx5p33_ASAP7_75t_R g4461 ( 
.A(n_3944),
.Y(n_4461)
);

NOR2xp33_ASAP7_75t_L g4462 ( 
.A(n_3980),
.B(n_3389),
.Y(n_4462)
);

CKINVDCx5p33_ASAP7_75t_R g4463 ( 
.A(n_4102),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_SL g4464 ( 
.A(n_4077),
.B(n_3639),
.Y(n_4464)
);

AND2x6_ASAP7_75t_L g4465 ( 
.A(n_4116),
.B(n_3856),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4090),
.B(n_3390),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4122),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4123),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_4173),
.B(n_3735),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4178),
.B(n_3393),
.Y(n_4470)
);

BUFx3_ASAP7_75t_L g4471 ( 
.A(n_4189),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4204),
.B(n_3421),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4219),
.Y(n_4473)
);

INVx3_ASAP7_75t_L g4474 ( 
.A(n_3996),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_4013),
.B(n_3428),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4098),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_3930),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_3949),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_3962),
.B(n_3457),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_3906),
.B(n_3459),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4151),
.Y(n_4481)
);

INVxp67_ASAP7_75t_L g4482 ( 
.A(n_4069),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4152),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_3955),
.B(n_3508),
.Y(n_4484)
);

BUFx6f_ASAP7_75t_L g4485 ( 
.A(n_3914),
.Y(n_4485)
);

INVx3_ASAP7_75t_L g4486 ( 
.A(n_3979),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4118),
.Y(n_4487)
);

BUFx3_ASAP7_75t_L g4488 ( 
.A(n_4000),
.Y(n_4488)
);

INVx3_ASAP7_75t_L g4489 ( 
.A(n_4074),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4079),
.B(n_3532),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_3929),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_SL g4492 ( 
.A(n_3971),
.B(n_3648),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4153),
.B(n_3509),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_4154),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4156),
.B(n_3548),
.Y(n_4495)
);

A2O1A1Ixp33_ASAP7_75t_L g4496 ( 
.A1(n_4033),
.A2(n_3665),
.B(n_3675),
.C(n_3664),
.Y(n_4496)
);

AOI22xp33_ASAP7_75t_L g4497 ( 
.A1(n_3879),
.A2(n_3705),
.B1(n_3708),
.B2(n_3678),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4082),
.B(n_3562),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4035),
.Y(n_4499)
);

OAI22xp5_ASAP7_75t_SL g4500 ( 
.A1(n_4100),
.A2(n_3723),
.B1(n_3729),
.B2(n_3709),
.Y(n_4500)
);

HB1xp67_ASAP7_75t_L g4501 ( 
.A(n_3902),
.Y(n_4501)
);

BUFx8_ASAP7_75t_L g4502 ( 
.A(n_4001),
.Y(n_4502)
);

AOI22xp33_ASAP7_75t_L g4503 ( 
.A1(n_4085),
.A2(n_3565),
.B1(n_3603),
.B2(n_3775),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4271),
.Y(n_4504)
);

CKINVDCx5p33_ASAP7_75t_R g4505 ( 
.A(n_3887),
.Y(n_4505)
);

CKINVDCx8_ASAP7_75t_R g4506 ( 
.A(n_3890),
.Y(n_4506)
);

BUFx3_ASAP7_75t_L g4507 ( 
.A(n_4002),
.Y(n_4507)
);

AND3x1_ASAP7_75t_SL g4508 ( 
.A(n_4200),
.B(n_345),
.C(n_346),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_3903),
.Y(n_4509)
);

BUFx6f_ASAP7_75t_L g4510 ( 
.A(n_4009),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_3977),
.Y(n_4511)
);

OAI22xp5_ASAP7_75t_SL g4512 ( 
.A1(n_4202),
.A2(n_3554),
.B1(n_348),
.B2(n_346),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_SL g4513 ( 
.A(n_3921),
.B(n_347),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4223),
.Y(n_4514)
);

BUFx3_ASAP7_75t_L g4515 ( 
.A(n_3982),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_R g4516 ( 
.A(n_4203),
.B(n_347),
.Y(n_4516)
);

INVx2_ASAP7_75t_L g4517 ( 
.A(n_3978),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4224),
.Y(n_4518)
);

BUFx2_ASAP7_75t_L g4519 ( 
.A(n_4197),
.Y(n_4519)
);

AOI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_4096),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_4004),
.Y(n_4521)
);

AOI22xp33_ASAP7_75t_L g4522 ( 
.A1(n_4186),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4225),
.Y(n_4523)
);

BUFx2_ASAP7_75t_L g4524 ( 
.A(n_4040),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4283),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4127),
.Y(n_4526)
);

BUFx6f_ASAP7_75t_L g4527 ( 
.A(n_3969),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_4285),
.Y(n_4528)
);

BUFx6f_ASAP7_75t_L g4529 ( 
.A(n_4070),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_SL g4530 ( 
.A(n_4205),
.B(n_351),
.Y(n_4530)
);

AND2x2_ASAP7_75t_L g4531 ( 
.A(n_4240),
.B(n_352),
.Y(n_4531)
);

AND2x4_ASAP7_75t_L g4532 ( 
.A(n_3858),
.B(n_352),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4244),
.B(n_353),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_3904),
.B(n_353),
.Y(n_4534)
);

AND3x1_ASAP7_75t_SL g4535 ( 
.A(n_4018),
.B(n_353),
.C(n_354),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4230),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4076),
.B(n_354),
.Y(n_4537)
);

AOI22xp33_ASAP7_75t_L g4538 ( 
.A1(n_4196),
.A2(n_4199),
.B1(n_4228),
.B2(n_4218),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_3934),
.Y(n_4539)
);

INVx2_ASAP7_75t_L g4540 ( 
.A(n_3935),
.Y(n_4540)
);

AND3x1_ASAP7_75t_SL g4541 ( 
.A(n_4141),
.B(n_355),
.C(n_356),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4231),
.B(n_355),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4083),
.B(n_356),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_3990),
.B(n_356),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_4031),
.B(n_357),
.Y(n_4545)
);

BUFx8_ASAP7_75t_L g4546 ( 
.A(n_3965),
.Y(n_4546)
);

BUFx12f_ASAP7_75t_L g4547 ( 
.A(n_3981),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_3991),
.B(n_357),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4220),
.Y(n_4549)
);

AOI22xp5_ASAP7_75t_L g4550 ( 
.A1(n_4063),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_4550)
);

INVx3_ASAP7_75t_L g4551 ( 
.A(n_3992),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_3993),
.B(n_358),
.Y(n_4552)
);

CKINVDCx5p33_ASAP7_75t_R g4553 ( 
.A(n_4142),
.Y(n_4553)
);

NAND2x1p5_ASAP7_75t_L g4554 ( 
.A(n_3995),
.B(n_358),
.Y(n_4554)
);

AND2x4_ASAP7_75t_L g4555 ( 
.A(n_4005),
.B(n_3997),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_3998),
.B(n_359),
.Y(n_4556)
);

INVx4_ASAP7_75t_L g4557 ( 
.A(n_4003),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_3939),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_3919),
.B(n_359),
.Y(n_4559)
);

CKINVDCx16_ASAP7_75t_R g4560 ( 
.A(n_4104),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4238),
.B(n_360),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_3964),
.B(n_3966),
.Y(n_4562)
);

A2O1A1Ixp33_ASAP7_75t_L g4563 ( 
.A1(n_4155),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_3868),
.B(n_361),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_4248),
.B(n_362),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4165),
.B(n_362),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_3945),
.Y(n_4567)
);

OR2x2_ASAP7_75t_L g4568 ( 
.A(n_4007),
.B(n_363),
.Y(n_4568)
);

INVx3_ASAP7_75t_L g4569 ( 
.A(n_4032),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_3947),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_3950),
.Y(n_4571)
);

OAI22xp5_ASAP7_75t_L g4572 ( 
.A1(n_3958),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_3953),
.Y(n_4573)
);

INVx3_ASAP7_75t_L g4574 ( 
.A(n_4034),
.Y(n_4574)
);

BUFx12f_ASAP7_75t_L g4575 ( 
.A(n_4128),
.Y(n_4575)
);

INVxp33_ASAP7_75t_L g4576 ( 
.A(n_3960),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4143),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4108),
.B(n_363),
.Y(n_4578)
);

OAI21x1_ASAP7_75t_L g4579 ( 
.A1(n_3940),
.A2(n_3943),
.B(n_3877),
.Y(n_4579)
);

INVx3_ASAP7_75t_L g4580 ( 
.A(n_3891),
.Y(n_4580)
);

AND3x1_ASAP7_75t_SL g4581 ( 
.A(n_4129),
.B(n_364),
.C(n_365),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4289),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4172),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_SL g4584 ( 
.A(n_3917),
.B(n_364),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4174),
.Y(n_4585)
);

AOI22xp33_ASAP7_75t_L g4586 ( 
.A1(n_4019),
.A2(n_4103),
.B1(n_4236),
.B2(n_4233),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4176),
.Y(n_4587)
);

AND2x4_ASAP7_75t_L g4588 ( 
.A(n_3923),
.B(n_365),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4099),
.B(n_366),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_4159),
.B(n_366),
.Y(n_4590)
);

BUFx8_ASAP7_75t_L g4591 ( 
.A(n_4131),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4291),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4111),
.B(n_367),
.Y(n_4593)
);

AND2x4_ASAP7_75t_L g4594 ( 
.A(n_3924),
.B(n_367),
.Y(n_4594)
);

BUFx6f_ASAP7_75t_L g4595 ( 
.A(n_3931),
.Y(n_4595)
);

INVxp67_ASAP7_75t_L g4596 ( 
.A(n_4158),
.Y(n_4596)
);

HB1xp67_ASAP7_75t_L g4597 ( 
.A(n_3873),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4161),
.B(n_368),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4181),
.Y(n_4599)
);

AND2x4_ASAP7_75t_L g4600 ( 
.A(n_3876),
.B(n_368),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4182),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4185),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4163),
.B(n_369),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_L g4604 ( 
.A(n_4164),
.B(n_369),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4227),
.B(n_370),
.Y(n_4605)
);

AND2x2_ASAP7_75t_L g4606 ( 
.A(n_4255),
.B(n_370),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4187),
.Y(n_4607)
);

BUFx2_ASAP7_75t_L g4608 ( 
.A(n_4239),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4256),
.B(n_371),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_3892),
.B(n_372),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4188),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4190),
.Y(n_4612)
);

AOI22xp33_ASAP7_75t_L g4613 ( 
.A1(n_4237),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_4613)
);

NOR2xp33_ASAP7_75t_L g4614 ( 
.A(n_4106),
.B(n_372),
.Y(n_4614)
);

NOR2xp67_ASAP7_75t_L g4615 ( 
.A(n_3888),
.B(n_4051),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4193),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4194),
.B(n_373),
.Y(n_4617)
);

INVx3_ASAP7_75t_L g4618 ( 
.A(n_3913),
.Y(n_4618)
);

CKINVDCx5p33_ASAP7_75t_R g4619 ( 
.A(n_4107),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4206),
.B(n_373),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4208),
.Y(n_4621)
);

INVx2_ASAP7_75t_L g4622 ( 
.A(n_4292),
.Y(n_4622)
);

INVx2_ASAP7_75t_SL g4623 ( 
.A(n_4054),
.Y(n_4623)
);

NOR2xp33_ASAP7_75t_L g4624 ( 
.A(n_3974),
.B(n_4241),
.Y(n_4624)
);

INVxp67_ASAP7_75t_L g4625 ( 
.A(n_4119),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4209),
.B(n_374),
.Y(n_4626)
);

AND2x2_ASAP7_75t_L g4627 ( 
.A(n_4261),
.B(n_375),
.Y(n_4627)
);

AND2x4_ASAP7_75t_L g4628 ( 
.A(n_3870),
.B(n_375),
.Y(n_4628)
);

NOR2xp67_ASAP7_75t_L g4629 ( 
.A(n_4136),
.B(n_375),
.Y(n_4629)
);

HB1xp67_ASAP7_75t_L g4630 ( 
.A(n_3912),
.Y(n_4630)
);

CKINVDCx5p33_ASAP7_75t_R g4631 ( 
.A(n_4138),
.Y(n_4631)
);

OAI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_3896),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4210),
.B(n_376),
.Y(n_4633)
);

AO21x2_ASAP7_75t_L g4634 ( 
.A1(n_4299),
.A2(n_3895),
.B(n_4109),
.Y(n_4634)
);

OAI21x1_ASAP7_75t_L g4635 ( 
.A1(n_4579),
.A2(n_4117),
.B(n_3963),
.Y(n_4635)
);

BUFx6f_ASAP7_75t_SL g4636 ( 
.A(n_4427),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4320),
.Y(n_4637)
);

OAI21x1_ASAP7_75t_L g4638 ( 
.A1(n_4336),
.A2(n_4088),
.B(n_4086),
.Y(n_4638)
);

AO21x2_ASAP7_75t_L g4639 ( 
.A1(n_4516),
.A2(n_4253),
.B(n_4075),
.Y(n_4639)
);

BUFx2_ASAP7_75t_L g4640 ( 
.A(n_4381),
.Y(n_4640)
);

INVx3_ASAP7_75t_L g4641 ( 
.A(n_4319),
.Y(n_4641)
);

OA21x2_ASAP7_75t_L g4642 ( 
.A1(n_4437),
.A2(n_4039),
.B(n_4037),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4305),
.B(n_4246),
.Y(n_4643)
);

INVx2_ASAP7_75t_L g4644 ( 
.A(n_4398),
.Y(n_4644)
);

INVx2_ASAP7_75t_SL g4645 ( 
.A(n_4319),
.Y(n_4645)
);

AOI22x1_ASAP7_75t_L g4646 ( 
.A1(n_4316),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4321),
.Y(n_4647)
);

INVx2_ASAP7_75t_SL g4648 ( 
.A(n_4298),
.Y(n_4648)
);

OAI21x1_ASAP7_75t_L g4649 ( 
.A1(n_4477),
.A2(n_4093),
.B(n_4091),
.Y(n_4649)
);

NOR2x1_ASAP7_75t_SL g4650 ( 
.A(n_4307),
.B(n_4311),
.Y(n_4650)
);

INVx1_ASAP7_75t_SL g4651 ( 
.A(n_4303),
.Y(n_4651)
);

OAI21x1_ASAP7_75t_L g4652 ( 
.A1(n_4492),
.A2(n_4094),
.B(n_3928),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4308),
.B(n_4280),
.Y(n_4653)
);

INVx3_ASAP7_75t_L g4654 ( 
.A(n_4431),
.Y(n_4654)
);

OAI21xp5_ASAP7_75t_L g4655 ( 
.A1(n_4437),
.A2(n_4050),
.B(n_4084),
.Y(n_4655)
);

INVx3_ASAP7_75t_L g4656 ( 
.A(n_4506),
.Y(n_4656)
);

INVx1_ASAP7_75t_SL g4657 ( 
.A(n_4306),
.Y(n_4657)
);

OA21x2_ASAP7_75t_L g4658 ( 
.A1(n_4345),
.A2(n_4043),
.B(n_4041),
.Y(n_4658)
);

INVx2_ASAP7_75t_SL g4659 ( 
.A(n_4345),
.Y(n_4659)
);

AOI21xp5_ASAP7_75t_L g4660 ( 
.A1(n_4404),
.A2(n_3918),
.B(n_4126),
.Y(n_4660)
);

OR2x6_ASAP7_75t_L g4661 ( 
.A(n_4328),
.B(n_4056),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_4312),
.Y(n_4662)
);

INVx2_ASAP7_75t_SL g4663 ( 
.A(n_4385),
.Y(n_4663)
);

AOI22x1_ASAP7_75t_L g4664 ( 
.A1(n_4316),
.A2(n_4560),
.B1(n_4368),
.B2(n_4394),
.Y(n_4664)
);

OAI21xp5_ASAP7_75t_L g4665 ( 
.A1(n_4497),
.A2(n_4148),
.B(n_4145),
.Y(n_4665)
);

INVx4_ASAP7_75t_L g4666 ( 
.A(n_4547),
.Y(n_4666)
);

HB1xp67_ASAP7_75t_SL g4667 ( 
.A(n_4443),
.Y(n_4667)
);

AO21x2_ASAP7_75t_L g4668 ( 
.A1(n_4408),
.A2(n_4046),
.B(n_4044),
.Y(n_4668)
);

OAI21xp5_ASAP7_75t_L g4669 ( 
.A1(n_4407),
.A2(n_4150),
.B(n_4110),
.Y(n_4669)
);

NAND2x1p5_ASAP7_75t_L g4670 ( 
.A(n_4474),
.B(n_4057),
.Y(n_4670)
);

BUFx5_ASAP7_75t_L g4671 ( 
.A(n_4302),
.Y(n_4671)
);

CKINVDCx5p33_ASAP7_75t_R g4672 ( 
.A(n_4318),
.Y(n_4672)
);

AND2x4_ASAP7_75t_L g4673 ( 
.A(n_4352),
.B(n_4059),
.Y(n_4673)
);

OAI21x1_ASAP7_75t_SL g4674 ( 
.A1(n_4310),
.A2(n_4175),
.B(n_4169),
.Y(n_4674)
);

OAI21x1_ASAP7_75t_L g4675 ( 
.A1(n_4421),
.A2(n_3926),
.B(n_4047),
.Y(n_4675)
);

OAI21x1_ASAP7_75t_L g4676 ( 
.A1(n_4504),
.A2(n_4049),
.B(n_4048),
.Y(n_4676)
);

AND2x4_ASAP7_75t_L g4677 ( 
.A(n_4302),
.B(n_4062),
.Y(n_4677)
);

BUFx6f_ASAP7_75t_L g4678 ( 
.A(n_4341),
.Y(n_4678)
);

OAI21x1_ASAP7_75t_L g4679 ( 
.A1(n_4487),
.A2(n_3909),
.B(n_4064),
.Y(n_4679)
);

INVx2_ASAP7_75t_SL g4680 ( 
.A(n_4385),
.Y(n_4680)
);

INVx2_ASAP7_75t_SL g4681 ( 
.A(n_4378),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4322),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4314),
.B(n_378),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4409),
.B(n_4262),
.Y(n_4684)
);

INVxp67_ASAP7_75t_SL g4685 ( 
.A(n_4386),
.Y(n_4685)
);

AND2x6_ASAP7_75t_L g4686 ( 
.A(n_4389),
.B(n_4133),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4390),
.Y(n_4687)
);

AO21x2_ASAP7_75t_L g4688 ( 
.A1(n_4513),
.A2(n_3894),
.B(n_3893),
.Y(n_4688)
);

AOI22x1_ASAP7_75t_L g4689 ( 
.A1(n_4461),
.A2(n_4393),
.B1(n_4505),
.B2(n_4463),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4400),
.B(n_4263),
.Y(n_4690)
);

NAND2x1p5_ASAP7_75t_L g4691 ( 
.A(n_4331),
.B(n_4066),
.Y(n_4691)
);

BUFx6f_ASAP7_75t_L g4692 ( 
.A(n_4341),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4342),
.B(n_4382),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4334),
.Y(n_4694)
);

CKINVDCx11_ASAP7_75t_R g4695 ( 
.A(n_4575),
.Y(n_4695)
);

BUFx12f_ASAP7_75t_L g4696 ( 
.A(n_4443),
.Y(n_4696)
);

BUFx2_ASAP7_75t_L g4697 ( 
.A(n_4515),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4315),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4339),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4353),
.Y(n_4700)
);

BUFx3_ASAP7_75t_L g4701 ( 
.A(n_4332),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4344),
.B(n_379),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4358),
.Y(n_4703)
);

AO21x2_ASAP7_75t_L g4704 ( 
.A1(n_4367),
.A2(n_4068),
.B(n_4067),
.Y(n_4704)
);

OAI21x1_ASAP7_75t_L g4705 ( 
.A1(n_4478),
.A2(n_4073),
.B(n_4071),
.Y(n_4705)
);

INVx3_ASAP7_75t_L g4706 ( 
.A(n_4502),
.Y(n_4706)
);

CKINVDCx5p33_ASAP7_75t_R g4707 ( 
.A(n_4313),
.Y(n_4707)
);

BUFx8_ASAP7_75t_L g4708 ( 
.A(n_4343),
.Y(n_4708)
);

BUFx6f_ASAP7_75t_L g4709 ( 
.A(n_4364),
.Y(n_4709)
);

AND2x4_ASAP7_75t_L g4710 ( 
.A(n_4359),
.B(n_3916),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4491),
.Y(n_4711)
);

OAI21x1_ASAP7_75t_L g4712 ( 
.A1(n_4489),
.A2(n_3885),
.B(n_3884),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4511),
.Y(n_4713)
);

AO21x2_ASAP7_75t_L g4714 ( 
.A1(n_4584),
.A2(n_4212),
.B(n_4211),
.Y(n_4714)
);

CKINVDCx5p33_ASAP7_75t_R g4715 ( 
.A(n_4313),
.Y(n_4715)
);

CKINVDCx20_ASAP7_75t_R g4716 ( 
.A(n_4411),
.Y(n_4716)
);

INVx1_ASAP7_75t_SL g4717 ( 
.A(n_4323),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4340),
.B(n_3897),
.Y(n_4718)
);

OAI21x1_ASAP7_75t_L g4719 ( 
.A1(n_4539),
.A2(n_4024),
.B(n_4022),
.Y(n_4719)
);

OAI21x1_ASAP7_75t_L g4720 ( 
.A1(n_4540),
.A2(n_3932),
.B(n_4268),
.Y(n_4720)
);

OR2x6_ASAP7_75t_L g4721 ( 
.A(n_4347),
.B(n_4232),
.Y(n_4721)
);

OAI21x1_ASAP7_75t_SL g4722 ( 
.A1(n_4338),
.A2(n_4168),
.B(n_4147),
.Y(n_4722)
);

OAI21x1_ASAP7_75t_L g4723 ( 
.A1(n_4558),
.A2(n_3933),
.B(n_4273),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4517),
.Y(n_4724)
);

CKINVDCx5p33_ASAP7_75t_R g4725 ( 
.A(n_4350),
.Y(n_4725)
);

BUFx6f_ASAP7_75t_L g4726 ( 
.A(n_4364),
.Y(n_4726)
);

AO21x2_ASAP7_75t_L g4727 ( 
.A1(n_4615),
.A2(n_4214),
.B(n_4213),
.Y(n_4727)
);

BUFx3_ASAP7_75t_L g4728 ( 
.A(n_4502),
.Y(n_4728)
);

BUFx4f_ASAP7_75t_SL g4729 ( 
.A(n_4546),
.Y(n_4729)
);

BUFx3_ASAP7_75t_L g4730 ( 
.A(n_4326),
.Y(n_4730)
);

HB1xp67_ASAP7_75t_L g4731 ( 
.A(n_4501),
.Y(n_4731)
);

AND2x4_ASAP7_75t_L g4732 ( 
.A(n_4374),
.B(n_3900),
.Y(n_4732)
);

OAI21x1_ASAP7_75t_L g4733 ( 
.A1(n_4567),
.A2(n_4279),
.B(n_4278),
.Y(n_4733)
);

BUFx2_ASAP7_75t_R g4734 ( 
.A(n_4366),
.Y(n_4734)
);

INVx1_ASAP7_75t_SL g4735 ( 
.A(n_4351),
.Y(n_4735)
);

OAI21x1_ASAP7_75t_L g4736 ( 
.A1(n_4570),
.A2(n_4276),
.B(n_4275),
.Y(n_4736)
);

AOI22x1_ASAP7_75t_L g4737 ( 
.A1(n_4608),
.A2(n_4453),
.B1(n_4524),
.B2(n_4519),
.Y(n_4737)
);

OAI21x1_ASAP7_75t_L g4738 ( 
.A1(n_4571),
.A2(n_4295),
.B(n_4294),
.Y(n_4738)
);

OR2x2_ASAP7_75t_L g4739 ( 
.A(n_4401),
.B(n_3901),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4376),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4402),
.B(n_379),
.Y(n_4741)
);

BUFx3_ASAP7_75t_L g4742 ( 
.A(n_4546),
.Y(n_4742)
);

NAND2x1p5_ASAP7_75t_L g4743 ( 
.A(n_4361),
.B(n_4120),
.Y(n_4743)
);

BUFx3_ASAP7_75t_L g4744 ( 
.A(n_4591),
.Y(n_4744)
);

OA21x2_ASAP7_75t_L g4745 ( 
.A1(n_4524),
.A2(n_4216),
.B(n_4215),
.Y(n_4745)
);

AND2x4_ASAP7_75t_L g4746 ( 
.A(n_4413),
.B(n_4557),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4456),
.Y(n_4747)
);

OAI21x1_ASAP7_75t_SL g4748 ( 
.A1(n_4452),
.A2(n_4258),
.B(n_4250),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_4333),
.B(n_379),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4392),
.B(n_4286),
.Y(n_4750)
);

OAI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_4370),
.A2(n_4121),
.B(n_4251),
.Y(n_4751)
);

BUFx3_ASAP7_75t_L g4752 ( 
.A(n_4591),
.Y(n_4752)
);

AO21x2_ASAP7_75t_L g4753 ( 
.A1(n_4629),
.A2(n_3886),
.B(n_4296),
.Y(n_4753)
);

INVx6_ASAP7_75t_L g4754 ( 
.A(n_4527),
.Y(n_4754)
);

INVx2_ASAP7_75t_L g4755 ( 
.A(n_4377),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4415),
.Y(n_4756)
);

OAI21x1_ASAP7_75t_L g4757 ( 
.A1(n_4573),
.A2(n_4113),
.B(n_4112),
.Y(n_4757)
);

AND2x4_ASAP7_75t_L g4758 ( 
.A(n_4405),
.B(n_4252),
.Y(n_4758)
);

AO21x2_ASAP7_75t_L g4759 ( 
.A1(n_4304),
.A2(n_4134),
.B(n_4171),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4509),
.Y(n_4760)
);

NAND2x1p5_ASAP7_75t_L g4761 ( 
.A(n_4608),
.B(n_4530),
.Y(n_4761)
);

OAI21x1_ASAP7_75t_L g4762 ( 
.A1(n_4486),
.A2(n_4115),
.B(n_4011),
.Y(n_4762)
);

BUFx12f_ASAP7_75t_L g4763 ( 
.A(n_4619),
.Y(n_4763)
);

OR2x2_ASAP7_75t_L g4764 ( 
.A(n_4396),
.B(n_380),
.Y(n_4764)
);

BUFx6f_ASAP7_75t_L g4765 ( 
.A(n_4527),
.Y(n_4765)
);

INVx3_ASAP7_75t_L g4766 ( 
.A(n_4488),
.Y(n_4766)
);

AO21x2_ASAP7_75t_L g4767 ( 
.A1(n_4564),
.A2(n_4281),
.B(n_4270),
.Y(n_4767)
);

BUFx8_ASAP7_75t_L g4768 ( 
.A(n_4600),
.Y(n_4768)
);

OAI21x1_ASAP7_75t_L g4769 ( 
.A1(n_4362),
.A2(n_4254),
.B(n_4012),
.Y(n_4769)
);

OAI21x1_ASAP7_75t_L g4770 ( 
.A1(n_4577),
.A2(n_4135),
.B(n_4016),
.Y(n_4770)
);

OAI21xp5_ASAP7_75t_L g4771 ( 
.A1(n_4444),
.A2(n_4027),
.B(n_4284),
.Y(n_4771)
);

OAI21x1_ASAP7_75t_L g4772 ( 
.A1(n_4451),
.A2(n_4015),
.B(n_4242),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4300),
.Y(n_4773)
);

NAND2x1p5_ASAP7_75t_L g4774 ( 
.A(n_4588),
.B(n_4243),
.Y(n_4774)
);

OR2x6_ASAP7_75t_L g4775 ( 
.A(n_4519),
.B(n_4264),
.Y(n_4775)
);

AO21x2_ASAP7_75t_L g4776 ( 
.A1(n_4475),
.A2(n_4267),
.B(n_4266),
.Y(n_4776)
);

CKINVDCx8_ASAP7_75t_R g4777 ( 
.A(n_4465),
.Y(n_4777)
);

INVx3_ASAP7_75t_L g4778 ( 
.A(n_4507),
.Y(n_4778)
);

BUFx3_ASAP7_75t_L g4779 ( 
.A(n_4434),
.Y(n_4779)
);

OR2x6_ASAP7_75t_L g4780 ( 
.A(n_4600),
.B(n_4269),
.Y(n_4780)
);

INVx6_ASAP7_75t_L g4781 ( 
.A(n_4510),
.Y(n_4781)
);

INVx1_ASAP7_75t_SL g4782 ( 
.A(n_4440),
.Y(n_4782)
);

INVx3_ASAP7_75t_L g4783 ( 
.A(n_4441),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4521),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4630),
.Y(n_4785)
);

AOI22x1_ASAP7_75t_L g4786 ( 
.A1(n_4423),
.A2(n_4553),
.B1(n_4631),
.B2(n_4425),
.Y(n_4786)
);

CKINVDCx16_ASAP7_75t_R g4787 ( 
.A(n_4384),
.Y(n_4787)
);

AOI22xp33_ASAP7_75t_L g4788 ( 
.A1(n_4512),
.A2(n_4235),
.B1(n_382),
.B2(n_380),
.Y(n_4788)
);

BUFx2_ASAP7_75t_SL g4789 ( 
.A(n_4383),
.Y(n_4789)
);

AO21x2_ASAP7_75t_L g4790 ( 
.A1(n_4388),
.A2(n_380),
.B(n_381),
.Y(n_4790)
);

INVx8_ASAP7_75t_L g4791 ( 
.A(n_4465),
.Y(n_4791)
);

INVx3_ASAP7_75t_L g4792 ( 
.A(n_4441),
.Y(n_4792)
);

CKINVDCx11_ASAP7_75t_R g4793 ( 
.A(n_4510),
.Y(n_4793)
);

BUFx3_ASAP7_75t_L g4794 ( 
.A(n_4471),
.Y(n_4794)
);

OAI21x1_ASAP7_75t_L g4795 ( 
.A1(n_4495),
.A2(n_594),
.B(n_593),
.Y(n_4795)
);

BUFx3_ASAP7_75t_L g4796 ( 
.A(n_4420),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4399),
.Y(n_4797)
);

AO21x2_ASAP7_75t_L g4798 ( 
.A1(n_4439),
.A2(n_381),
.B(n_382),
.Y(n_4798)
);

INVx2_ASAP7_75t_SL g4799 ( 
.A(n_4395),
.Y(n_4799)
);

BUFx10_ASAP7_75t_L g4800 ( 
.A(n_4324),
.Y(n_4800)
);

INVx3_ASAP7_75t_L g4801 ( 
.A(n_4418),
.Y(n_4801)
);

AO21x2_ASAP7_75t_L g4802 ( 
.A1(n_4432),
.A2(n_381),
.B(n_382),
.Y(n_4802)
);

BUFx6f_ASAP7_75t_L g4803 ( 
.A(n_4395),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4297),
.Y(n_4804)
);

BUFx12f_ASAP7_75t_L g4805 ( 
.A(n_4588),
.Y(n_4805)
);

INVx2_ASAP7_75t_L g4806 ( 
.A(n_4412),
.Y(n_4806)
);

INVx2_ASAP7_75t_SL g4807 ( 
.A(n_4529),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4325),
.Y(n_4808)
);

OAI21x1_ASAP7_75t_L g4809 ( 
.A1(n_4582),
.A2(n_595),
.B(n_593),
.Y(n_4809)
);

INVx3_ASAP7_75t_L g4810 ( 
.A(n_4551),
.Y(n_4810)
);

AND2x4_ASAP7_75t_L g4811 ( 
.A(n_4429),
.B(n_383),
.Y(n_4811)
);

OAI21x1_ASAP7_75t_L g4812 ( 
.A1(n_4592),
.A2(n_596),
.B(n_595),
.Y(n_4812)
);

NAND2x1p5_ASAP7_75t_L g4813 ( 
.A(n_4594),
.B(n_383),
.Y(n_4813)
);

AO21x2_ASAP7_75t_L g4814 ( 
.A1(n_4481),
.A2(n_384),
.B(n_385),
.Y(n_4814)
);

CKINVDCx20_ASAP7_75t_R g4815 ( 
.A(n_4355),
.Y(n_4815)
);

OA21x2_ASAP7_75t_L g4816 ( 
.A1(n_4483),
.A2(n_385),
.B(n_386),
.Y(n_4816)
);

AOI22x1_ASAP7_75t_L g4817 ( 
.A1(n_4554),
.A2(n_388),
.B1(n_385),
.B2(n_387),
.Y(n_4817)
);

BUFx4_ASAP7_75t_SL g4818 ( 
.A(n_4476),
.Y(n_4818)
);

INVx4_ASAP7_75t_L g4819 ( 
.A(n_4465),
.Y(n_4819)
);

AOI22x1_ASAP7_75t_L g4820 ( 
.A1(n_4532),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_4820)
);

AOI22x1_ASAP7_75t_L g4821 ( 
.A1(n_4532),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4329),
.Y(n_4822)
);

BUFx2_ASAP7_75t_R g4823 ( 
.A(n_4369),
.Y(n_4823)
);

NAND2x1p5_ASAP7_75t_L g4824 ( 
.A(n_4594),
.B(n_390),
.Y(n_4824)
);

BUFx2_ASAP7_75t_L g4825 ( 
.A(n_4391),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4458),
.Y(n_4826)
);

AND2x4_ASAP7_75t_L g4827 ( 
.A(n_4555),
.B(n_390),
.Y(n_4827)
);

NAND2x1p5_ASAP7_75t_L g4828 ( 
.A(n_4628),
.B(n_390),
.Y(n_4828)
);

OAI21x1_ASAP7_75t_L g4829 ( 
.A1(n_4622),
.A2(n_597),
.B(n_596),
.Y(n_4829)
);

INVx3_ASAP7_75t_SL g4830 ( 
.A(n_4555),
.Y(n_4830)
);

OAI21x1_ASAP7_75t_L g4831 ( 
.A1(n_4494),
.A2(n_599),
.B(n_598),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_L g4832 ( 
.A(n_4330),
.B(n_391),
.Y(n_4832)
);

OAI21xp5_ASAP7_75t_L g4833 ( 
.A1(n_4563),
.A2(n_391),
.B(n_392),
.Y(n_4833)
);

BUFx24_ASAP7_75t_L g4834 ( 
.A(n_4628),
.Y(n_4834)
);

BUFx12f_ASAP7_75t_L g4835 ( 
.A(n_4485),
.Y(n_4835)
);

OR2x6_ASAP7_75t_L g4836 ( 
.A(n_4482),
.B(n_391),
.Y(n_4836)
);

BUFx2_ASAP7_75t_SL g4837 ( 
.A(n_4562),
.Y(n_4837)
);

BUFx2_ASAP7_75t_L g4838 ( 
.A(n_4485),
.Y(n_4838)
);

AND2x2_ASAP7_75t_L g4839 ( 
.A(n_4335),
.B(n_392),
.Y(n_4839)
);

OAI21x1_ASAP7_75t_L g4840 ( 
.A1(n_4499),
.A2(n_599),
.B(n_598),
.Y(n_4840)
);

BUFx12f_ASAP7_75t_L g4841 ( 
.A(n_4623),
.Y(n_4841)
);

INVx2_ASAP7_75t_L g4842 ( 
.A(n_4416),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4468),
.Y(n_4843)
);

OAI21x1_ASAP7_75t_L g4844 ( 
.A1(n_4514),
.A2(n_601),
.B(n_600),
.Y(n_4844)
);

BUFx6f_ASAP7_75t_L g4845 ( 
.A(n_4529),
.Y(n_4845)
);

NAND2x1p5_ASAP7_75t_L g4846 ( 
.A(n_4544),
.B(n_4552),
.Y(n_4846)
);

INVx3_ASAP7_75t_L g4847 ( 
.A(n_4529),
.Y(n_4847)
);

OAI21x1_ASAP7_75t_L g4848 ( 
.A1(n_4518),
.A2(n_601),
.B(n_600),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4473),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4337),
.Y(n_4850)
);

AND2x4_ASAP7_75t_L g4851 ( 
.A(n_4580),
.B(n_392),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4597),
.Y(n_4852)
);

OAI21x1_ASAP7_75t_L g4853 ( 
.A1(n_4523),
.A2(n_603),
.B(n_602),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4406),
.Y(n_4854)
);

INVx1_ASAP7_75t_SL g4855 ( 
.A(n_4410),
.Y(n_4855)
);

INVx6_ASAP7_75t_SL g4856 ( 
.A(n_4327),
.Y(n_4856)
);

AO21x2_ASAP7_75t_L g4857 ( 
.A1(n_4357),
.A2(n_393),
.B(n_394),
.Y(n_4857)
);

BUFx2_ASAP7_75t_L g4858 ( 
.A(n_4730),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4854),
.Y(n_4859)
);

AOI22xp33_ASAP7_75t_SL g4860 ( 
.A1(n_4737),
.A2(n_4791),
.B1(n_4837),
.B2(n_4805),
.Y(n_4860)
);

AOI22xp33_ASAP7_75t_L g4861 ( 
.A1(n_4791),
.A2(n_4301),
.B1(n_4500),
.B2(n_4576),
.Y(n_4861)
);

BUFx2_ASAP7_75t_L g4862 ( 
.A(n_4716),
.Y(n_4862)
);

AOI22xp33_ASAP7_75t_L g4863 ( 
.A1(n_4780),
.A2(n_4538),
.B1(n_4356),
.B2(n_4586),
.Y(n_4863)
);

BUFx4f_ASAP7_75t_SL g4864 ( 
.A(n_4696),
.Y(n_4864)
);

AOI22xp33_ASAP7_75t_SL g4865 ( 
.A1(n_4768),
.A2(n_4569),
.B1(n_4574),
.B2(n_4618),
.Y(n_4865)
);

AOI22xp5_ASAP7_75t_L g4866 ( 
.A1(n_4815),
.A2(n_4721),
.B1(n_4780),
.B2(n_4424),
.Y(n_4866)
);

AOI22xp33_ASAP7_75t_L g4867 ( 
.A1(n_4722),
.A2(n_4348),
.B1(n_4464),
.B2(n_4438),
.Y(n_4867)
);

OAI22xp5_ASAP7_75t_L g4868 ( 
.A1(n_4777),
.A2(n_4596),
.B1(n_4503),
.B2(n_4625),
.Y(n_4868)
);

AOI22xp33_ASAP7_75t_SL g4869 ( 
.A1(n_4786),
.A2(n_4556),
.B1(n_4433),
.B2(n_4595),
.Y(n_4869)
);

CKINVDCx6p67_ASAP7_75t_R g4870 ( 
.A(n_4744),
.Y(n_4870)
);

CKINVDCx11_ASAP7_75t_R g4871 ( 
.A(n_4695),
.Y(n_4871)
);

NAND2x1p5_ASAP7_75t_L g4872 ( 
.A(n_4742),
.B(n_4752),
.Y(n_4872)
);

BUFx3_ASAP7_75t_L g4873 ( 
.A(n_4794),
.Y(n_4873)
);

OAI22xp5_ASAP7_75t_L g4874 ( 
.A1(n_4777),
.A2(n_4446),
.B1(n_4371),
.B2(n_4455),
.Y(n_4874)
);

AOI22xp33_ASAP7_75t_L g4875 ( 
.A1(n_4646),
.A2(n_4526),
.B1(n_4583),
.B2(n_4536),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4647),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4682),
.Y(n_4877)
);

AOI22xp33_ASAP7_75t_L g4878 ( 
.A1(n_4775),
.A2(n_4585),
.B1(n_4599),
.B2(n_4587),
.Y(n_4878)
);

INVx3_ASAP7_75t_L g4879 ( 
.A(n_4729),
.Y(n_4879)
);

OAI22xp5_ASAP7_75t_L g4880 ( 
.A1(n_4775),
.A2(n_4520),
.B1(n_4496),
.B2(n_4550),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4806),
.Y(n_4881)
);

AOI22xp5_ASAP7_75t_L g4882 ( 
.A1(n_4721),
.A2(n_4414),
.B1(n_4535),
.B2(n_4581),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4842),
.Y(n_4883)
);

OAI21xp5_ASAP7_75t_SL g4884 ( 
.A1(n_4706),
.A2(n_4614),
.B(n_4522),
.Y(n_4884)
);

BUFx8_ASAP7_75t_L g4885 ( 
.A(n_4636),
.Y(n_4885)
);

CKINVDCx11_ASAP7_75t_R g4886 ( 
.A(n_4793),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4826),
.Y(n_4887)
);

AOI22xp33_ASAP7_75t_L g4888 ( 
.A1(n_4674),
.A2(n_4601),
.B1(n_4607),
.B2(n_4602),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4843),
.Y(n_4889)
);

AOI22xp33_ASAP7_75t_L g4890 ( 
.A1(n_4820),
.A2(n_4611),
.B1(n_4616),
.B2(n_4612),
.Y(n_4890)
);

BUFx2_ASAP7_75t_L g4891 ( 
.A(n_4701),
.Y(n_4891)
);

NAND2x1p5_ASAP7_75t_L g4892 ( 
.A(n_4728),
.B(n_4578),
.Y(n_4892)
);

OAI22xp33_ASAP7_75t_L g4893 ( 
.A1(n_4787),
.A2(n_4568),
.B1(n_4621),
.B2(n_4559),
.Y(n_4893)
);

INVx2_ASAP7_75t_L g4894 ( 
.A(n_4713),
.Y(n_4894)
);

AOI22xp33_ASAP7_75t_L g4895 ( 
.A1(n_4821),
.A2(n_4449),
.B1(n_4605),
.B2(n_4624),
.Y(n_4895)
);

INVx2_ASAP7_75t_SL g4896 ( 
.A(n_4708),
.Y(n_4896)
);

CKINVDCx5p33_ASAP7_75t_R g4897 ( 
.A(n_4667),
.Y(n_4897)
);

AOI22xp33_ASAP7_75t_L g4898 ( 
.A1(n_4748),
.A2(n_4533),
.B1(n_4542),
.B2(n_4531),
.Y(n_4898)
);

AND2x2_ASAP7_75t_L g4899 ( 
.A(n_4657),
.B(n_4735),
.Y(n_4899)
);

INVx1_ASAP7_75t_SL g4900 ( 
.A(n_4782),
.Y(n_4900)
);

NAND2x1p5_ASAP7_75t_L g4901 ( 
.A(n_4666),
.B(n_4593),
.Y(n_4901)
);

CKINVDCx11_ASAP7_75t_R g4902 ( 
.A(n_4651),
.Y(n_4902)
);

AOI22xp33_ASAP7_75t_L g4903 ( 
.A1(n_4759),
.A2(n_4525),
.B1(n_4528),
.B2(n_4606),
.Y(n_4903)
);

CKINVDCx11_ASAP7_75t_R g4904 ( 
.A(n_4800),
.Y(n_4904)
);

BUFx6f_ASAP7_75t_L g4905 ( 
.A(n_4678),
.Y(n_4905)
);

BUFx12f_ASAP7_75t_L g4906 ( 
.A(n_4707),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4808),
.B(n_4417),
.Y(n_4907)
);

CKINVDCx20_ASAP7_75t_R g4908 ( 
.A(n_4672),
.Y(n_4908)
);

BUFx8_ASAP7_75t_L g4909 ( 
.A(n_4763),
.Y(n_4909)
);

AOI22xp33_ASAP7_75t_L g4910 ( 
.A1(n_4661),
.A2(n_4595),
.B1(n_4462),
.B2(n_4627),
.Y(n_4910)
);

AOI22xp33_ASAP7_75t_L g4911 ( 
.A1(n_4661),
.A2(n_4549),
.B1(n_4543),
.B2(n_4565),
.Y(n_4911)
);

INVx2_ASAP7_75t_L g4912 ( 
.A(n_4724),
.Y(n_4912)
);

CKINVDCx11_ASAP7_75t_R g4913 ( 
.A(n_4640),
.Y(n_4913)
);

AOI22xp33_ASAP7_75t_L g4914 ( 
.A1(n_4639),
.A2(n_4387),
.B1(n_4572),
.B2(n_4537),
.Y(n_4914)
);

AOI22xp33_ASAP7_75t_L g4915 ( 
.A1(n_4686),
.A2(n_4435),
.B1(n_4534),
.B2(n_4436),
.Y(n_4915)
);

CKINVDCx5p33_ASAP7_75t_R g4916 ( 
.A(n_4715),
.Y(n_4916)
);

HB1xp67_ASAP7_75t_L g4917 ( 
.A(n_4717),
.Y(n_4917)
);

INVx2_ASAP7_75t_L g4918 ( 
.A(n_4711),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4849),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_SL g4920 ( 
.A1(n_4819),
.A2(n_4309),
.B(n_4447),
.Y(n_4920)
);

BUFx2_ASAP7_75t_L g4921 ( 
.A(n_4697),
.Y(n_4921)
);

AOI22xp33_ASAP7_75t_L g4922 ( 
.A1(n_4686),
.A2(n_4422),
.B1(n_4445),
.B2(n_4442),
.Y(n_4922)
);

BUFx6f_ASAP7_75t_L g4923 ( 
.A(n_4678),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4804),
.B(n_4460),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4797),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4773),
.Y(n_4926)
);

INVx6_ASAP7_75t_L g4927 ( 
.A(n_4835),
.Y(n_4927)
);

BUFx10_ASAP7_75t_L g4928 ( 
.A(n_4836),
.Y(n_4928)
);

INVx1_ASAP7_75t_SL g4929 ( 
.A(n_4818),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4687),
.Y(n_4930)
);

BUFx3_ASAP7_75t_L g4931 ( 
.A(n_4662),
.Y(n_4931)
);

BUFx6f_ASAP7_75t_L g4932 ( 
.A(n_4692),
.Y(n_4932)
);

OAI21xp5_ASAP7_75t_SL g4933 ( 
.A1(n_4656),
.A2(n_4613),
.B(n_4632),
.Y(n_4933)
);

BUFx4_ASAP7_75t_SL g4934 ( 
.A(n_4725),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4694),
.Y(n_4935)
);

AOI22xp33_ASAP7_75t_L g4936 ( 
.A1(n_4686),
.A2(n_4467),
.B1(n_4454),
.B2(n_4561),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4699),
.Y(n_4937)
);

BUFx8_ASAP7_75t_L g4938 ( 
.A(n_4841),
.Y(n_4938)
);

BUFx2_ASAP7_75t_L g4939 ( 
.A(n_4766),
.Y(n_4939)
);

HB1xp67_ASAP7_75t_L g4940 ( 
.A(n_4731),
.Y(n_4940)
);

BUFx6f_ASAP7_75t_L g4941 ( 
.A(n_4692),
.Y(n_4941)
);

AND2x4_ASAP7_75t_SL g4942 ( 
.A(n_4641),
.B(n_4457),
.Y(n_4942)
);

BUFx2_ASAP7_75t_L g4943 ( 
.A(n_4778),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4700),
.Y(n_4944)
);

BUFx2_ASAP7_75t_L g4945 ( 
.A(n_4856),
.Y(n_4945)
);

AOI22xp5_ASAP7_75t_L g4946 ( 
.A1(n_4855),
.A2(n_4541),
.B1(n_4508),
.B2(n_4430),
.Y(n_4946)
);

AOI22xp5_ASAP7_75t_L g4947 ( 
.A1(n_4836),
.A2(n_4448),
.B1(n_4450),
.B2(n_4480),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4703),
.Y(n_4948)
);

BUFx10_ASAP7_75t_L g4949 ( 
.A(n_4851),
.Y(n_4949)
);

INVx2_ASAP7_75t_L g4950 ( 
.A(n_4637),
.Y(n_4950)
);

AOI22xp33_ASAP7_75t_L g4951 ( 
.A1(n_4796),
.A2(n_4589),
.B1(n_4490),
.B2(n_4566),
.Y(n_4951)
);

AND2x2_ASAP7_75t_L g4952 ( 
.A(n_4740),
.B(n_4346),
.Y(n_4952)
);

INVx2_ASAP7_75t_L g4953 ( 
.A(n_4644),
.Y(n_4953)
);

CKINVDCx5p33_ASAP7_75t_R g4954 ( 
.A(n_4734),
.Y(n_4954)
);

AOI22xp33_ASAP7_75t_L g4955 ( 
.A1(n_4827),
.A2(n_4372),
.B1(n_4609),
.B2(n_4363),
.Y(n_4955)
);

BUFx8_ASAP7_75t_SL g4956 ( 
.A(n_4654),
.Y(n_4956)
);

INVx3_ASAP7_75t_L g4957 ( 
.A(n_4779),
.Y(n_4957)
);

CKINVDCx11_ASAP7_75t_R g4958 ( 
.A(n_4830),
.Y(n_4958)
);

AOI22xp33_ASAP7_75t_SL g4959 ( 
.A1(n_4789),
.A2(n_4469),
.B1(n_4459),
.B2(n_4354),
.Y(n_4959)
);

BUFx2_ASAP7_75t_L g4960 ( 
.A(n_4645),
.Y(n_4960)
);

AOI22xp33_ASAP7_75t_SL g4961 ( 
.A1(n_4664),
.A2(n_4365),
.B1(n_4373),
.B2(n_4375),
.Y(n_4961)
);

BUFx6f_ASAP7_75t_L g4962 ( 
.A(n_4709),
.Y(n_4962)
);

INVx6_ASAP7_75t_L g4963 ( 
.A(n_4709),
.Y(n_4963)
);

AOI22xp33_ASAP7_75t_SL g4964 ( 
.A1(n_4671),
.A2(n_4379),
.B1(n_4380),
.B2(n_4317),
.Y(n_4964)
);

AOI22xp33_ASAP7_75t_SL g4965 ( 
.A1(n_4671),
.A2(n_4650),
.B1(n_4761),
.B2(n_4828),
.Y(n_4965)
);

INVx5_ASAP7_75t_L g4966 ( 
.A(n_4765),
.Y(n_4966)
);

HB1xp67_ASAP7_75t_L g4967 ( 
.A(n_4755),
.Y(n_4967)
);

BUFx2_ASAP7_75t_L g4968 ( 
.A(n_4645),
.Y(n_4968)
);

CKINVDCx16_ASAP7_75t_R g4969 ( 
.A(n_4702),
.Y(n_4969)
);

CKINVDCx11_ASAP7_75t_R g4970 ( 
.A(n_4726),
.Y(n_4970)
);

OAI22xp5_ASAP7_75t_L g4971 ( 
.A1(n_4813),
.A2(n_4479),
.B1(n_4403),
.B2(n_4426),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4698),
.Y(n_4972)
);

AOI22xp33_ASAP7_75t_L g4973 ( 
.A1(n_4817),
.A2(n_4811),
.B1(n_4758),
.B2(n_4788),
.Y(n_4973)
);

INVx4_ASAP7_75t_L g4974 ( 
.A(n_4726),
.Y(n_4974)
);

BUFx2_ASAP7_75t_SL g4975 ( 
.A(n_4671),
.Y(n_4975)
);

INVx4_ASAP7_75t_L g4976 ( 
.A(n_4781),
.Y(n_4976)
);

AOI22xp5_ASAP7_75t_L g4977 ( 
.A1(n_4677),
.A2(n_4349),
.B1(n_4472),
.B2(n_4470),
.Y(n_4977)
);

AOI22xp5_ASAP7_75t_L g4978 ( 
.A1(n_4669),
.A2(n_4493),
.B1(n_4466),
.B2(n_4484),
.Y(n_4978)
);

INVx8_ASAP7_75t_L g4979 ( 
.A(n_4834),
.Y(n_4979)
);

AOI22xp33_ASAP7_75t_L g4980 ( 
.A1(n_4767),
.A2(n_4545),
.B1(n_4598),
.B2(n_4590),
.Y(n_4980)
);

CKINVDCx11_ASAP7_75t_R g4981 ( 
.A(n_4825),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4760),
.Y(n_4982)
);

BUFx4_ASAP7_75t_R g4983 ( 
.A(n_4823),
.Y(n_4983)
);

AOI22xp33_ASAP7_75t_SL g4984 ( 
.A1(n_4824),
.A2(n_4548),
.B1(n_4360),
.B2(n_4428),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_4852),
.Y(n_4985)
);

AOI22xp33_ASAP7_75t_L g4986 ( 
.A1(n_4776),
.A2(n_4774),
.B1(n_4771),
.B2(n_4710),
.Y(n_4986)
);

INVx6_ASAP7_75t_L g4987 ( 
.A(n_4803),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4784),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4747),
.Y(n_4989)
);

BUFx3_ASAP7_75t_L g4990 ( 
.A(n_4838),
.Y(n_4990)
);

BUFx2_ASAP7_75t_SL g4991 ( 
.A(n_4648),
.Y(n_4991)
);

AOI22xp33_ASAP7_75t_L g4992 ( 
.A1(n_4746),
.A2(n_4604),
.B1(n_4603),
.B2(n_4617),
.Y(n_4992)
);

BUFx2_ASAP7_75t_SL g4993 ( 
.A(n_4648),
.Y(n_4993)
);

BUFx2_ASAP7_75t_SL g4994 ( 
.A(n_4681),
.Y(n_4994)
);

CKINVDCx5p33_ASAP7_75t_R g4995 ( 
.A(n_4689),
.Y(n_4995)
);

INVx2_ASAP7_75t_SL g4996 ( 
.A(n_4754),
.Y(n_4996)
);

CKINVDCx5p33_ASAP7_75t_R g4997 ( 
.A(n_4702),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4935),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4937),
.Y(n_4999)
);

AND2x2_ASAP7_75t_L g5000 ( 
.A(n_4858),
.B(n_4822),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4967),
.B(n_4989),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4944),
.Y(n_5002)
);

CKINVDCx11_ASAP7_75t_R g5003 ( 
.A(n_4871),
.Y(n_5003)
);

AOI22xp33_ASAP7_75t_L g5004 ( 
.A1(n_4863),
.A2(n_4655),
.B1(n_4846),
.B2(n_4634),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_L g5005 ( 
.A(n_4917),
.B(n_4785),
.Y(n_5005)
);

OAI21x1_ASAP7_75t_L g5006 ( 
.A1(n_4878),
.A2(n_4712),
.B(n_4635),
.Y(n_5006)
);

BUFx6f_ASAP7_75t_L g5007 ( 
.A(n_4958),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4948),
.Y(n_5008)
);

AOI21xp5_ASAP7_75t_L g5009 ( 
.A1(n_4920),
.A2(n_4660),
.B(n_4659),
.Y(n_5009)
);

OAI31xp33_ASAP7_75t_L g5010 ( 
.A1(n_4874),
.A2(n_4691),
.A3(n_4743),
.B(n_4670),
.Y(n_5010)
);

OA21x2_ASAP7_75t_L g5011 ( 
.A1(n_4986),
.A2(n_4762),
.B(n_4652),
.Y(n_5011)
);

INVx2_ASAP7_75t_L g5012 ( 
.A(n_4899),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4891),
.Y(n_5013)
);

OA21x2_ASAP7_75t_L g5014 ( 
.A1(n_4888),
.A2(n_4693),
.B(n_4720),
.Y(n_5014)
);

AO21x1_ASAP7_75t_L g5015 ( 
.A1(n_4942),
.A2(n_4685),
.B(n_4741),
.Y(n_5015)
);

OA21x2_ASAP7_75t_L g5016 ( 
.A1(n_4866),
.A2(n_4675),
.B(n_4659),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4982),
.Y(n_5017)
);

AO31x2_ASAP7_75t_L g5018 ( 
.A1(n_4939),
.A2(n_4756),
.A3(n_4850),
.B(n_4643),
.Y(n_5018)
);

AOI21xp5_ASAP7_75t_L g5019 ( 
.A1(n_4965),
.A2(n_4745),
.B(n_4658),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_4930),
.B(n_4653),
.Y(n_5020)
);

OAI21x1_ASAP7_75t_L g5021 ( 
.A1(n_4903),
.A2(n_4922),
.B(n_4936),
.Y(n_5021)
);

OR2x2_ASAP7_75t_L g5022 ( 
.A(n_4940),
.B(n_4739),
.Y(n_5022)
);

A2O1A1Ixp33_ASAP7_75t_L g5023 ( 
.A1(n_4979),
.A2(n_4751),
.B(n_4665),
.C(n_4833),
.Y(n_5023)
);

AOI21x1_ASAP7_75t_L g5024 ( 
.A1(n_4896),
.A2(n_4816),
.B(n_4642),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4926),
.B(n_4653),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_4988),
.B(n_4810),
.Y(n_5026)
);

AOI22xp33_ASAP7_75t_L g5027 ( 
.A1(n_4880),
.A2(n_4790),
.B1(n_4704),
.B2(n_4673),
.Y(n_5027)
);

HB1xp67_ASAP7_75t_L g5028 ( 
.A(n_4921),
.Y(n_5028)
);

AOI22xp33_ASAP7_75t_L g5029 ( 
.A1(n_4861),
.A2(n_4668),
.B1(n_4727),
.B2(n_4732),
.Y(n_5029)
);

OA21x2_ASAP7_75t_L g5030 ( 
.A1(n_4943),
.A2(n_4723),
.B(n_4679),
.Y(n_5030)
);

OR2x6_ASAP7_75t_L g5031 ( 
.A(n_4979),
.B(n_4681),
.Y(n_5031)
);

HB1xp67_ASAP7_75t_L g5032 ( 
.A(n_4900),
.Y(n_5032)
);

INVx2_ASAP7_75t_L g5033 ( 
.A(n_4894),
.Y(n_5033)
);

HB1xp67_ASAP7_75t_L g5034 ( 
.A(n_4873),
.Y(n_5034)
);

NAND3xp33_ASAP7_75t_L g5035 ( 
.A(n_4867),
.B(n_4832),
.C(n_4764),
.Y(n_5035)
);

AOI221xp5_ASAP7_75t_L g5036 ( 
.A1(n_4893),
.A2(n_4690),
.B1(n_4750),
.B2(n_4684),
.C(n_4610),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_4985),
.B(n_4718),
.Y(n_5037)
);

NOR2xp33_ASAP7_75t_L g5038 ( 
.A(n_4902),
.B(n_4801),
.Y(n_5038)
);

OA21x2_ASAP7_75t_L g5039 ( 
.A1(n_4980),
.A2(n_4638),
.B(n_4772),
.Y(n_5039)
);

AOI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4860),
.A2(n_4753),
.B(n_4688),
.Y(n_5040)
);

HB1xp67_ASAP7_75t_L g5041 ( 
.A(n_4969),
.Y(n_5041)
);

AOI21xp5_ASAP7_75t_L g5042 ( 
.A1(n_4869),
.A2(n_4807),
.B(n_4680),
.Y(n_5042)
);

HB1xp67_ASAP7_75t_L g5043 ( 
.A(n_4960),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4859),
.Y(n_5044)
);

CKINVDCx16_ASAP7_75t_R g5045 ( 
.A(n_4929),
.Y(n_5045)
);

OAI21x1_ASAP7_75t_L g5046 ( 
.A1(n_4971),
.A2(n_4847),
.B(n_4705),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4881),
.B(n_4683),
.Y(n_5047)
);

OAI21xp5_ASAP7_75t_L g5048 ( 
.A1(n_4882),
.A2(n_4676),
.B(n_4831),
.Y(n_5048)
);

OR2x2_ASAP7_75t_L g5049 ( 
.A(n_4883),
.B(n_4807),
.Y(n_5049)
);

OR2x2_ASAP7_75t_L g5050 ( 
.A(n_4887),
.B(n_4683),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4968),
.B(n_4783),
.Y(n_5051)
);

INVx2_ASAP7_75t_L g5052 ( 
.A(n_4912),
.Y(n_5052)
);

HB1xp67_ASAP7_75t_L g5053 ( 
.A(n_4950),
.Y(n_5053)
);

AOI221xp5_ASAP7_75t_L g5054 ( 
.A1(n_4914),
.A2(n_4397),
.B1(n_4620),
.B2(n_4633),
.C(n_4626),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4889),
.B(n_4749),
.Y(n_5055)
);

AO31x2_ASAP7_75t_L g5056 ( 
.A1(n_4868),
.A2(n_4419),
.A3(n_4498),
.B(n_4754),
.Y(n_5056)
);

AND2x4_ASAP7_75t_L g5057 ( 
.A(n_4990),
.B(n_4792),
.Y(n_5057)
);

BUFx6f_ASAP7_75t_L g5058 ( 
.A(n_4905),
.Y(n_5058)
);

OAI22xp33_ASAP7_75t_L g5059 ( 
.A1(n_4997),
.A2(n_4946),
.B1(n_4995),
.B2(n_4947),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4876),
.Y(n_5060)
);

OA21x2_ASAP7_75t_L g5061 ( 
.A1(n_4915),
.A2(n_4757),
.B(n_4649),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_4919),
.B(n_4749),
.Y(n_5062)
);

OAI21x1_ASAP7_75t_L g5063 ( 
.A1(n_4872),
.A2(n_4769),
.B(n_4738),
.Y(n_5063)
);

CKINVDCx11_ASAP7_75t_R g5064 ( 
.A(n_4908),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_SL g5065 ( 
.A(n_4959),
.B(n_4765),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_L g5066 ( 
.A(n_4907),
.B(n_4839),
.Y(n_5066)
);

OAI21x1_ASAP7_75t_L g5067 ( 
.A1(n_4957),
.A2(n_4736),
.B(n_4733),
.Y(n_5067)
);

AO21x2_ASAP7_75t_L g5068 ( 
.A1(n_4924),
.A2(n_4798),
.B(n_4857),
.Y(n_5068)
);

OR2x6_ASAP7_75t_L g5069 ( 
.A(n_4994),
.B(n_4663),
.Y(n_5069)
);

AOI21xp5_ASAP7_75t_L g5070 ( 
.A1(n_4890),
.A2(n_4875),
.B(n_4961),
.Y(n_5070)
);

OAI21x1_ASAP7_75t_L g5071 ( 
.A1(n_4901),
.A2(n_4719),
.B(n_4770),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4877),
.Y(n_5072)
);

AND2x2_ASAP7_75t_L g5073 ( 
.A(n_4952),
.B(n_4663),
.Y(n_5073)
);

OA21x2_ASAP7_75t_L g5074 ( 
.A1(n_4911),
.A2(n_4925),
.B(n_4910),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4953),
.Y(n_5075)
);

AO21x2_ASAP7_75t_L g5076 ( 
.A1(n_4978),
.A2(n_4814),
.B(n_4795),
.Y(n_5076)
);

OAI21x1_ASAP7_75t_L g5077 ( 
.A1(n_4892),
.A2(n_4844),
.B(n_4840),
.Y(n_5077)
);

A2O1A1Ixp33_ASAP7_75t_L g5078 ( 
.A1(n_4884),
.A2(n_4839),
.B(n_4853),
.C(n_4848),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4972),
.Y(n_5079)
);

CKINVDCx5p33_ASAP7_75t_R g5080 ( 
.A(n_4897),
.Y(n_5080)
);

INVx2_ASAP7_75t_L g5081 ( 
.A(n_4918),
.Y(n_5081)
);

OR2x2_ASAP7_75t_L g5082 ( 
.A(n_4991),
.B(n_4993),
.Y(n_5082)
);

AOI22xp5_ASAP7_75t_L g5083 ( 
.A1(n_4898),
.A2(n_4802),
.B1(n_4714),
.B2(n_4680),
.Y(n_5083)
);

INVx2_ASAP7_75t_L g5084 ( 
.A(n_4981),
.Y(n_5084)
);

BUFx3_ASAP7_75t_L g5085 ( 
.A(n_4870),
.Y(n_5085)
);

INVx2_ASAP7_75t_L g5086 ( 
.A(n_4987),
.Y(n_5086)
);

AOI22xp5_ASAP7_75t_SL g5087 ( 
.A1(n_4954),
.A2(n_4799),
.B1(n_4845),
.B2(n_4803),
.Y(n_5087)
);

HB1xp67_ASAP7_75t_L g5088 ( 
.A(n_4996),
.Y(n_5088)
);

AND2x4_ASAP7_75t_L g5089 ( 
.A(n_4974),
.B(n_4799),
.Y(n_5089)
);

OR2x6_ASAP7_75t_L g5090 ( 
.A(n_4927),
.B(n_4862),
.Y(n_5090)
);

OAI21x1_ASAP7_75t_L g5091 ( 
.A1(n_4879),
.A2(n_4812),
.B(n_4809),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_4928),
.B(n_4945),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4977),
.Y(n_5093)
);

OR2x2_ASAP7_75t_L g5094 ( 
.A(n_4976),
.B(n_4845),
.Y(n_5094)
);

A2O1A1Ixp33_ASAP7_75t_L g5095 ( 
.A1(n_4865),
.A2(n_4933),
.B(n_4973),
.C(n_4984),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4964),
.A2(n_4829),
.B(n_393),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_L g5097 ( 
.A(n_4951),
.B(n_393),
.Y(n_5097)
);

AOI21x1_ASAP7_75t_L g5098 ( 
.A1(n_4983),
.A2(n_394),
.B(n_395),
.Y(n_5098)
);

AOI222xp33_ASAP7_75t_L g5099 ( 
.A1(n_4895),
.A2(n_396),
.B1(n_398),
.B2(n_394),
.C1(n_395),
.C2(n_397),
.Y(n_5099)
);

OA21x2_ASAP7_75t_L g5100 ( 
.A1(n_4992),
.A2(n_395),
.B(n_396),
.Y(n_5100)
);

AOI21xp5_ASAP7_75t_L g5101 ( 
.A1(n_4955),
.A2(n_396),
.B(n_397),
.Y(n_5101)
);

OR2x2_ASAP7_75t_L g5102 ( 
.A(n_5022),
.B(n_4975),
.Y(n_5102)
);

AOI22xp33_ASAP7_75t_L g5103 ( 
.A1(n_5059),
.A2(n_4913),
.B1(n_4904),
.B2(n_4949),
.Y(n_5103)
);

AO31x2_ASAP7_75t_L g5104 ( 
.A1(n_5095),
.A2(n_5015),
.A3(n_5040),
.B(n_5019),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5001),
.Y(n_5105)
);

AND2x2_ASAP7_75t_L g5106 ( 
.A(n_5073),
.B(n_4931),
.Y(n_5106)
);

AOI22xp33_ASAP7_75t_L g5107 ( 
.A1(n_5004),
.A2(n_4927),
.B1(n_4885),
.B2(n_4987),
.Y(n_5107)
);

OR2x2_ASAP7_75t_L g5108 ( 
.A(n_5053),
.B(n_4905),
.Y(n_5108)
);

OAI22xp5_ASAP7_75t_L g5109 ( 
.A1(n_5031),
.A2(n_4864),
.B1(n_4963),
.B2(n_4966),
.Y(n_5109)
);

AO31x2_ASAP7_75t_L g5110 ( 
.A1(n_5013),
.A2(n_5023),
.A3(n_5070),
.B(n_5038),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_4998),
.Y(n_5111)
);

AOI221xp5_ASAP7_75t_L g5112 ( 
.A1(n_5093),
.A2(n_4916),
.B1(n_4932),
.B2(n_4941),
.C(n_4923),
.Y(n_5112)
);

AOI22xp33_ASAP7_75t_L g5113 ( 
.A1(n_5010),
.A2(n_4970),
.B1(n_4963),
.B2(n_4886),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5025),
.B(n_4923),
.Y(n_5114)
);

BUFx4f_ASAP7_75t_SL g5115 ( 
.A(n_5007),
.Y(n_5115)
);

OA21x2_ASAP7_75t_L g5116 ( 
.A1(n_5048),
.A2(n_5046),
.B(n_5021),
.Y(n_5116)
);

INVxp67_ASAP7_75t_L g5117 ( 
.A(n_5034),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_5012),
.B(n_4932),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4999),
.Y(n_5119)
);

AOI22xp33_ASAP7_75t_SL g5120 ( 
.A1(n_5041),
.A2(n_4938),
.B1(n_4909),
.B2(n_4966),
.Y(n_5120)
);

OAI221xp5_ASAP7_75t_L g5121 ( 
.A1(n_5029),
.A2(n_4941),
.B1(n_4962),
.B2(n_4966),
.C(n_4934),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_5020),
.B(n_4962),
.Y(n_5122)
);

AOI22xp5_ASAP7_75t_L g5123 ( 
.A1(n_5036),
.A2(n_4906),
.B1(n_4956),
.B2(n_399),
.Y(n_5123)
);

AOI22xp33_ASAP7_75t_L g5124 ( 
.A1(n_5074),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_5124)
);

OAI22xp5_ASAP7_75t_L g5125 ( 
.A1(n_5031),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_5125)
);

OR2x2_ASAP7_75t_L g5126 ( 
.A(n_5037),
.B(n_5028),
.Y(n_5126)
);

OAI21x1_ASAP7_75t_L g5127 ( 
.A1(n_5006),
.A2(n_400),
.B(n_401),
.Y(n_5127)
);

AOI22xp33_ASAP7_75t_L g5128 ( 
.A1(n_5027),
.A2(n_403),
.B1(n_400),
.B2(n_402),
.Y(n_5128)
);

OAI22xp33_ASAP7_75t_L g5129 ( 
.A1(n_5069),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_5129)
);

OAI221xp5_ASAP7_75t_SL g5130 ( 
.A1(n_5083),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.C(n_407),
.Y(n_5130)
);

CKINVDCx6p67_ASAP7_75t_R g5131 ( 
.A(n_5003),
.Y(n_5131)
);

OAI22xp5_ASAP7_75t_L g5132 ( 
.A1(n_5069),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_5132)
);

AOI221xp5_ASAP7_75t_SL g5133 ( 
.A1(n_5009),
.A2(n_5042),
.B1(n_5078),
.B2(n_5065),
.C(n_5000),
.Y(n_5133)
);

AOI221xp5_ASAP7_75t_L g5134 ( 
.A1(n_5035),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.C(n_410),
.Y(n_5134)
);

OAI21x1_ASAP7_75t_L g5135 ( 
.A1(n_5024),
.A2(n_407),
.B(n_408),
.Y(n_5135)
);

OR2x2_ASAP7_75t_L g5136 ( 
.A(n_5005),
.B(n_408),
.Y(n_5136)
);

OR2x2_ASAP7_75t_L g5137 ( 
.A(n_5066),
.B(n_409),
.Y(n_5137)
);

OAI221xp5_ASAP7_75t_L g5138 ( 
.A1(n_5098),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.C(n_412),
.Y(n_5138)
);

NOR2x1_ASAP7_75t_SL g5139 ( 
.A(n_5082),
.B(n_410),
.Y(n_5139)
);

AOI22xp33_ASAP7_75t_L g5140 ( 
.A1(n_5054),
.A2(n_414),
.B1(n_411),
.B2(n_412),
.Y(n_5140)
);

AOI22xp33_ASAP7_75t_L g5141 ( 
.A1(n_5100),
.A2(n_414),
.B1(n_411),
.B2(n_412),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_5002),
.Y(n_5142)
);

OAI22xp5_ASAP7_75t_L g5143 ( 
.A1(n_5090),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_5143)
);

BUFx4f_ASAP7_75t_SL g5144 ( 
.A(n_5007),
.Y(n_5144)
);

OAI211xp5_ASAP7_75t_L g5145 ( 
.A1(n_5099),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_5145)
);

INVx3_ASAP7_75t_L g5146 ( 
.A(n_5090),
.Y(n_5146)
);

AOI22xp33_ASAP7_75t_L g5147 ( 
.A1(n_5096),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_5075),
.B(n_418),
.Y(n_5148)
);

AOI22xp33_ASAP7_75t_SL g5149 ( 
.A1(n_5016),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_5149)
);

INVx2_ASAP7_75t_L g5150 ( 
.A(n_5018),
.Y(n_5150)
);

OAI211xp5_ASAP7_75t_SL g5151 ( 
.A1(n_5097),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5008),
.Y(n_5152)
);

OAI221xp5_ASAP7_75t_L g5153 ( 
.A1(n_5014),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_5153)
);

AOI21xp5_ASAP7_75t_L g5154 ( 
.A1(n_5087),
.A2(n_422),
.B(n_423),
.Y(n_5154)
);

BUFx4f_ASAP7_75t_SL g5155 ( 
.A(n_5085),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_5017),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_5044),
.Y(n_5157)
);

A2O1A1Ixp33_ASAP7_75t_L g5158 ( 
.A1(n_5092),
.A2(n_425),
.B(n_422),
.C(n_424),
.Y(n_5158)
);

INVx2_ASAP7_75t_L g5159 ( 
.A(n_5018),
.Y(n_5159)
);

AOI221xp5_ASAP7_75t_L g5160 ( 
.A1(n_5101),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.C(n_428),
.Y(n_5160)
);

NOR2xp33_ASAP7_75t_SL g5161 ( 
.A(n_5045),
.B(n_427),
.Y(n_5161)
);

A2O1A1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_5063),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_5162)
);

BUFx3_ASAP7_75t_L g5163 ( 
.A(n_5064),
.Y(n_5163)
);

INVx8_ASAP7_75t_L g5164 ( 
.A(n_5080),
.Y(n_5164)
);

A2O1A1Ixp33_ASAP7_75t_L g5165 ( 
.A1(n_5084),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_5165)
);

AND2x2_ASAP7_75t_L g5166 ( 
.A(n_5043),
.B(n_429),
.Y(n_5166)
);

AOI22xp33_ASAP7_75t_L g5167 ( 
.A1(n_5076),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_5167)
);

AOI22xp33_ASAP7_75t_L g5168 ( 
.A1(n_5032),
.A2(n_434),
.B1(n_431),
.B2(n_432),
.Y(n_5168)
);

AND2x2_ASAP7_75t_L g5169 ( 
.A(n_5051),
.B(n_431),
.Y(n_5169)
);

OAI22xp33_ASAP7_75t_L g5170 ( 
.A1(n_5088),
.A2(n_435),
.B1(n_432),
.B2(n_434),
.Y(n_5170)
);

AND2x2_ASAP7_75t_L g5171 ( 
.A(n_5057),
.B(n_435),
.Y(n_5171)
);

INVx4_ASAP7_75t_L g5172 ( 
.A(n_5058),
.Y(n_5172)
);

AOI22xp33_ASAP7_75t_L g5173 ( 
.A1(n_5068),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_5173)
);

INVx2_ASAP7_75t_SL g5174 ( 
.A(n_5089),
.Y(n_5174)
);

INVx2_ASAP7_75t_L g5175 ( 
.A(n_5033),
.Y(n_5175)
);

OAI21xp33_ASAP7_75t_L g5176 ( 
.A1(n_5026),
.A2(n_436),
.B(n_437),
.Y(n_5176)
);

AOI22xp33_ASAP7_75t_L g5177 ( 
.A1(n_5011),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_5177)
);

AOI22xp33_ASAP7_75t_L g5178 ( 
.A1(n_5061),
.A2(n_440),
.B1(n_438),
.B2(n_439),
.Y(n_5178)
);

AND2x2_ASAP7_75t_L g5179 ( 
.A(n_5086),
.B(n_439),
.Y(n_5179)
);

OR2x2_ASAP7_75t_L g5180 ( 
.A(n_5050),
.B(n_440),
.Y(n_5180)
);

CKINVDCx5p33_ASAP7_75t_R g5181 ( 
.A(n_5058),
.Y(n_5181)
);

OAI22xp33_ASAP7_75t_L g5182 ( 
.A1(n_5094),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5060),
.Y(n_5183)
);

OAI21xp5_ASAP7_75t_SL g5184 ( 
.A1(n_5047),
.A2(n_441),
.B(n_442),
.Y(n_5184)
);

AND2x4_ASAP7_75t_L g5185 ( 
.A(n_5067),
.B(n_441),
.Y(n_5185)
);

AOI22xp33_ASAP7_75t_L g5186 ( 
.A1(n_5077),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_5186)
);

INVx2_ASAP7_75t_L g5187 ( 
.A(n_5052),
.Y(n_5187)
);

AOI22xp33_ASAP7_75t_SL g5188 ( 
.A1(n_5039),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_5188)
);

OAI221xp5_ASAP7_75t_L g5189 ( 
.A1(n_5055),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.C(n_446),
.Y(n_5189)
);

HB1xp67_ASAP7_75t_L g5190 ( 
.A(n_5117),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_5111),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5119),
.Y(n_5192)
);

OR2x2_ASAP7_75t_L g5193 ( 
.A(n_5126),
.B(n_5062),
.Y(n_5193)
);

AND2x2_ASAP7_75t_L g5194 ( 
.A(n_5146),
.B(n_5056),
.Y(n_5194)
);

AND2x2_ASAP7_75t_L g5195 ( 
.A(n_5174),
.B(n_5056),
.Y(n_5195)
);

AOI22xp33_ASAP7_75t_L g5196 ( 
.A1(n_5123),
.A2(n_5039),
.B1(n_5072),
.B2(n_5030),
.Y(n_5196)
);

AND2x2_ASAP7_75t_L g5197 ( 
.A(n_5118),
.B(n_5079),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5142),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_5152),
.Y(n_5199)
);

OR2x2_ASAP7_75t_L g5200 ( 
.A(n_5105),
.B(n_5081),
.Y(n_5200)
);

AND2x2_ASAP7_75t_L g5201 ( 
.A(n_5106),
.B(n_5049),
.Y(n_5201)
);

AND2x4_ASAP7_75t_SL g5202 ( 
.A(n_5131),
.B(n_5071),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5156),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_5175),
.Y(n_5204)
);

INVx2_ASAP7_75t_L g5205 ( 
.A(n_5187),
.Y(n_5205)
);

INVx3_ASAP7_75t_L g5206 ( 
.A(n_5172),
.Y(n_5206)
);

NOR2xp67_ASAP7_75t_L g5207 ( 
.A(n_5109),
.B(n_5121),
.Y(n_5207)
);

AND2x2_ASAP7_75t_L g5208 ( 
.A(n_5108),
.B(n_5091),
.Y(n_5208)
);

OA21x2_ASAP7_75t_L g5209 ( 
.A1(n_5133),
.A2(n_445),
.B(n_446),
.Y(n_5209)
);

OR2x2_ASAP7_75t_L g5210 ( 
.A(n_5157),
.B(n_447),
.Y(n_5210)
);

AND2x2_ASAP7_75t_L g5211 ( 
.A(n_5102),
.B(n_447),
.Y(n_5211)
);

INVx2_ASAP7_75t_SL g5212 ( 
.A(n_5155),
.Y(n_5212)
);

BUFx4f_ASAP7_75t_SL g5213 ( 
.A(n_5163),
.Y(n_5213)
);

AND2x2_ASAP7_75t_L g5214 ( 
.A(n_5116),
.B(n_448),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5116),
.B(n_448),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_5183),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_5122),
.B(n_448),
.Y(n_5217)
);

AND2x2_ASAP7_75t_L g5218 ( 
.A(n_5114),
.B(n_449),
.Y(n_5218)
);

AND2x4_ASAP7_75t_L g5219 ( 
.A(n_5185),
.B(n_450),
.Y(n_5219)
);

OAI221xp5_ASAP7_75t_L g5220 ( 
.A1(n_5184),
.A2(n_5161),
.B1(n_5149),
.B2(n_5103),
.C(n_5107),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_5148),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_5166),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_5150),
.B(n_450),
.Y(n_5223)
);

INVx2_ASAP7_75t_L g5224 ( 
.A(n_5159),
.Y(n_5224)
);

INVx2_ASAP7_75t_L g5225 ( 
.A(n_5180),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5136),
.Y(n_5226)
);

AOI22xp33_ASAP7_75t_L g5227 ( 
.A1(n_5153),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_5227)
);

INVx2_ASAP7_75t_SL g5228 ( 
.A(n_5181),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_5137),
.Y(n_5229)
);

INVx2_ASAP7_75t_L g5230 ( 
.A(n_5127),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5104),
.B(n_451),
.Y(n_5231)
);

HB1xp67_ASAP7_75t_L g5232 ( 
.A(n_5104),
.Y(n_5232)
);

HB1xp67_ASAP7_75t_L g5233 ( 
.A(n_5110),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_5169),
.Y(n_5234)
);

INVx2_ASAP7_75t_SL g5235 ( 
.A(n_5164),
.Y(n_5235)
);

INVx4_ASAP7_75t_R g5236 ( 
.A(n_5120),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_5135),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_5179),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_5171),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_L g5240 ( 
.A(n_5178),
.B(n_451),
.Y(n_5240)
);

AND2x4_ASAP7_75t_L g5241 ( 
.A(n_5110),
.B(n_452),
.Y(n_5241)
);

AND2x2_ASAP7_75t_L g5242 ( 
.A(n_5113),
.B(n_452),
.Y(n_5242)
);

OAI211xp5_ASAP7_75t_L g5243 ( 
.A1(n_5154),
.A2(n_455),
.B(n_453),
.C(n_454),
.Y(n_5243)
);

INVx2_ASAP7_75t_SL g5244 ( 
.A(n_5164),
.Y(n_5244)
);

INVx2_ASAP7_75t_L g5245 ( 
.A(n_5139),
.Y(n_5245)
);

INVx3_ASAP7_75t_L g5246 ( 
.A(n_5115),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_5132),
.Y(n_5247)
);

AND2x2_ASAP7_75t_L g5248 ( 
.A(n_5112),
.B(n_454),
.Y(n_5248)
);

OR2x2_ASAP7_75t_L g5249 ( 
.A(n_5177),
.B(n_454),
.Y(n_5249)
);

AOI221xp5_ASAP7_75t_L g5250 ( 
.A1(n_5189),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.C(n_458),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_5143),
.Y(n_5251)
);

AOI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_5209),
.A2(n_5162),
.B(n_5124),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_5214),
.B(n_5188),
.Y(n_5253)
);

AND2x2_ASAP7_75t_L g5254 ( 
.A(n_5206),
.B(n_5167),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_5206),
.B(n_5128),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_5204),
.Y(n_5256)
);

BUFx6f_ASAP7_75t_L g5257 ( 
.A(n_5246),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5190),
.Y(n_5258)
);

INVx1_ASAP7_75t_SL g5259 ( 
.A(n_5213),
.Y(n_5259)
);

OAI22xp33_ASAP7_75t_L g5260 ( 
.A1(n_5209),
.A2(n_5138),
.B1(n_5125),
.B2(n_5144),
.Y(n_5260)
);

INVxp67_ASAP7_75t_SL g5261 ( 
.A(n_5231),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_5205),
.Y(n_5262)
);

INVx2_ASAP7_75t_L g5263 ( 
.A(n_5190),
.Y(n_5263)
);

AOI21xp5_ASAP7_75t_L g5264 ( 
.A1(n_5241),
.A2(n_5220),
.B(n_5231),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_SL g5265 ( 
.A(n_5241),
.B(n_5129),
.Y(n_5265)
);

HB1xp67_ASAP7_75t_L g5266 ( 
.A(n_5215),
.Y(n_5266)
);

INVxp67_ASAP7_75t_L g5267 ( 
.A(n_5242),
.Y(n_5267)
);

INVxp67_ASAP7_75t_L g5268 ( 
.A(n_5248),
.Y(n_5268)
);

AOI21x1_ASAP7_75t_L g5269 ( 
.A1(n_5232),
.A2(n_5145),
.B(n_5130),
.Y(n_5269)
);

OAI22xp5_ASAP7_75t_L g5270 ( 
.A1(n_5220),
.A2(n_5173),
.B1(n_5141),
.B2(n_5158),
.Y(n_5270)
);

INVx2_ASAP7_75t_L g5271 ( 
.A(n_5200),
.Y(n_5271)
);

A2O1A1Ixp33_ASAP7_75t_L g5272 ( 
.A1(n_5207),
.A2(n_5176),
.B(n_5134),
.C(n_5165),
.Y(n_5272)
);

AO21x2_ASAP7_75t_L g5273 ( 
.A1(n_5232),
.A2(n_5170),
.B(n_5182),
.Y(n_5273)
);

OR2x2_ASAP7_75t_L g5274 ( 
.A(n_5193),
.B(n_5186),
.Y(n_5274)
);

HB1xp67_ASAP7_75t_L g5275 ( 
.A(n_5191),
.Y(n_5275)
);

OA21x2_ASAP7_75t_L g5276 ( 
.A1(n_5233),
.A2(n_5147),
.B(n_5140),
.Y(n_5276)
);

A2O1A1Ixp33_ASAP7_75t_L g5277 ( 
.A1(n_5207),
.A2(n_5151),
.B(n_5160),
.C(n_5168),
.Y(n_5277)
);

INVx2_ASAP7_75t_L g5278 ( 
.A(n_5224),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5192),
.Y(n_5279)
);

INVx2_ASAP7_75t_L g5280 ( 
.A(n_5237),
.Y(n_5280)
);

INVx2_ASAP7_75t_L g5281 ( 
.A(n_5230),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5198),
.Y(n_5282)
);

INVx2_ASAP7_75t_L g5283 ( 
.A(n_5199),
.Y(n_5283)
);

AOI21x1_ASAP7_75t_L g5284 ( 
.A1(n_5233),
.A2(n_456),
.B(n_457),
.Y(n_5284)
);

OR2x2_ASAP7_75t_L g5285 ( 
.A(n_5221),
.B(n_457),
.Y(n_5285)
);

AND2x4_ASAP7_75t_L g5286 ( 
.A(n_5202),
.B(n_458),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_5203),
.Y(n_5287)
);

NAND4xp25_ASAP7_75t_L g5288 ( 
.A(n_5196),
.B(n_460),
.C(n_458),
.D(n_459),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5216),
.Y(n_5289)
);

INVx2_ASAP7_75t_L g5290 ( 
.A(n_5219),
.Y(n_5290)
);

INVx2_ASAP7_75t_L g5291 ( 
.A(n_5219),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5223),
.Y(n_5292)
);

INVx3_ASAP7_75t_L g5293 ( 
.A(n_5213),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5225),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5229),
.Y(n_5295)
);

OAI22xp33_ASAP7_75t_L g5296 ( 
.A1(n_5245),
.A2(n_462),
.B1(n_459),
.B2(n_461),
.Y(n_5296)
);

INVx2_ASAP7_75t_L g5297 ( 
.A(n_5197),
.Y(n_5297)
);

INVxp67_ASAP7_75t_SL g5298 ( 
.A(n_5211),
.Y(n_5298)
);

OAI21xp33_ASAP7_75t_SL g5299 ( 
.A1(n_5196),
.A2(n_459),
.B(n_461),
.Y(n_5299)
);

O2A1O1Ixp33_ASAP7_75t_L g5300 ( 
.A1(n_5247),
.A2(n_463),
.B(n_461),
.C(n_462),
.Y(n_5300)
);

BUFx6f_ASAP7_75t_SL g5301 ( 
.A(n_5212),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_5208),
.Y(n_5302)
);

OAI22xp33_ASAP7_75t_L g5303 ( 
.A1(n_5195),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_5303)
);

OAI21x1_ASAP7_75t_L g5304 ( 
.A1(n_5194),
.A2(n_463),
.B(n_464),
.Y(n_5304)
);

BUFx2_ASAP7_75t_L g5305 ( 
.A(n_5228),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_L g5306 ( 
.A1(n_5235),
.A2(n_465),
.B(n_466),
.Y(n_5306)
);

BUFx2_ASAP7_75t_L g5307 ( 
.A(n_5246),
.Y(n_5307)
);

INVxp67_ASAP7_75t_SL g5308 ( 
.A(n_5251),
.Y(n_5308)
);

AOI222xp33_ASAP7_75t_L g5309 ( 
.A1(n_5226),
.A2(n_467),
.B1(n_469),
.B2(n_465),
.C1(n_466),
.C2(n_468),
.Y(n_5309)
);

BUFx2_ASAP7_75t_L g5310 ( 
.A(n_5244),
.Y(n_5310)
);

INVx2_ASAP7_75t_L g5311 ( 
.A(n_5201),
.Y(n_5311)
);

OAI22xp5_ASAP7_75t_L g5312 ( 
.A1(n_5222),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_5312)
);

BUFx2_ASAP7_75t_L g5313 ( 
.A(n_5239),
.Y(n_5313)
);

OA21x2_ASAP7_75t_L g5314 ( 
.A1(n_5238),
.A2(n_467),
.B(n_468),
.Y(n_5314)
);

OA21x2_ASAP7_75t_L g5315 ( 
.A1(n_5234),
.A2(n_5218),
.B(n_5217),
.Y(n_5315)
);

OAI22xp5_ASAP7_75t_L g5316 ( 
.A1(n_5210),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_5316)
);

OR2x2_ASAP7_75t_L g5317 ( 
.A(n_5240),
.B(n_469),
.Y(n_5317)
);

NOR2xp33_ASAP7_75t_R g5318 ( 
.A(n_5236),
.B(n_5249),
.Y(n_5318)
);

OAI22xp5_ASAP7_75t_L g5319 ( 
.A1(n_5308),
.A2(n_5236),
.B1(n_5227),
.B2(n_5243),
.Y(n_5319)
);

INVx1_ASAP7_75t_SL g5320 ( 
.A(n_5259),
.Y(n_5320)
);

HB1xp67_ASAP7_75t_L g5321 ( 
.A(n_5263),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_5258),
.Y(n_5322)
);

AO21x2_ASAP7_75t_L g5323 ( 
.A1(n_5264),
.A2(n_5318),
.B(n_5273),
.Y(n_5323)
);

AND2x4_ASAP7_75t_L g5324 ( 
.A(n_5307),
.B(n_5240),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_5266),
.B(n_5227),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_5261),
.B(n_5250),
.Y(n_5326)
);

AND2x2_ASAP7_75t_L g5327 ( 
.A(n_5310),
.B(n_5250),
.Y(n_5327)
);

AND2x2_ASAP7_75t_L g5328 ( 
.A(n_5305),
.B(n_5243),
.Y(n_5328)
);

HB1xp67_ASAP7_75t_L g5329 ( 
.A(n_5314),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5275),
.Y(n_5330)
);

OR2x2_ASAP7_75t_L g5331 ( 
.A(n_5295),
.B(n_470),
.Y(n_5331)
);

AND2x2_ASAP7_75t_L g5332 ( 
.A(n_5286),
.B(n_470),
.Y(n_5332)
);

AND2x2_ASAP7_75t_L g5333 ( 
.A(n_5286),
.B(n_5254),
.Y(n_5333)
);

NAND3xp33_ASAP7_75t_L g5334 ( 
.A(n_5299),
.B(n_471),
.C(n_472),
.Y(n_5334)
);

OR2x2_ASAP7_75t_L g5335 ( 
.A(n_5274),
.B(n_472),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_5276),
.B(n_473),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_L g5337 ( 
.A(n_5276),
.B(n_473),
.Y(n_5337)
);

AND2x2_ASAP7_75t_L g5338 ( 
.A(n_5255),
.B(n_474),
.Y(n_5338)
);

AOI222xp33_ASAP7_75t_L g5339 ( 
.A1(n_5270),
.A2(n_476),
.B1(n_478),
.B2(n_474),
.C1(n_475),
.C2(n_477),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_L g5340 ( 
.A(n_5303),
.B(n_474),
.Y(n_5340)
);

AND2x2_ASAP7_75t_L g5341 ( 
.A(n_5257),
.B(n_475),
.Y(n_5341)
);

OAI22xp5_ASAP7_75t_L g5342 ( 
.A1(n_5315),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_5314),
.Y(n_5343)
);

AND2x2_ASAP7_75t_L g5344 ( 
.A(n_5257),
.B(n_5315),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_5268),
.B(n_476),
.Y(n_5345)
);

OR2x2_ASAP7_75t_L g5346 ( 
.A(n_5294),
.B(n_477),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5284),
.Y(n_5347)
);

BUFx3_ASAP7_75t_L g5348 ( 
.A(n_5293),
.Y(n_5348)
);

INVx3_ASAP7_75t_L g5349 ( 
.A(n_5257),
.Y(n_5349)
);

BUFx3_ASAP7_75t_L g5350 ( 
.A(n_5304),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5292),
.Y(n_5351)
);

OR2x2_ASAP7_75t_L g5352 ( 
.A(n_5271),
.B(n_478),
.Y(n_5352)
);

HB1xp67_ASAP7_75t_L g5353 ( 
.A(n_5281),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5279),
.Y(n_5354)
);

BUFx6f_ASAP7_75t_L g5355 ( 
.A(n_5317),
.Y(n_5355)
);

AND2x2_ASAP7_75t_L g5356 ( 
.A(n_5313),
.B(n_478),
.Y(n_5356)
);

OR2x2_ASAP7_75t_L g5357 ( 
.A(n_5282),
.B(n_479),
.Y(n_5357)
);

AND2x2_ASAP7_75t_L g5358 ( 
.A(n_5311),
.B(n_479),
.Y(n_5358)
);

AND2x2_ASAP7_75t_L g5359 ( 
.A(n_5298),
.B(n_479),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_5267),
.B(n_5253),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5287),
.Y(n_5361)
);

AND2x2_ASAP7_75t_L g5362 ( 
.A(n_5297),
.B(n_480),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5289),
.Y(n_5363)
);

INVx2_ASAP7_75t_L g5364 ( 
.A(n_5290),
.Y(n_5364)
);

OR2x2_ASAP7_75t_L g5365 ( 
.A(n_5283),
.B(n_481),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_5291),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_5280),
.Y(n_5367)
);

OAI22xp5_ASAP7_75t_L g5368 ( 
.A1(n_5302),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_5285),
.Y(n_5369)
);

AOI21xp33_ASAP7_75t_L g5370 ( 
.A1(n_5260),
.A2(n_483),
.B(n_484),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_5269),
.Y(n_5371)
);

INVx2_ASAP7_75t_L g5372 ( 
.A(n_5256),
.Y(n_5372)
);

AND2x2_ASAP7_75t_L g5373 ( 
.A(n_5265),
.B(n_483),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_5269),
.Y(n_5374)
);

INVxp67_ASAP7_75t_L g5375 ( 
.A(n_5301),
.Y(n_5375)
);

OR2x6_ASAP7_75t_L g5376 ( 
.A(n_5306),
.B(n_484),
.Y(n_5376)
);

AND2x2_ASAP7_75t_L g5377 ( 
.A(n_5262),
.B(n_485),
.Y(n_5377)
);

OAI31xp33_ASAP7_75t_SL g5378 ( 
.A1(n_5288),
.A2(n_5296),
.A3(n_5316),
.B(n_5312),
.Y(n_5378)
);

AND2x4_ASAP7_75t_L g5379 ( 
.A(n_5272),
.B(n_485),
.Y(n_5379)
);

INVx2_ASAP7_75t_L g5380 ( 
.A(n_5278),
.Y(n_5380)
);

BUFx2_ASAP7_75t_L g5381 ( 
.A(n_5277),
.Y(n_5381)
);

AOI221xp5_ASAP7_75t_L g5382 ( 
.A1(n_5252),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.C(n_488),
.Y(n_5382)
);

INVx2_ASAP7_75t_SL g5383 ( 
.A(n_5300),
.Y(n_5383)
);

AND2x2_ASAP7_75t_L g5384 ( 
.A(n_5309),
.B(n_486),
.Y(n_5384)
);

OR2x2_ASAP7_75t_L g5385 ( 
.A(n_5308),
.B(n_487),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_5310),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_5263),
.Y(n_5387)
);

AND2x2_ASAP7_75t_L g5388 ( 
.A(n_5307),
.B(n_487),
.Y(n_5388)
);

NAND2xp33_ASAP7_75t_L g5389 ( 
.A(n_5318),
.B(n_488),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_5263),
.Y(n_5390)
);

OAI22xp5_ASAP7_75t_L g5391 ( 
.A1(n_5308),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5263),
.Y(n_5392)
);

INVx2_ASAP7_75t_SL g5393 ( 
.A(n_5293),
.Y(n_5393)
);

BUFx2_ASAP7_75t_L g5394 ( 
.A(n_5286),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5263),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_L g5396 ( 
.A(n_5308),
.B(n_489),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5310),
.Y(n_5397)
);

AOI33xp33_ASAP7_75t_L g5398 ( 
.A1(n_5260),
.A2(n_492),
.A3(n_494),
.B1(n_489),
.B2(n_490),
.B3(n_493),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5263),
.Y(n_5399)
);

CKINVDCx5p33_ASAP7_75t_R g5400 ( 
.A(n_5301),
.Y(n_5400)
);

AND2x2_ASAP7_75t_L g5401 ( 
.A(n_5307),
.B(n_490),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5263),
.Y(n_5402)
);

OR2x2_ASAP7_75t_L g5403 ( 
.A(n_5308),
.B(n_492),
.Y(n_5403)
);

INVx2_ASAP7_75t_SL g5404 ( 
.A(n_5293),
.Y(n_5404)
);

AND2x2_ASAP7_75t_L g5405 ( 
.A(n_5307),
.B(n_492),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_5310),
.Y(n_5406)
);

CKINVDCx5p33_ASAP7_75t_R g5407 ( 
.A(n_5301),
.Y(n_5407)
);

NAND3xp33_ASAP7_75t_L g5408 ( 
.A(n_5264),
.B(n_493),
.C(n_494),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5329),
.Y(n_5409)
);

AND2x4_ASAP7_75t_L g5410 ( 
.A(n_5375),
.B(n_494),
.Y(n_5410)
);

AND2x2_ASAP7_75t_L g5411 ( 
.A(n_5348),
.B(n_5320),
.Y(n_5411)
);

NAND2xp5_ASAP7_75t_L g5412 ( 
.A(n_5371),
.B(n_495),
.Y(n_5412)
);

AND2x2_ASAP7_75t_L g5413 ( 
.A(n_5393),
.B(n_495),
.Y(n_5413)
);

HB1xp67_ASAP7_75t_L g5414 ( 
.A(n_5321),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5343),
.Y(n_5415)
);

NAND2x1p5_ASAP7_75t_L g5416 ( 
.A(n_5332),
.B(n_603),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5386),
.Y(n_5417)
);

AND2x2_ASAP7_75t_L g5418 ( 
.A(n_5404),
.B(n_495),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5388),
.Y(n_5419)
);

AND2x2_ASAP7_75t_L g5420 ( 
.A(n_5397),
.B(n_496),
.Y(n_5420)
);

NOR2x1_ASAP7_75t_L g5421 ( 
.A(n_5408),
.B(n_496),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5401),
.Y(n_5422)
);

AND2x2_ASAP7_75t_L g5423 ( 
.A(n_5406),
.B(n_496),
.Y(n_5423)
);

INVx2_ASAP7_75t_SL g5424 ( 
.A(n_5400),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5405),
.Y(n_5425)
);

AND2x2_ASAP7_75t_L g5426 ( 
.A(n_5394),
.B(n_497),
.Y(n_5426)
);

AND2x2_ASAP7_75t_L g5427 ( 
.A(n_5333),
.B(n_497),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_5356),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_5396),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_5341),
.Y(n_5430)
);

OR2x2_ASAP7_75t_SL g5431 ( 
.A(n_5374),
.B(n_497),
.Y(n_5431)
);

NOR2xp33_ASAP7_75t_L g5432 ( 
.A(n_5407),
.B(n_498),
.Y(n_5432)
);

AND2x2_ASAP7_75t_L g5433 ( 
.A(n_5328),
.B(n_498),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_5373),
.Y(n_5434)
);

AND2x2_ASAP7_75t_L g5435 ( 
.A(n_5327),
.B(n_498),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_5364),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5324),
.B(n_499),
.Y(n_5437)
);

OR2x2_ASAP7_75t_L g5438 ( 
.A(n_5336),
.B(n_499),
.Y(n_5438)
);

INVx1_ASAP7_75t_SL g5439 ( 
.A(n_5344),
.Y(n_5439)
);

AND2x2_ASAP7_75t_L g5440 ( 
.A(n_5324),
.B(n_500),
.Y(n_5440)
);

AND2x2_ASAP7_75t_L g5441 ( 
.A(n_5355),
.B(n_500),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_5387),
.Y(n_5442)
);

INVx2_ASAP7_75t_L g5443 ( 
.A(n_5372),
.Y(n_5443)
);

AND2x2_ASAP7_75t_L g5444 ( 
.A(n_5355),
.B(n_500),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_5366),
.Y(n_5445)
);

INVx1_ASAP7_75t_L g5446 ( 
.A(n_5390),
.Y(n_5446)
);

NOR2xp33_ASAP7_75t_L g5447 ( 
.A(n_5319),
.B(n_501),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5392),
.Y(n_5448)
);

AND2x2_ASAP7_75t_SL g5449 ( 
.A(n_5381),
.B(n_501),
.Y(n_5449)
);

NAND3xp33_ASAP7_75t_L g5450 ( 
.A(n_5339),
.B(n_501),
.C(n_502),
.Y(n_5450)
);

AND2x2_ASAP7_75t_L g5451 ( 
.A(n_5355),
.B(n_502),
.Y(n_5451)
);

OR2x2_ASAP7_75t_L g5452 ( 
.A(n_5337),
.B(n_502),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5395),
.Y(n_5453)
);

NAND2x1p5_ASAP7_75t_L g5454 ( 
.A(n_5379),
.B(n_604),
.Y(n_5454)
);

HB1xp67_ASAP7_75t_L g5455 ( 
.A(n_5399),
.Y(n_5455)
);

OR2x2_ASAP7_75t_L g5456 ( 
.A(n_5335),
.B(n_5325),
.Y(n_5456)
);

OR2x2_ASAP7_75t_L g5457 ( 
.A(n_5326),
.B(n_503),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_5402),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5330),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5359),
.Y(n_5460)
);

INVx1_ASAP7_75t_SL g5461 ( 
.A(n_5377),
.Y(n_5461)
);

AND2x2_ASAP7_75t_L g5462 ( 
.A(n_5349),
.B(n_503),
.Y(n_5462)
);

AND2x2_ASAP7_75t_L g5463 ( 
.A(n_5349),
.B(n_504),
.Y(n_5463)
);

AND2x2_ASAP7_75t_L g5464 ( 
.A(n_5383),
.B(n_504),
.Y(n_5464)
);

OR2x2_ASAP7_75t_L g5465 ( 
.A(n_5385),
.B(n_504),
.Y(n_5465)
);

AND2x2_ASAP7_75t_SL g5466 ( 
.A(n_5389),
.B(n_505),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_5322),
.Y(n_5467)
);

OR2x2_ASAP7_75t_L g5468 ( 
.A(n_5403),
.B(n_505),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5345),
.Y(n_5469)
);

AND2x2_ASAP7_75t_L g5470 ( 
.A(n_5379),
.B(n_505),
.Y(n_5470)
);

AND2x2_ASAP7_75t_L g5471 ( 
.A(n_5369),
.B(n_506),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_L g5472 ( 
.A(n_5447),
.B(n_5323),
.Y(n_5472)
);

AND2x2_ASAP7_75t_L g5473 ( 
.A(n_5424),
.B(n_5338),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5414),
.Y(n_5474)
);

OR2x2_ASAP7_75t_L g5475 ( 
.A(n_5412),
.B(n_5360),
.Y(n_5475)
);

HB1xp67_ASAP7_75t_L g5476 ( 
.A(n_5455),
.Y(n_5476)
);

INVx2_ASAP7_75t_L g5477 ( 
.A(n_5411),
.Y(n_5477)
);

XOR2x2_ASAP7_75t_L g5478 ( 
.A(n_5466),
.B(n_5382),
.Y(n_5478)
);

AND2x2_ASAP7_75t_L g5479 ( 
.A(n_5464),
.B(n_5350),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5415),
.Y(n_5480)
);

XNOR2xp5_ASAP7_75t_L g5481 ( 
.A(n_5433),
.B(n_5384),
.Y(n_5481)
);

INVx4_ASAP7_75t_L g5482 ( 
.A(n_5410),
.Y(n_5482)
);

XNOR2xp5_ASAP7_75t_L g5483 ( 
.A(n_5416),
.B(n_5334),
.Y(n_5483)
);

INVxp67_ASAP7_75t_L g5484 ( 
.A(n_5432),
.Y(n_5484)
);

AND2x2_ASAP7_75t_SL g5485 ( 
.A(n_5449),
.B(n_5398),
.Y(n_5485)
);

AND2x2_ASAP7_75t_L g5486 ( 
.A(n_5417),
.B(n_5370),
.Y(n_5486)
);

INVx1_ASAP7_75t_SL g5487 ( 
.A(n_5439),
.Y(n_5487)
);

AND2x2_ASAP7_75t_L g5488 ( 
.A(n_5426),
.B(n_5351),
.Y(n_5488)
);

BUFx2_ASAP7_75t_SL g5489 ( 
.A(n_5410),
.Y(n_5489)
);

NOR2xp33_ASAP7_75t_R g5490 ( 
.A(n_5413),
.B(n_5340),
.Y(n_5490)
);

NAND2xp5_ASAP7_75t_L g5491 ( 
.A(n_5435),
.B(n_5347),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5462),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5463),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5415),
.Y(n_5494)
);

NAND2xp5_ASAP7_75t_L g5495 ( 
.A(n_5461),
.B(n_5378),
.Y(n_5495)
);

INVx2_ASAP7_75t_L g5496 ( 
.A(n_5441),
.Y(n_5496)
);

INVx2_ASAP7_75t_L g5497 ( 
.A(n_5444),
.Y(n_5497)
);

NAND2xp5_ASAP7_75t_L g5498 ( 
.A(n_5460),
.B(n_5342),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_5434),
.B(n_5354),
.Y(n_5499)
);

NAND3xp33_ASAP7_75t_L g5500 ( 
.A(n_5409),
.B(n_5391),
.C(n_5368),
.Y(n_5500)
);

AND2x2_ASAP7_75t_L g5501 ( 
.A(n_5420),
.B(n_5358),
.Y(n_5501)
);

OR2x2_ASAP7_75t_L g5502 ( 
.A(n_5457),
.B(n_5331),
.Y(n_5502)
);

AOI22xp5_ASAP7_75t_L g5503 ( 
.A1(n_5428),
.A2(n_5376),
.B1(n_5362),
.B2(n_5380),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_5419),
.B(n_5361),
.Y(n_5504)
);

XOR2xp5_ASAP7_75t_L g5505 ( 
.A(n_5450),
.B(n_5352),
.Y(n_5505)
);

OR2x2_ASAP7_75t_L g5506 ( 
.A(n_5431),
.B(n_5357),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5451),
.Y(n_5507)
);

XNOR2xp5_ASAP7_75t_L g5508 ( 
.A(n_5454),
.B(n_5376),
.Y(n_5508)
);

NOR2x1p5_ASAP7_75t_L g5509 ( 
.A(n_5456),
.B(n_5409),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_5418),
.Y(n_5510)
);

NAND4xp75_ASAP7_75t_SL g5511 ( 
.A(n_5423),
.B(n_5353),
.C(n_5346),
.D(n_5365),
.Y(n_5511)
);

NAND4xp75_ASAP7_75t_L g5512 ( 
.A(n_5421),
.B(n_5367),
.C(n_5363),
.D(n_508),
.Y(n_5512)
);

XOR2xp5_ASAP7_75t_L g5513 ( 
.A(n_5427),
.B(n_506),
.Y(n_5513)
);

AND2x4_ASAP7_75t_L g5514 ( 
.A(n_5430),
.B(n_509),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_5436),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5437),
.Y(n_5516)
);

NOR4xp25_ASAP7_75t_L g5517 ( 
.A(n_5459),
.B(n_510),
.C(n_507),
.D(n_509),
.Y(n_5517)
);

AND2x2_ASAP7_75t_L g5518 ( 
.A(n_5440),
.B(n_507),
.Y(n_5518)
);

NAND2xp5_ASAP7_75t_L g5519 ( 
.A(n_5422),
.B(n_510),
.Y(n_5519)
);

AND2x2_ASAP7_75t_L g5520 ( 
.A(n_5425),
.B(n_510),
.Y(n_5520)
);

NOR3xp33_ASAP7_75t_SL g5521 ( 
.A(n_5429),
.B(n_511),
.C(n_512),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_5443),
.Y(n_5522)
);

AND2x2_ASAP7_75t_L g5523 ( 
.A(n_5471),
.B(n_511),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_5469),
.B(n_511),
.Y(n_5524)
);

INVxp67_ASAP7_75t_SL g5525 ( 
.A(n_5465),
.Y(n_5525)
);

AND2x2_ASAP7_75t_L g5526 ( 
.A(n_5469),
.B(n_513),
.Y(n_5526)
);

AND2x2_ASAP7_75t_L g5527 ( 
.A(n_5470),
.B(n_513),
.Y(n_5527)
);

INVx2_ASAP7_75t_SL g5528 ( 
.A(n_5468),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_5442),
.Y(n_5529)
);

NAND4xp75_ASAP7_75t_SL g5530 ( 
.A(n_5442),
.B(n_516),
.C(n_514),
.D(n_515),
.Y(n_5530)
);

NAND3xp33_ASAP7_75t_L g5531 ( 
.A(n_5445),
.B(n_514),
.C(n_515),
.Y(n_5531)
);

NAND4xp75_ASAP7_75t_SL g5532 ( 
.A(n_5446),
.B(n_517),
.C(n_515),
.D(n_516),
.Y(n_5532)
);

HB1xp67_ASAP7_75t_L g5533 ( 
.A(n_5446),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5448),
.Y(n_5534)
);

INVxp67_ASAP7_75t_L g5535 ( 
.A(n_5438),
.Y(n_5535)
);

INVxp67_ASAP7_75t_L g5536 ( 
.A(n_5452),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5448),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_5453),
.Y(n_5538)
);

XNOR2xp5_ASAP7_75t_L g5539 ( 
.A(n_5458),
.B(n_516),
.Y(n_5539)
);

NAND4xp75_ASAP7_75t_SL g5540 ( 
.A(n_5467),
.B(n_520),
.C(n_518),
.D(n_519),
.Y(n_5540)
);

XOR2x2_ASAP7_75t_L g5541 ( 
.A(n_5467),
.B(n_518),
.Y(n_5541)
);

NOR3xp33_ASAP7_75t_SL g5542 ( 
.A(n_5447),
.B(n_518),
.C(n_519),
.Y(n_5542)
);

AOI211xp5_ASAP7_75t_SL g5543 ( 
.A1(n_5447),
.A2(n_522),
.B(n_520),
.C(n_521),
.Y(n_5543)
);

NOR2x1_ASAP7_75t_L g5544 ( 
.A(n_5447),
.B(n_520),
.Y(n_5544)
);

XNOR2xp5_ASAP7_75t_L g5545 ( 
.A(n_5424),
.B(n_521),
.Y(n_5545)
);

BUFx3_ASAP7_75t_L g5546 ( 
.A(n_5411),
.Y(n_5546)
);

XNOR2x2_ASAP7_75t_L g5547 ( 
.A(n_5411),
.B(n_522),
.Y(n_5547)
);

NAND3xp33_ASAP7_75t_L g5548 ( 
.A(n_5447),
.B(n_522),
.C(n_523),
.Y(n_5548)
);

AND2x2_ASAP7_75t_L g5549 ( 
.A(n_5546),
.B(n_523),
.Y(n_5549)
);

AOI21xp5_ASAP7_75t_L g5550 ( 
.A1(n_5472),
.A2(n_5495),
.B(n_5508),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5476),
.Y(n_5551)
);

NAND2x1p5_ASAP7_75t_L g5552 ( 
.A(n_5482),
.B(n_523),
.Y(n_5552)
);

INVx2_ASAP7_75t_L g5553 ( 
.A(n_5477),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5474),
.Y(n_5554)
);

AOI22xp5_ASAP7_75t_L g5555 ( 
.A1(n_5485),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5515),
.Y(n_5556)
);

OR2x2_ASAP7_75t_L g5557 ( 
.A(n_5487),
.B(n_524),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5522),
.Y(n_5558)
);

AND2x4_ASAP7_75t_L g5559 ( 
.A(n_5473),
.B(n_524),
.Y(n_5559)
);

AND2x2_ASAP7_75t_L g5560 ( 
.A(n_5479),
.B(n_526),
.Y(n_5560)
);

OR2x2_ASAP7_75t_L g5561 ( 
.A(n_5498),
.B(n_5500),
.Y(n_5561)
);

INVxp67_ASAP7_75t_L g5562 ( 
.A(n_5489),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_5489),
.Y(n_5563)
);

OR2x2_ASAP7_75t_L g5564 ( 
.A(n_5528),
.B(n_526),
.Y(n_5564)
);

OAI22xp33_ASAP7_75t_L g5565 ( 
.A1(n_5503),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_L g5566 ( 
.A(n_5481),
.B(n_527),
.Y(n_5566)
);

NAND2xp67_ASAP7_75t_L g5567 ( 
.A(n_5486),
.B(n_527),
.Y(n_5567)
);

AND2x2_ASAP7_75t_L g5568 ( 
.A(n_5501),
.B(n_528),
.Y(n_5568)
);

INVx4_ASAP7_75t_L g5569 ( 
.A(n_5482),
.Y(n_5569)
);

INVxp67_ASAP7_75t_L g5570 ( 
.A(n_5523),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5533),
.Y(n_5571)
);

AOI22xp5_ASAP7_75t_L g5572 ( 
.A1(n_5483),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_5572)
);

AND2x2_ASAP7_75t_L g5573 ( 
.A(n_5488),
.B(n_529),
.Y(n_5573)
);

NOR2x1_ASAP7_75t_L g5574 ( 
.A(n_5512),
.B(n_530),
.Y(n_5574)
);

AND2x2_ASAP7_75t_L g5575 ( 
.A(n_5520),
.B(n_531),
.Y(n_5575)
);

OR2x2_ASAP7_75t_L g5576 ( 
.A(n_5525),
.B(n_531),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_5543),
.B(n_532),
.Y(n_5577)
);

OR2x2_ASAP7_75t_L g5578 ( 
.A(n_5524),
.B(n_532),
.Y(n_5578)
);

OR2x2_ASAP7_75t_L g5579 ( 
.A(n_5519),
.B(n_532),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5514),
.Y(n_5580)
);

INVx2_ASAP7_75t_L g5581 ( 
.A(n_5514),
.Y(n_5581)
);

AND2x2_ASAP7_75t_L g5582 ( 
.A(n_5526),
.B(n_533),
.Y(n_5582)
);

NAND2xp5_ASAP7_75t_L g5583 ( 
.A(n_5545),
.B(n_533),
.Y(n_5583)
);

INVxp67_ASAP7_75t_SL g5584 ( 
.A(n_5484),
.Y(n_5584)
);

AND2x4_ASAP7_75t_L g5585 ( 
.A(n_5496),
.B(n_533),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_SL g5586 ( 
.A(n_5544),
.B(n_534),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5518),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_L g5588 ( 
.A(n_5517),
.B(n_534),
.Y(n_5588)
);

NAND2x1p5_ASAP7_75t_L g5589 ( 
.A(n_5527),
.B(n_535),
.Y(n_5589)
);

AOI22xp5_ASAP7_75t_L g5590 ( 
.A1(n_5478),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5480),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5494),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_5492),
.B(n_5493),
.Y(n_5593)
);

NAND2x1_ASAP7_75t_L g5594 ( 
.A(n_5497),
.B(n_535),
.Y(n_5594)
);

AND2x2_ASAP7_75t_L g5595 ( 
.A(n_5509),
.B(n_536),
.Y(n_5595)
);

NAND2xp5_ASAP7_75t_L g5596 ( 
.A(n_5510),
.B(n_537),
.Y(n_5596)
);

NOR2xp67_ASAP7_75t_L g5597 ( 
.A(n_5516),
.B(n_5506),
.Y(n_5597)
);

INVx1_ASAP7_75t_SL g5598 ( 
.A(n_5530),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5507),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_5539),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5505),
.B(n_537),
.Y(n_5601)
);

AND2x2_ASAP7_75t_SL g5602 ( 
.A(n_5475),
.B(n_538),
.Y(n_5602)
);

NAND2xp5_ASAP7_75t_L g5603 ( 
.A(n_5542),
.B(n_538),
.Y(n_5603)
);

OR4x1_ASAP7_75t_L g5604 ( 
.A(n_5529),
.B(n_5537),
.C(n_5534),
.D(n_5547),
.Y(n_5604)
);

AND2x4_ASAP7_75t_L g5605 ( 
.A(n_5521),
.B(n_538),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5504),
.Y(n_5606)
);

NAND2xp5_ASAP7_75t_L g5607 ( 
.A(n_5513),
.B(n_5535),
.Y(n_5607)
);

AND2x4_ASAP7_75t_L g5608 ( 
.A(n_5536),
.B(n_539),
.Y(n_5608)
);

NOR2xp33_ASAP7_75t_L g5609 ( 
.A(n_5491),
.B(n_539),
.Y(n_5609)
);

NAND2x1p5_ASAP7_75t_L g5610 ( 
.A(n_5502),
.B(n_540),
.Y(n_5610)
);

AND2x2_ASAP7_75t_L g5611 ( 
.A(n_5490),
.B(n_540),
.Y(n_5611)
);

NAND2xp5_ASAP7_75t_L g5612 ( 
.A(n_5541),
.B(n_540),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5499),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5538),
.Y(n_5614)
);

OR2x2_ASAP7_75t_L g5615 ( 
.A(n_5531),
.B(n_542),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5548),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5532),
.Y(n_5617)
);

NOR2xp33_ASAP7_75t_L g5618 ( 
.A(n_5511),
.B(n_5540),
.Y(n_5618)
);

CKINVDCx16_ASAP7_75t_R g5619 ( 
.A(n_5569),
.Y(n_5619)
);

OAI21xp33_ASAP7_75t_SL g5620 ( 
.A1(n_5563),
.A2(n_542),
.B(n_543),
.Y(n_5620)
);

OAI22xp33_ASAP7_75t_L g5621 ( 
.A1(n_5562),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_5621)
);

OAI21xp33_ASAP7_75t_L g5622 ( 
.A1(n_5561),
.A2(n_544),
.B(n_545),
.Y(n_5622)
);

OAI21xp33_ASAP7_75t_L g5623 ( 
.A1(n_5618),
.A2(n_544),
.B(n_546),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5549),
.Y(n_5624)
);

INVx1_ASAP7_75t_SL g5625 ( 
.A(n_5585),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5557),
.Y(n_5626)
);

INVxp67_ASAP7_75t_SL g5627 ( 
.A(n_5552),
.Y(n_5627)
);

INVx2_ASAP7_75t_L g5628 ( 
.A(n_5553),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5581),
.Y(n_5629)
);

AND2x2_ASAP7_75t_L g5630 ( 
.A(n_5560),
.B(n_546),
.Y(n_5630)
);

XNOR2x1_ASAP7_75t_L g5631 ( 
.A(n_5574),
.B(n_546),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_5595),
.Y(n_5632)
);

AOI21xp33_ASAP7_75t_L g5633 ( 
.A1(n_5556),
.A2(n_547),
.B(n_548),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_5558),
.Y(n_5634)
);

INVx2_ASAP7_75t_L g5635 ( 
.A(n_5585),
.Y(n_5635)
);

AOI22xp5_ASAP7_75t_L g5636 ( 
.A1(n_5598),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.Y(n_5636)
);

OAI21xp5_ASAP7_75t_L g5637 ( 
.A1(n_5550),
.A2(n_548),
.B(n_549),
.Y(n_5637)
);

OR2x2_ASAP7_75t_L g5638 ( 
.A(n_5601),
.B(n_549),
.Y(n_5638)
);

OAI21xp5_ASAP7_75t_L g5639 ( 
.A1(n_5597),
.A2(n_550),
.B(n_551),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_5605),
.B(n_551),
.Y(n_5640)
);

OAI21xp5_ASAP7_75t_L g5641 ( 
.A1(n_5570),
.A2(n_552),
.B(n_553),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_5611),
.Y(n_5642)
);

AOI22xp5_ASAP7_75t_L g5643 ( 
.A1(n_5617),
.A2(n_5609),
.B1(n_5573),
.B2(n_5584),
.Y(n_5643)
);

INVxp67_ASAP7_75t_L g5644 ( 
.A(n_5575),
.Y(n_5644)
);

OR4x1_ASAP7_75t_L g5645 ( 
.A(n_5551),
.B(n_554),
.C(n_552),
.D(n_553),
.Y(n_5645)
);

NAND2xp5_ASAP7_75t_L g5646 ( 
.A(n_5559),
.B(n_552),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5564),
.Y(n_5647)
);

INVx2_ASAP7_75t_SL g5648 ( 
.A(n_5580),
.Y(n_5648)
);

INVx1_ASAP7_75t_SL g5649 ( 
.A(n_5608),
.Y(n_5649)
);

OA21x2_ASAP7_75t_L g5650 ( 
.A1(n_5566),
.A2(n_553),
.B(n_554),
.Y(n_5650)
);

OAI211xp5_ASAP7_75t_SL g5651 ( 
.A1(n_5554),
.A2(n_564),
.B(n_572),
.C(n_556),
.Y(n_5651)
);

NAND3xp33_ASAP7_75t_SL g5652 ( 
.A(n_5555),
.B(n_5590),
.C(n_5572),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_5582),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5615),
.Y(n_5654)
);

NAND2xp5_ASAP7_75t_L g5655 ( 
.A(n_5568),
.B(n_556),
.Y(n_5655)
);

AOI22xp5_ASAP7_75t_L g5656 ( 
.A1(n_5600),
.A2(n_5616),
.B1(n_5612),
.B2(n_5565),
.Y(n_5656)
);

OAI221xp5_ASAP7_75t_L g5657 ( 
.A1(n_5594),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.C(n_560),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5610),
.Y(n_5658)
);

O2A1O1Ixp33_ASAP7_75t_L g5659 ( 
.A1(n_5607),
.A2(n_5588),
.B(n_5586),
.C(n_5571),
.Y(n_5659)
);

NAND2x1p5_ASAP7_75t_L g5660 ( 
.A(n_5578),
.B(n_557),
.Y(n_5660)
);

NAND3xp33_ASAP7_75t_L g5661 ( 
.A(n_5576),
.B(n_5614),
.C(n_5577),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5579),
.Y(n_5662)
);

NAND3xp33_ASAP7_75t_L g5663 ( 
.A(n_5596),
.B(n_557),
.C(n_558),
.Y(n_5663)
);

NAND3xp33_ASAP7_75t_L g5664 ( 
.A(n_5606),
.B(n_558),
.C(n_559),
.Y(n_5664)
);

AOI22xp33_ASAP7_75t_L g5665 ( 
.A1(n_5613),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.Y(n_5665)
);

OAI22xp5_ASAP7_75t_L g5666 ( 
.A1(n_5587),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.Y(n_5666)
);

A2O1A1Ixp33_ASAP7_75t_L g5667 ( 
.A1(n_5599),
.A2(n_565),
.B(n_563),
.C(n_564),
.Y(n_5667)
);

INVxp67_ASAP7_75t_L g5668 ( 
.A(n_5583),
.Y(n_5668)
);

OAI21xp33_ASAP7_75t_L g5669 ( 
.A1(n_5567),
.A2(n_563),
.B(n_564),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_5593),
.Y(n_5670)
);

INVxp67_ASAP7_75t_L g5671 ( 
.A(n_5603),
.Y(n_5671)
);

AOI21xp33_ASAP7_75t_L g5672 ( 
.A1(n_5602),
.A2(n_565),
.B(n_566),
.Y(n_5672)
);

AOI21xp5_ASAP7_75t_L g5673 ( 
.A1(n_5591),
.A2(n_5592),
.B(n_5589),
.Y(n_5673)
);

OAI21xp33_ASAP7_75t_SL g5674 ( 
.A1(n_5604),
.A2(n_565),
.B(n_566),
.Y(n_5674)
);

AOI22xp5_ASAP7_75t_L g5675 ( 
.A1(n_5598),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5563),
.Y(n_5676)
);

A2O1A1Ixp33_ASAP7_75t_L g5677 ( 
.A1(n_5618),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_5677)
);

NAND2xp5_ASAP7_75t_L g5678 ( 
.A(n_5563),
.B(n_567),
.Y(n_5678)
);

INVx2_ASAP7_75t_L g5679 ( 
.A(n_5563),
.Y(n_5679)
);

OAI22xp33_ASAP7_75t_L g5680 ( 
.A1(n_5569),
.A2(n_570),
.B1(n_568),
.B2(n_569),
.Y(n_5680)
);

INVx2_ASAP7_75t_SL g5681 ( 
.A(n_5563),
.Y(n_5681)
);

XNOR2x1_ASAP7_75t_L g5682 ( 
.A(n_5574),
.B(n_570),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5563),
.Y(n_5683)
);

AOI22xp33_ASAP7_75t_L g5684 ( 
.A1(n_5569),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_5563),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_5563),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5563),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5563),
.Y(n_5688)
);

INVx2_ASAP7_75t_L g5689 ( 
.A(n_5563),
.Y(n_5689)
);

OAI211xp5_ASAP7_75t_L g5690 ( 
.A1(n_5674),
.A2(n_573),
.B(n_571),
.C(n_572),
.Y(n_5690)
);

AOI22xp33_ASAP7_75t_SL g5691 ( 
.A1(n_5619),
.A2(n_575),
.B1(n_573),
.B2(n_574),
.Y(n_5691)
);

NOR2xp33_ASAP7_75t_L g5692 ( 
.A(n_5620),
.B(n_573),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5681),
.Y(n_5693)
);

AOI211xp5_ASAP7_75t_L g5694 ( 
.A1(n_5637),
.A2(n_574),
.B(n_576),
.C(n_604),
.Y(n_5694)
);

AND2x2_ASAP7_75t_L g5695 ( 
.A(n_5630),
.B(n_576),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_5679),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5686),
.Y(n_5697)
);

OAI31xp33_ASAP7_75t_L g5698 ( 
.A1(n_5631),
.A2(n_607),
.A3(n_605),
.B(n_606),
.Y(n_5698)
);

AND2x2_ASAP7_75t_L g5699 ( 
.A(n_5627),
.B(n_605),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_5689),
.Y(n_5700)
);

NAND2xp5_ASAP7_75t_L g5701 ( 
.A(n_5676),
.B(n_606),
.Y(n_5701)
);

NAND2xp5_ASAP7_75t_L g5702 ( 
.A(n_5683),
.B(n_607),
.Y(n_5702)
);

AO21x1_ASAP7_75t_L g5703 ( 
.A1(n_5685),
.A2(n_608),
.B(n_609),
.Y(n_5703)
);

AOI22xp33_ASAP7_75t_SL g5704 ( 
.A1(n_5687),
.A2(n_611),
.B1(n_608),
.B2(n_610),
.Y(n_5704)
);

NAND2xp5_ASAP7_75t_L g5705 ( 
.A(n_5688),
.B(n_610),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5640),
.Y(n_5706)
);

AOI221xp5_ASAP7_75t_L g5707 ( 
.A1(n_5652),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.C(n_614),
.Y(n_5707)
);

NOR2xp33_ASAP7_75t_L g5708 ( 
.A(n_5625),
.B(n_613),
.Y(n_5708)
);

OAI21xp5_ASAP7_75t_SL g5709 ( 
.A1(n_5682),
.A2(n_615),
.B(n_616),
.Y(n_5709)
);

AOI22xp5_ASAP7_75t_L g5710 ( 
.A1(n_5670),
.A2(n_619),
.B1(n_617),
.B2(n_618),
.Y(n_5710)
);

OAI32xp33_ASAP7_75t_L g5711 ( 
.A1(n_5628),
.A2(n_619),
.A3(n_617),
.B1(n_618),
.B2(n_620),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5678),
.Y(n_5712)
);

OR2x2_ASAP7_75t_L g5713 ( 
.A(n_5629),
.B(n_981),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5646),
.Y(n_5714)
);

AND2x2_ASAP7_75t_L g5715 ( 
.A(n_5649),
.B(n_620),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_5635),
.Y(n_5716)
);

INVx2_ASAP7_75t_SL g5717 ( 
.A(n_5648),
.Y(n_5717)
);

OAI22xp33_ASAP7_75t_L g5718 ( 
.A1(n_5643),
.A2(n_623),
.B1(n_621),
.B2(n_622),
.Y(n_5718)
);

AO21x1_ASAP7_75t_L g5719 ( 
.A1(n_5634),
.A2(n_621),
.B(n_622),
.Y(n_5719)
);

AND2x2_ASAP7_75t_L g5720 ( 
.A(n_5653),
.B(n_624),
.Y(n_5720)
);

AOI21xp5_ASAP7_75t_L g5721 ( 
.A1(n_5672),
.A2(n_625),
.B(n_626),
.Y(n_5721)
);

NOR2xp33_ASAP7_75t_L g5722 ( 
.A(n_5622),
.B(n_626),
.Y(n_5722)
);

AOI221xp5_ASAP7_75t_L g5723 ( 
.A1(n_5659),
.A2(n_629),
.B1(n_627),
.B2(n_628),
.C(n_630),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5660),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5655),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_5636),
.Y(n_5726)
);

INVx2_ASAP7_75t_SL g5727 ( 
.A(n_5658),
.Y(n_5727)
);

AND2x2_ASAP7_75t_L g5728 ( 
.A(n_5624),
.B(n_628),
.Y(n_5728)
);

NAND2xp5_ASAP7_75t_L g5729 ( 
.A(n_5684),
.B(n_629),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_5675),
.Y(n_5730)
);

OAI22xp5_ASAP7_75t_L g5731 ( 
.A1(n_5656),
.A2(n_633),
.B1(n_630),
.B2(n_631),
.Y(n_5731)
);

AND2x2_ASAP7_75t_L g5732 ( 
.A(n_5642),
.B(n_631),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5638),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5666),
.Y(n_5734)
);

AND2x2_ASAP7_75t_L g5735 ( 
.A(n_5644),
.B(n_633),
.Y(n_5735)
);

AND2x2_ASAP7_75t_L g5736 ( 
.A(n_5632),
.B(n_634),
.Y(n_5736)
);

NAND2xp5_ASAP7_75t_L g5737 ( 
.A(n_5680),
.B(n_634),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5647),
.Y(n_5738)
);

OAI21xp33_ASAP7_75t_L g5739 ( 
.A1(n_5654),
.A2(n_635),
.B(n_636),
.Y(n_5739)
);

INVx2_ASAP7_75t_SL g5740 ( 
.A(n_5716),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5699),
.Y(n_5741)
);

AOI22xp5_ASAP7_75t_L g5742 ( 
.A1(n_5717),
.A2(n_5623),
.B1(n_5669),
.B2(n_5626),
.Y(n_5742)
);

INVxp67_ASAP7_75t_L g5743 ( 
.A(n_5708),
.Y(n_5743)
);

OR2x2_ASAP7_75t_L g5744 ( 
.A(n_5693),
.B(n_5664),
.Y(n_5744)
);

INVx1_ASAP7_75t_SL g5745 ( 
.A(n_5713),
.Y(n_5745)
);

AOI22xp5_ASAP7_75t_L g5746 ( 
.A1(n_5727),
.A2(n_5671),
.B1(n_5661),
.B2(n_5668),
.Y(n_5746)
);

AOI211x1_ASAP7_75t_L g5747 ( 
.A1(n_5690),
.A2(n_5673),
.B(n_5639),
.C(n_5662),
.Y(n_5747)
);

AOI22xp5_ASAP7_75t_L g5748 ( 
.A1(n_5692),
.A2(n_5663),
.B1(n_5621),
.B2(n_5657),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5715),
.Y(n_5749)
);

O2A1O1Ixp33_ASAP7_75t_L g5750 ( 
.A1(n_5731),
.A2(n_5677),
.B(n_5667),
.C(n_5633),
.Y(n_5750)
);

AND2x2_ASAP7_75t_L g5751 ( 
.A(n_5695),
.B(n_5650),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5696),
.Y(n_5752)
);

OAI22xp5_ASAP7_75t_L g5753 ( 
.A1(n_5697),
.A2(n_5665),
.B1(n_5650),
.B2(n_5641),
.Y(n_5753)
);

NAND2xp5_ASAP7_75t_L g5754 ( 
.A(n_5691),
.B(n_5645),
.Y(n_5754)
);

INVx2_ASAP7_75t_L g5755 ( 
.A(n_5700),
.Y(n_5755)
);

OAI221xp5_ASAP7_75t_L g5756 ( 
.A1(n_5698),
.A2(n_5651),
.B1(n_639),
.B2(n_637),
.C(n_638),
.Y(n_5756)
);

XOR2x2_ASAP7_75t_L g5757 ( 
.A(n_5694),
.B(n_637),
.Y(n_5757)
);

INVx2_ASAP7_75t_L g5758 ( 
.A(n_5724),
.Y(n_5758)
);

INVx2_ASAP7_75t_SL g5759 ( 
.A(n_5738),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5703),
.Y(n_5760)
);

AND2x2_ASAP7_75t_L g5761 ( 
.A(n_5735),
.B(n_638),
.Y(n_5761)
);

NAND4xp25_ASAP7_75t_SL g5762 ( 
.A(n_5726),
.B(n_642),
.C(n_639),
.D(n_640),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5728),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5737),
.Y(n_5764)
);

AND2x2_ASAP7_75t_L g5765 ( 
.A(n_5720),
.B(n_640),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5719),
.Y(n_5766)
);

NAND3xp33_ASAP7_75t_L g5767 ( 
.A(n_5707),
.B(n_642),
.C(n_643),
.Y(n_5767)
);

INVxp67_ASAP7_75t_SL g5768 ( 
.A(n_5701),
.Y(n_5768)
);

AOI21xp33_ASAP7_75t_L g5769 ( 
.A1(n_5730),
.A2(n_5718),
.B(n_5705),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5736),
.Y(n_5770)
);

AND2x2_ASAP7_75t_L g5771 ( 
.A(n_5732),
.B(n_5730),
.Y(n_5771)
);

AOI22xp5_ASAP7_75t_L g5772 ( 
.A1(n_5734),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.Y(n_5772)
);

OAI221xp5_ASAP7_75t_L g5773 ( 
.A1(n_5709),
.A2(n_649),
.B1(n_647),
.B2(n_648),
.C(n_650),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5702),
.Y(n_5774)
);

INVxp67_ASAP7_75t_L g5775 ( 
.A(n_5722),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5733),
.Y(n_5776)
);

NAND2xp5_ASAP7_75t_L g5777 ( 
.A(n_5704),
.B(n_647),
.Y(n_5777)
);

AOI222xp33_ASAP7_75t_L g5778 ( 
.A1(n_5723),
.A2(n_651),
.B1(n_653),
.B2(n_648),
.C1(n_650),
.C2(n_652),
.Y(n_5778)
);

O2A1O1Ixp33_ASAP7_75t_L g5779 ( 
.A1(n_5729),
.A2(n_653),
.B(n_651),
.C(n_652),
.Y(n_5779)
);

NOR4xp25_ASAP7_75t_L g5780 ( 
.A(n_5706),
.B(n_5712),
.C(n_5714),
.D(n_5725),
.Y(n_5780)
);

INVxp67_ASAP7_75t_L g5781 ( 
.A(n_5721),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5711),
.Y(n_5782)
);

AND2x2_ASAP7_75t_L g5783 ( 
.A(n_5739),
.B(n_981),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5710),
.Y(n_5784)
);

AOI31xp33_ASAP7_75t_L g5785 ( 
.A1(n_5723),
.A2(n_658),
.A3(n_654),
.B(n_655),
.Y(n_5785)
);

AND2x2_ASAP7_75t_L g5786 ( 
.A(n_5699),
.B(n_979),
.Y(n_5786)
);

OR2x2_ASAP7_75t_L g5787 ( 
.A(n_5717),
.B(n_654),
.Y(n_5787)
);

NOR3xp33_ASAP7_75t_L g5788 ( 
.A(n_5762),
.B(n_655),
.C(n_660),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_5740),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5787),
.Y(n_5790)
);

NAND2xp5_ASAP7_75t_SL g5791 ( 
.A(n_5758),
.B(n_661),
.Y(n_5791)
);

INVx2_ASAP7_75t_L g5792 ( 
.A(n_5755),
.Y(n_5792)
);

AND2x2_ASAP7_75t_L g5793 ( 
.A(n_5786),
.B(n_662),
.Y(n_5793)
);

NOR2xp33_ASAP7_75t_L g5794 ( 
.A(n_5760),
.B(n_662),
.Y(n_5794)
);

OR2x2_ASAP7_75t_L g5795 ( 
.A(n_5744),
.B(n_663),
.Y(n_5795)
);

NOR2xp33_ASAP7_75t_L g5796 ( 
.A(n_5766),
.B(n_666),
.Y(n_5796)
);

AND2x2_ASAP7_75t_L g5797 ( 
.A(n_5765),
.B(n_668),
.Y(n_5797)
);

XNOR2x1_ASAP7_75t_L g5798 ( 
.A(n_5757),
.B(n_668),
.Y(n_5798)
);

AOI211xp5_ASAP7_75t_L g5799 ( 
.A1(n_5773),
.A2(n_5769),
.B(n_5756),
.C(n_5753),
.Y(n_5799)
);

NAND2xp5_ASAP7_75t_SL g5800 ( 
.A(n_5772),
.B(n_669),
.Y(n_5800)
);

OAI211xp5_ASAP7_75t_L g5801 ( 
.A1(n_5778),
.A2(n_671),
.B(n_669),
.C(n_670),
.Y(n_5801)
);

NAND2xp5_ASAP7_75t_L g5802 ( 
.A(n_5751),
.B(n_671),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_5761),
.B(n_5771),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5783),
.Y(n_5804)
);

NAND3xp33_ASAP7_75t_SL g5805 ( 
.A(n_5779),
.B(n_672),
.C(n_673),
.Y(n_5805)
);

XOR2x2_ASAP7_75t_L g5806 ( 
.A(n_5747),
.B(n_672),
.Y(n_5806)
);

INVx2_ASAP7_75t_L g5807 ( 
.A(n_5752),
.Y(n_5807)
);

NOR2xp33_ASAP7_75t_L g5808 ( 
.A(n_5754),
.B(n_674),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5777),
.Y(n_5809)
);

NAND2xp5_ASAP7_75t_SL g5810 ( 
.A(n_5748),
.B(n_675),
.Y(n_5810)
);

NOR3x1_ASAP7_75t_L g5811 ( 
.A(n_5767),
.B(n_675),
.C(n_676),
.Y(n_5811)
);

AOI21xp5_ASAP7_75t_L g5812 ( 
.A1(n_5750),
.A2(n_677),
.B(n_679),
.Y(n_5812)
);

OAI21xp5_ASAP7_75t_SL g5813 ( 
.A1(n_5785),
.A2(n_680),
.B(n_681),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5782),
.Y(n_5814)
);

INVx2_ASAP7_75t_SL g5815 ( 
.A(n_5776),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5742),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_5741),
.Y(n_5817)
);

AOI21xp5_ASAP7_75t_L g5818 ( 
.A1(n_5781),
.A2(n_682),
.B(n_683),
.Y(n_5818)
);

NOR2xp33_ASAP7_75t_L g5819 ( 
.A(n_5745),
.B(n_682),
.Y(n_5819)
);

NOR2xp33_ASAP7_75t_L g5820 ( 
.A(n_5749),
.B(n_684),
.Y(n_5820)
);

INVxp67_ASAP7_75t_L g5821 ( 
.A(n_5759),
.Y(n_5821)
);

NAND3xp33_ASAP7_75t_L g5822 ( 
.A(n_5746),
.B(n_685),
.C(n_686),
.Y(n_5822)
);

OAI21xp33_ASAP7_75t_L g5823 ( 
.A1(n_5780),
.A2(n_686),
.B(n_687),
.Y(n_5823)
);

NOR2xp33_ASAP7_75t_L g5824 ( 
.A(n_5784),
.B(n_687),
.Y(n_5824)
);

NOR2xp33_ASAP7_75t_SL g5825 ( 
.A(n_5743),
.B(n_688),
.Y(n_5825)
);

AND2x2_ASAP7_75t_L g5826 ( 
.A(n_5803),
.B(n_5763),
.Y(n_5826)
);

AOI22xp5_ASAP7_75t_L g5827 ( 
.A1(n_5789),
.A2(n_5764),
.B1(n_5770),
.B2(n_5775),
.Y(n_5827)
);

NAND3xp33_ASAP7_75t_L g5828 ( 
.A(n_5808),
.B(n_5764),
.C(n_5774),
.Y(n_5828)
);

OAI211xp5_ASAP7_75t_L g5829 ( 
.A1(n_5799),
.A2(n_5768),
.B(n_691),
.C(n_688),
.Y(n_5829)
);

AOI211x1_ASAP7_75t_L g5830 ( 
.A1(n_5812),
.A2(n_692),
.B(n_689),
.C(n_691),
.Y(n_5830)
);

AND2x2_ASAP7_75t_L g5831 ( 
.A(n_5797),
.B(n_692),
.Y(n_5831)
);

NAND3xp33_ASAP7_75t_L g5832 ( 
.A(n_5822),
.B(n_693),
.C(n_694),
.Y(n_5832)
);

AOI221xp5_ASAP7_75t_L g5833 ( 
.A1(n_5823),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.C(n_699),
.Y(n_5833)
);

AOI21xp5_ASAP7_75t_SL g5834 ( 
.A1(n_5823),
.A2(n_695),
.B(n_696),
.Y(n_5834)
);

AOI221xp5_ASAP7_75t_L g5835 ( 
.A1(n_5814),
.A2(n_701),
.B1(n_697),
.B2(n_700),
.C(n_702),
.Y(n_5835)
);

OAI311xp33_ASAP7_75t_L g5836 ( 
.A1(n_5813),
.A2(n_702),
.A3(n_700),
.B1(n_701),
.C1(n_703),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5792),
.Y(n_5837)
);

OAI221xp5_ASAP7_75t_L g5838 ( 
.A1(n_5788),
.A2(n_5821),
.B1(n_5816),
.B2(n_5815),
.C(n_5801),
.Y(n_5838)
);

OAI22xp5_ASAP7_75t_L g5839 ( 
.A1(n_5802),
.A2(n_706),
.B1(n_704),
.B2(n_705),
.Y(n_5839)
);

OAI21xp5_ASAP7_75t_L g5840 ( 
.A1(n_5818),
.A2(n_705),
.B(n_706),
.Y(n_5840)
);

NAND2xp33_ASAP7_75t_SL g5841 ( 
.A(n_5798),
.B(n_978),
.Y(n_5841)
);

NOR2xp33_ASAP7_75t_L g5842 ( 
.A(n_5805),
.B(n_708),
.Y(n_5842)
);

AOI22xp33_ASAP7_75t_L g5843 ( 
.A1(n_5807),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_5843)
);

NOR2xp33_ASAP7_75t_L g5844 ( 
.A(n_5825),
.B(n_709),
.Y(n_5844)
);

HB1xp67_ASAP7_75t_L g5845 ( 
.A(n_5795),
.Y(n_5845)
);

AOI221x1_ASAP7_75t_L g5846 ( 
.A1(n_5817),
.A2(n_5796),
.B1(n_5794),
.B2(n_5819),
.C(n_5824),
.Y(n_5846)
);

OAI221xp5_ASAP7_75t_SL g5847 ( 
.A1(n_5790),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.C(n_713),
.Y(n_5847)
);

NAND2xp5_ASAP7_75t_L g5848 ( 
.A(n_5793),
.B(n_712),
.Y(n_5848)
);

OAI32xp33_ASAP7_75t_L g5849 ( 
.A1(n_5820),
.A2(n_5804),
.A3(n_5809),
.B1(n_5810),
.B2(n_5791),
.Y(n_5849)
);

NOR3x1_ASAP7_75t_L g5850 ( 
.A(n_5800),
.B(n_713),
.C(n_714),
.Y(n_5850)
);

AOI221xp5_ASAP7_75t_L g5851 ( 
.A1(n_5806),
.A2(n_717),
.B1(n_715),
.B2(n_716),
.C(n_719),
.Y(n_5851)
);

AOI21xp5_ASAP7_75t_L g5852 ( 
.A1(n_5811),
.A2(n_715),
.B(n_716),
.Y(n_5852)
);

NAND2xp5_ASAP7_75t_L g5853 ( 
.A(n_5789),
.B(n_719),
.Y(n_5853)
);

NAND2xp5_ASAP7_75t_L g5854 ( 
.A(n_5789),
.B(n_720),
.Y(n_5854)
);

OAI21xp5_ASAP7_75t_SL g5855 ( 
.A1(n_5813),
.A2(n_721),
.B(n_722),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5789),
.Y(n_5856)
);

AOI21xp5_ASAP7_75t_L g5857 ( 
.A1(n_5812),
.A2(n_721),
.B(n_723),
.Y(n_5857)
);

OAI22x1_ASAP7_75t_L g5858 ( 
.A1(n_5837),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5856),
.Y(n_5859)
);

OAI22xp5_ASAP7_75t_L g5860 ( 
.A1(n_5838),
.A2(n_729),
.B1(n_727),
.B2(n_728),
.Y(n_5860)
);

INVx1_ASAP7_75t_SL g5861 ( 
.A(n_5853),
.Y(n_5861)
);

AOI22xp5_ASAP7_75t_L g5862 ( 
.A1(n_5842),
.A2(n_732),
.B1(n_730),
.B2(n_731),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5854),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5826),
.Y(n_5864)
);

INVxp33_ASAP7_75t_L g5865 ( 
.A(n_5844),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5848),
.Y(n_5866)
);

BUFx2_ASAP7_75t_L g5867 ( 
.A(n_5845),
.Y(n_5867)
);

AOI31xp33_ASAP7_75t_L g5868 ( 
.A1(n_5835),
.A2(n_733),
.A3(n_730),
.B(n_732),
.Y(n_5868)
);

INVx2_ASAP7_75t_L g5869 ( 
.A(n_5850),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5831),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_L g5871 ( 
.A(n_5852),
.B(n_733),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5839),
.Y(n_5872)
);

A2O1A1Ixp33_ASAP7_75t_SL g5873 ( 
.A1(n_5829),
.A2(n_737),
.B(n_734),
.C(n_735),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5830),
.Y(n_5874)
);

AOI22xp5_ASAP7_75t_L g5875 ( 
.A1(n_5855),
.A2(n_738),
.B1(n_735),
.B2(n_737),
.Y(n_5875)
);

OA22x2_ASAP7_75t_L g5876 ( 
.A1(n_5827),
.A2(n_740),
.B1(n_738),
.B2(n_739),
.Y(n_5876)
);

AND4x1_ASAP7_75t_L g5877 ( 
.A(n_5851),
.B(n_742),
.C(n_739),
.D(n_741),
.Y(n_5877)
);

AOI22xp5_ASAP7_75t_L g5878 ( 
.A1(n_5841),
.A2(n_5828),
.B1(n_5832),
.B2(n_5833),
.Y(n_5878)
);

NAND4xp25_ASAP7_75t_SL g5879 ( 
.A(n_5846),
.B(n_744),
.C(n_741),
.D(n_743),
.Y(n_5879)
);

AOI22xp5_ASAP7_75t_L g5880 ( 
.A1(n_5840),
.A2(n_746),
.B1(n_743),
.B2(n_745),
.Y(n_5880)
);

AOI221xp5_ASAP7_75t_L g5881 ( 
.A1(n_5860),
.A2(n_5847),
.B1(n_5849),
.B2(n_5834),
.C(n_5857),
.Y(n_5881)
);

AOI221xp5_ASAP7_75t_L g5882 ( 
.A1(n_5868),
.A2(n_5836),
.B1(n_5843),
.B2(n_749),
.C(n_747),
.Y(n_5882)
);

NAND2xp5_ASAP7_75t_L g5883 ( 
.A(n_5864),
.B(n_977),
.Y(n_5883)
);

AOI221xp5_ASAP7_75t_L g5884 ( 
.A1(n_5858),
.A2(n_749),
.B1(n_747),
.B2(n_748),
.C(n_750),
.Y(n_5884)
);

NOR3xp33_ASAP7_75t_L g5885 ( 
.A(n_5879),
.B(n_748),
.C(n_751),
.Y(n_5885)
);

OAI21xp5_ASAP7_75t_SL g5886 ( 
.A1(n_5875),
.A2(n_752),
.B(n_753),
.Y(n_5886)
);

O2A1O1Ixp33_ASAP7_75t_L g5887 ( 
.A1(n_5873),
.A2(n_754),
.B(n_752),
.C(n_753),
.Y(n_5887)
);

O2A1O1Ixp33_ASAP7_75t_L g5888 ( 
.A1(n_5871),
.A2(n_758),
.B(n_755),
.C(n_756),
.Y(n_5888)
);

AOI221xp5_ASAP7_75t_L g5889 ( 
.A1(n_5859),
.A2(n_760),
.B1(n_758),
.B2(n_759),
.C(n_761),
.Y(n_5889)
);

OAI221xp5_ASAP7_75t_SL g5890 ( 
.A1(n_5862),
.A2(n_762),
.B1(n_759),
.B2(n_761),
.C(n_763),
.Y(n_5890)
);

AOI22xp5_ASAP7_75t_L g5891 ( 
.A1(n_5874),
.A2(n_765),
.B1(n_762),
.B2(n_764),
.Y(n_5891)
);

AOI221xp5_ASAP7_75t_L g5892 ( 
.A1(n_5867),
.A2(n_766),
.B1(n_764),
.B2(n_765),
.C(n_767),
.Y(n_5892)
);

NAND3xp33_ASAP7_75t_SL g5893 ( 
.A(n_5880),
.B(n_767),
.C(n_768),
.Y(n_5893)
);

OAI21xp33_ASAP7_75t_L g5894 ( 
.A1(n_5865),
.A2(n_768),
.B(n_769),
.Y(n_5894)
);

NOR3xp33_ASAP7_75t_SL g5895 ( 
.A(n_5872),
.B(n_770),
.C(n_771),
.Y(n_5895)
);

OAI21xp5_ASAP7_75t_L g5896 ( 
.A1(n_5878),
.A2(n_771),
.B(n_772),
.Y(n_5896)
);

OAI211xp5_ASAP7_75t_SL g5897 ( 
.A1(n_5881),
.A2(n_5861),
.B(n_5863),
.C(n_5866),
.Y(n_5897)
);

AOI211xp5_ASAP7_75t_L g5898 ( 
.A1(n_5890),
.A2(n_5869),
.B(n_5870),
.C(n_5877),
.Y(n_5898)
);

HB1xp67_ASAP7_75t_L g5899 ( 
.A(n_5883),
.Y(n_5899)
);

AOI211x1_ASAP7_75t_SL g5900 ( 
.A1(n_5893),
.A2(n_5896),
.B(n_5882),
.C(n_5895),
.Y(n_5900)
);

NAND3x1_ASAP7_75t_SL g5901 ( 
.A(n_5884),
.B(n_5892),
.C(n_5889),
.Y(n_5901)
);

AOI211xp5_ASAP7_75t_L g5902 ( 
.A1(n_5894),
.A2(n_5887),
.B(n_5888),
.C(n_5886),
.Y(n_5902)
);

INVx2_ASAP7_75t_SL g5903 ( 
.A(n_5891),
.Y(n_5903)
);

OAI221xp5_ASAP7_75t_SL g5904 ( 
.A1(n_5885),
.A2(n_5876),
.B1(n_775),
.B2(n_773),
.C(n_774),
.Y(n_5904)
);

NAND4xp25_ASAP7_75t_SL g5905 ( 
.A(n_5881),
.B(n_776),
.C(n_773),
.D(n_775),
.Y(n_5905)
);

NAND3xp33_ASAP7_75t_SL g5906 ( 
.A(n_5881),
.B(n_777),
.C(n_778),
.Y(n_5906)
);

OAI211xp5_ASAP7_75t_L g5907 ( 
.A1(n_5881),
.A2(n_779),
.B(n_777),
.C(n_778),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5883),
.Y(n_5908)
);

NAND3xp33_ASAP7_75t_SL g5909 ( 
.A(n_5881),
.B(n_779),
.C(n_780),
.Y(n_5909)
);

OAI221xp5_ASAP7_75t_L g5910 ( 
.A1(n_5892),
.A2(n_783),
.B1(n_781),
.B2(n_782),
.C(n_784),
.Y(n_5910)
);

INVx1_ASAP7_75t_L g5911 ( 
.A(n_5883),
.Y(n_5911)
);

AND3x4_ASAP7_75t_L g5912 ( 
.A(n_5901),
.B(n_782),
.C(n_784),
.Y(n_5912)
);

O2A1O1Ixp33_ASAP7_75t_L g5913 ( 
.A1(n_5910),
.A2(n_787),
.B(n_785),
.C(n_786),
.Y(n_5913)
);

NOR2x1_ASAP7_75t_L g5914 ( 
.A(n_5906),
.B(n_785),
.Y(n_5914)
);

NOR2x1_ASAP7_75t_L g5915 ( 
.A(n_5909),
.B(n_5897),
.Y(n_5915)
);

OAI321xp33_ASAP7_75t_L g5916 ( 
.A1(n_5904),
.A2(n_977),
.A3(n_788),
.B1(n_790),
.B2(n_786),
.C(n_787),
.Y(n_5916)
);

NOR2xp33_ASAP7_75t_L g5917 ( 
.A(n_5907),
.B(n_789),
.Y(n_5917)
);

NAND2x1p5_ASAP7_75t_L g5918 ( 
.A(n_5903),
.B(n_789),
.Y(n_5918)
);

NAND3x1_ASAP7_75t_SL g5919 ( 
.A(n_5905),
.B(n_790),
.C(n_791),
.Y(n_5919)
);

NOR3xp33_ASAP7_75t_L g5920 ( 
.A(n_5898),
.B(n_792),
.C(n_793),
.Y(n_5920)
);

AND3x1_ASAP7_75t_L g5921 ( 
.A(n_5902),
.B(n_792),
.C(n_793),
.Y(n_5921)
);

XNOR2xp5_ASAP7_75t_L g5922 ( 
.A(n_5900),
.B(n_794),
.Y(n_5922)
);

HB1xp67_ASAP7_75t_L g5923 ( 
.A(n_5899),
.Y(n_5923)
);

AOI221xp5_ASAP7_75t_L g5924 ( 
.A1(n_5916),
.A2(n_5911),
.B1(n_5908),
.B2(n_796),
.C(n_794),
.Y(n_5924)
);

NOR3xp33_ASAP7_75t_L g5925 ( 
.A(n_5915),
.B(n_976),
.C(n_795),
.Y(n_5925)
);

NOR2xp33_ASAP7_75t_L g5926 ( 
.A(n_5922),
.B(n_796),
.Y(n_5926)
);

AOI31xp33_ASAP7_75t_L g5927 ( 
.A1(n_5918),
.A2(n_800),
.A3(n_797),
.B(n_798),
.Y(n_5927)
);

OR2x2_ASAP7_75t_L g5928 ( 
.A(n_5923),
.B(n_797),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5912),
.Y(n_5929)
);

NAND3x1_ASAP7_75t_L g5930 ( 
.A(n_5914),
.B(n_800),
.C(n_801),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5921),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_5920),
.B(n_802),
.Y(n_5932)
);

NOR2x1_ASAP7_75t_L g5933 ( 
.A(n_5917),
.B(n_803),
.Y(n_5933)
);

NOR3x1_ASAP7_75t_L g5934 ( 
.A(n_5919),
.B(n_804),
.C(n_805),
.Y(n_5934)
);

NOR3xp33_ASAP7_75t_SL g5935 ( 
.A(n_5913),
.B(n_804),
.C(n_805),
.Y(n_5935)
);

NOR2x1p5_ASAP7_75t_L g5936 ( 
.A(n_5922),
.B(n_806),
.Y(n_5936)
);

INVx1_ASAP7_75t_L g5937 ( 
.A(n_5922),
.Y(n_5937)
);

NAND2xp5_ASAP7_75t_L g5938 ( 
.A(n_5922),
.B(n_806),
.Y(n_5938)
);

AOI21xp5_ASAP7_75t_SL g5939 ( 
.A1(n_5913),
.A2(n_807),
.B(n_808),
.Y(n_5939)
);

NAND2x1p5_ASAP7_75t_L g5940 ( 
.A(n_5915),
.B(n_807),
.Y(n_5940)
);

AND2x4_ASAP7_75t_L g5941 ( 
.A(n_5923),
.B(n_808),
.Y(n_5941)
);

NOR2xp33_ASAP7_75t_L g5942 ( 
.A(n_5922),
.B(n_809),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5922),
.Y(n_5943)
);

NAND5xp2_ASAP7_75t_L g5944 ( 
.A(n_5926),
.B(n_812),
.C(n_810),
.D(n_811),
.E(n_813),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5932),
.Y(n_5945)
);

NAND3xp33_ASAP7_75t_SL g5946 ( 
.A(n_5925),
.B(n_813),
.C(n_814),
.Y(n_5946)
);

AOI21xp5_ASAP7_75t_L g5947 ( 
.A1(n_5939),
.A2(n_815),
.B(n_817),
.Y(n_5947)
);

INVxp67_ASAP7_75t_L g5948 ( 
.A(n_5942),
.Y(n_5948)
);

OAI211xp5_ASAP7_75t_SL g5949 ( 
.A1(n_5938),
.A2(n_820),
.B(n_818),
.C(n_819),
.Y(n_5949)
);

NOR3xp33_ASAP7_75t_L g5950 ( 
.A(n_5937),
.B(n_818),
.C(n_820),
.Y(n_5950)
);

NAND4xp25_ASAP7_75t_SL g5951 ( 
.A(n_5924),
.B(n_823),
.C(n_821),
.D(n_822),
.Y(n_5951)
);

NAND5xp2_ASAP7_75t_L g5952 ( 
.A(n_5943),
.B(n_823),
.C(n_821),
.D(n_822),
.E(n_824),
.Y(n_5952)
);

AOI21xp5_ASAP7_75t_L g5953 ( 
.A1(n_5927),
.A2(n_824),
.B(n_825),
.Y(n_5953)
);

AOI22xp5_ASAP7_75t_L g5954 ( 
.A1(n_5929),
.A2(n_829),
.B1(n_827),
.B2(n_828),
.Y(n_5954)
);

XNOR2xp5_ASAP7_75t_L g5955 ( 
.A(n_5954),
.B(n_5936),
.Y(n_5955)
);

AND3x4_ASAP7_75t_L g5956 ( 
.A(n_5950),
.B(n_5935),
.C(n_5933),
.Y(n_5956)
);

HB1xp67_ASAP7_75t_L g5957 ( 
.A(n_5951),
.Y(n_5957)
);

NAND2x1p5_ASAP7_75t_L g5958 ( 
.A(n_5945),
.B(n_5931),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5948),
.Y(n_5959)
);

XNOR2xp5_ASAP7_75t_L g5960 ( 
.A(n_5946),
.B(n_5930),
.Y(n_5960)
);

NOR2xp67_ASAP7_75t_L g5961 ( 
.A(n_5944),
.B(n_5928),
.Y(n_5961)
);

AOI21xp5_ASAP7_75t_L g5962 ( 
.A1(n_5947),
.A2(n_5941),
.B(n_5940),
.Y(n_5962)
);

AOI211xp5_ASAP7_75t_SL g5963 ( 
.A1(n_5961),
.A2(n_5949),
.B(n_5953),
.C(n_5952),
.Y(n_5963)
);

AOI22xp33_ASAP7_75t_L g5964 ( 
.A1(n_5959),
.A2(n_5934),
.B1(n_831),
.B2(n_829),
.Y(n_5964)
);

INVxp67_ASAP7_75t_SL g5965 ( 
.A(n_5958),
.Y(n_5965)
);

AOI22xp5_ASAP7_75t_L g5966 ( 
.A1(n_5956),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.Y(n_5966)
);

INVx3_ASAP7_75t_L g5967 ( 
.A(n_5965),
.Y(n_5967)
);

AOI31xp33_ASAP7_75t_L g5968 ( 
.A1(n_5963),
.A2(n_5960),
.A3(n_5955),
.B(n_5957),
.Y(n_5968)
);

NAND2xp5_ASAP7_75t_L g5969 ( 
.A(n_5967),
.B(n_5962),
.Y(n_5969)
);

AOI22xp33_ASAP7_75t_L g5970 ( 
.A1(n_5969),
.A2(n_5968),
.B1(n_5964),
.B2(n_5966),
.Y(n_5970)
);

AOI22xp5_ASAP7_75t_L g5971 ( 
.A1(n_5970),
.A2(n_833),
.B1(n_830),
.B2(n_832),
.Y(n_5971)
);

AOI22xp5_ASAP7_75t_L g5972 ( 
.A1(n_5971),
.A2(n_836),
.B1(n_834),
.B2(n_835),
.Y(n_5972)
);

OAI22xp5_ASAP7_75t_L g5973 ( 
.A1(n_5972),
.A2(n_838),
.B1(n_835),
.B2(n_837),
.Y(n_5973)
);

XNOR2xp5_ASAP7_75t_SL g5974 ( 
.A(n_5973),
.B(n_838),
.Y(n_5974)
);

AOI22xp33_ASAP7_75t_L g5975 ( 
.A1(n_5974),
.A2(n_841),
.B1(n_839),
.B2(n_840),
.Y(n_5975)
);

O2A1O1Ixp33_ASAP7_75t_L g5976 ( 
.A1(n_5975),
.A2(n_843),
.B(n_839),
.C(n_840),
.Y(n_5976)
);

AOI211xp5_ASAP7_75t_L g5977 ( 
.A1(n_5976),
.A2(n_845),
.B(n_843),
.C(n_844),
.Y(n_5977)
);


endmodule