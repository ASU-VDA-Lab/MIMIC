module fake_ibex_189_n_377 (n_85, n_84, n_64, n_3, n_73, n_65, n_95, n_55, n_63, n_98, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_97, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_96, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_377);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_95;
input n_55;
input n_63;
input n_98;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_97;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_96;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_377;

wire n_151;
wire n_171;
wire n_103;
wire n_204;
wire n_274;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_193;
wire n_108;
wire n_350;
wire n_165;
wire n_255;
wire n_175;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_239;
wire n_134;
wire n_371;
wire n_357;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_176;
wire n_216;
wire n_166;
wire n_163;
wire n_114;
wire n_236;
wire n_376;
wire n_189;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_187;
wire n_105;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_113;
wire n_117;
wire n_265;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_210;
wire n_348;
wire n_220;
wire n_287;
wire n_243;
wire n_228;
wire n_147;
wire n_251;
wire n_373;
wire n_244;
wire n_343;
wire n_310;
wire n_323;
wire n_143;
wire n_106;
wire n_224;
wire n_183;
wire n_333;
wire n_110;
wire n_306;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_109;
wire n_127;
wire n_121;
wire n_325;
wire n_301;
wire n_296;
wire n_120;
wire n_168;
wire n_155;
wire n_315;
wire n_122;
wire n_116;
wire n_370;
wire n_289;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_136;
wire n_261;
wire n_367;
wire n_221;
wire n_355;
wire n_102;
wire n_99;
wire n_269;
wire n_156;
wire n_126;
wire n_356;
wire n_104;
wire n_141;
wire n_222;
wire n_186;
wire n_349;
wire n_295;
wire n_331;
wire n_230;
wire n_185;
wire n_352;
wire n_290;
wire n_174;
wire n_157;
wire n_219;
wire n_246;
wire n_146;
wire n_207;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_139;
wire n_275;
wire n_129;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_347;
wire n_335;
wire n_263;
wire n_353;
wire n_359;
wire n_262;
wire n_299;
wire n_137;
wire n_338;
wire n_173;
wire n_363;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_257;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_365;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_329;
wire n_188;
wire n_200;
wire n_199;
wire n_308;
wire n_135;
wire n_283;
wire n_366;
wire n_111;
wire n_322;
wire n_227;
wire n_115;
wire n_248;
wire n_101;
wire n_190;
wire n_138;
wire n_214;
wire n_238;
wire n_332;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_225;
wire n_360;
wire n_272;
wire n_223;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_148;
wire n_342;
wire n_233;
wire n_118;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_178;
wire n_303;
wire n_362;
wire n_162;
wire n_240;
wire n_282;
wire n_266;
wire n_294;
wire n_112;
wire n_284;
wire n_172;
wire n_250;
wire n_313;
wire n_345;
wire n_119;
wire n_361;
wire n_319;
wire n_195;
wire n_212;
wire n_311;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_302;
wire n_344;
wire n_297;
wire n_252;
wire n_107;
wire n_149;
wire n_254;
wire n_213;
wire n_271;
wire n_241;
wire n_292;
wire n_364;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_160;
wire n_184;
wire n_232;
wire n_281;

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_43),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_8),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_41),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_40),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_0),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_12),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_54),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_21),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_18),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_17),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_34),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_44),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_13),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_46),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_50),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_24),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_22),
.Y(n_145)
);

INVxp33_ASAP7_75t_SL g146 ( 
.A(n_76),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_23),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_36),
.Y(n_154)
);

INVxp33_ASAP7_75t_SL g155 ( 
.A(n_25),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_52),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_32),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_19),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_5),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_15),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_0),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_27),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_73),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

INVxp33_ASAP7_75t_SL g171 ( 
.A(n_47),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_65),
.Y(n_173)
);

INVxp33_ASAP7_75t_SL g174 ( 
.A(n_63),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_45),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_26),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_95),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_4),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_56),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_10),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_30),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_98),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_71),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_33),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_62),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_103),
.A2(n_188),
.B1(n_111),
.B2(n_142),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_100),
.B(n_57),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_117),
.B(n_1),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_143),
.B(n_3),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_3),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g204 ( 
.A(n_110),
.B(n_4),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_112),
.A2(n_6),
.B1(n_7),
.B2(n_29),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_7),
.B1(n_58),
.B2(n_61),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_118),
.B(n_68),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_122),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_128),
.A2(n_72),
.B1(n_80),
.B2(n_87),
.Y(n_217)
);

AND3x1_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_146),
.A2(n_171),
.B1(n_155),
.B2(n_174),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_163),
.A2(n_175),
.B1(n_182),
.B2(n_190),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_115),
.A2(n_190),
.B1(n_139),
.B2(n_182),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_102),
.B(n_176),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_115),
.A2(n_139),
.B1(n_168),
.B2(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_102),
.A2(n_176),
.B1(n_124),
.B2(n_114),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_126),
.B(n_152),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_99),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_124),
.B(n_154),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_133),
.A2(n_157),
.B1(n_186),
.B2(n_134),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_137),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_R g240 ( 
.A1(n_140),
.A2(n_159),
.B1(n_184),
.B2(n_141),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_147),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_153),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_150),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_151),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_156),
.B(n_166),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_167),
.B1(n_181),
.B2(n_179),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_105),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_197),
.Y(n_253)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_200),
.A2(n_161),
.B(n_173),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_160),
.Y(n_257)
);

OAI221xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_169),
.B1(n_170),
.B2(n_109),
.C(n_149),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

OAI221xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_153),
.B1(n_185),
.B2(n_206),
.C(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_206),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_218),
.B1(n_226),
.B2(n_229),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_234),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

AO22x2_ASAP7_75t_L g270 ( 
.A1(n_217),
.A2(n_203),
.B1(n_216),
.B2(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_196),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

OAI221xp5_ASAP7_75t_L g277 ( 
.A1(n_237),
.A2(n_232),
.B1(n_242),
.B2(n_239),
.C(n_235),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_216),
.B(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_199),
.A2(n_217),
.B1(n_205),
.B2(n_222),
.Y(n_280)
);

AO22x2_ASAP7_75t_L g281 ( 
.A1(n_199),
.A2(n_225),
.B1(n_232),
.B2(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_201),
.Y(n_285)
);

AO22x2_ASAP7_75t_L g286 ( 
.A1(n_249),
.A2(n_221),
.B1(n_247),
.B2(n_207),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_211),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_212),
.B(n_223),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_250),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_215),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_194),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_210),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_215),
.B(n_244),
.Y(n_299)
);

AO22x2_ASAP7_75t_L g300 ( 
.A1(n_209),
.A2(n_226),
.B1(n_217),
.B2(n_229),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_194),
.Y(n_302)
);

AO22x2_ASAP7_75t_L g303 ( 
.A1(n_194),
.A2(n_226),
.B1(n_217),
.B2(n_229),
.Y(n_303)
);

AND2x4_ASAP7_75t_SL g304 ( 
.A(n_267),
.B(n_244),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_274),
.Y(n_306)
);

CKINVDCx8_ASAP7_75t_R g307 ( 
.A(n_267),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_257),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_253),
.B1(n_261),
.B2(n_254),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_268),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_268),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_255),
.B(n_277),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_280),
.Y(n_315)
);

BUFx2_ASAP7_75t_SL g316 ( 
.A(n_264),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_257),
.B(n_297),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_275),
.B(n_266),
.C(n_272),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_252),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_290),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_262),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_286),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_300),
.B1(n_270),
.B2(n_258),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_289),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_281),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_259),
.B(n_286),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_307),
.A2(n_287),
.B1(n_300),
.B2(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_305),
.B(n_302),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_318),
.A2(n_288),
.B(n_294),
.C(n_284),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_293),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_313),
.A2(n_301),
.B(n_265),
.C(n_295),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_289),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_299),
.B(n_269),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_308),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_270),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_310),
.A2(n_265),
.B(n_271),
.C(n_251),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_320),
.A2(n_256),
.B(n_322),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_317),
.Y(n_345)
);

BUFx8_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

O2A1O1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_320),
.B(n_323),
.C(n_327),
.Y(n_349)
);

AOI221xp5_ASAP7_75t_L g350 ( 
.A1(n_328),
.A2(n_324),
.B1(n_317),
.B2(n_323),
.C(n_304),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_309),
.Y(n_351)
);

AO32x2_ASAP7_75t_L g352 ( 
.A1(n_337),
.A2(n_343),
.A3(n_342),
.B1(n_340),
.B2(n_335),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_316),
.Y(n_353)
);

BUFx4f_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_319),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_347),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_329),
.B(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

AOI21x1_ASAP7_75t_L g360 ( 
.A1(n_352),
.A2(n_340),
.B(n_337),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_355),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_357),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_356),
.Y(n_364)
);

NAND4xp75_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_345),
.C(n_361),
.D(n_350),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_362),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_364),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_366),
.A2(n_362),
.B1(n_363),
.B2(n_353),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_367),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_369),
.B(n_367),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_370),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_368),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_365),
.C(n_335),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_346),
.B1(n_358),
.B2(n_340),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_374),
.A2(n_346),
.B1(n_358),
.B2(n_348),
.Y(n_375)
);

OAI222xp33_ASAP7_75t_L g376 ( 
.A1(n_375),
.A2(n_360),
.B1(n_351),
.B2(n_352),
.C1(n_314),
.C2(n_334),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_256),
.B1(n_321),
.B2(n_326),
.Y(n_377)
);


endmodule