module fake_jpeg_24749_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_21),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g16 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_4),
.C(n_13),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_7),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_23),
.B(n_8),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_28),
.C(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_21),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_38),
.B(n_39),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_29),
.B(n_17),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_19),
.C1(n_20),
.C2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);


endmodule