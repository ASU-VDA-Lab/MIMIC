module fake_jpeg_8789_n_33 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_33);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_1),
.A2(n_5),
.B1(n_0),
.B2(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_12),
.B(n_15),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_26),
.B(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_21),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_16),
.B1(n_6),
.B2(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_20),
.B1(n_2),
.B2(n_22),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_30),
.B1(n_25),
.B2(n_14),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_10),
.B(n_13),
.Y(n_33)
);


endmodule