module fake_jpeg_11792_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_11),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_52),
.Y(n_88)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_48),
.B(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_2),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_65),
.C(n_26),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_25),
.B(n_2),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_5),
.B(n_6),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_61),
.Y(n_100)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_23),
.B(n_10),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_12),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_14),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_67),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_14),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_27),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_70),
.B(n_79),
.Y(n_120)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_74),
.Y(n_118)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_22),
.B(n_33),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_22),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_80),
.Y(n_127)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_31),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_16),
.B(n_20),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_76),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_24),
.B(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_24),
.B(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_26),
.B(n_39),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_56),
.A2(n_20),
.B1(n_44),
.B2(n_42),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_89),
.A2(n_97),
.B1(n_103),
.B2(n_130),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_90),
.B(n_91),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_34),
.C(n_38),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_34),
.B1(n_38),
.B2(n_42),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_74),
.B1(n_80),
.B2(n_99),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_44),
.B1(n_32),
.B2(n_39),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_107),
.B1(n_111),
.B2(n_119),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_29),
.B1(n_32),
.B2(n_54),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_52),
.B1(n_61),
.B2(n_60),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_70),
.B1(n_53),
.B2(n_50),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_70),
.B1(n_53),
.B2(n_50),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_51),
.C(n_62),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_116),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_79),
.B(n_78),
.C(n_83),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_57),
.A2(n_68),
.B1(n_63),
.B2(n_45),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_47),
.B(n_73),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_58),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_59),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_80),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_71),
.B1(n_43),
.B2(n_41),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_87),
.B1(n_96),
.B2(n_117),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_56),
.B1(n_37),
.B2(n_61),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_133),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_142),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_139),
.B(n_148),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_104),
.B1(n_90),
.B2(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_104),
.B1(n_92),
.B2(n_126),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_91),
.A2(n_123),
.B1(n_130),
.B2(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_93),
.B1(n_88),
.B2(n_109),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_166),
.B1(n_157),
.B2(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_149),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_152),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_153),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_87),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_112),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_159),
.Y(n_175)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_137),
.B1(n_169),
.B2(n_134),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_106),
.B(n_112),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_109),
.A2(n_98),
.B1(n_105),
.B2(n_101),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_98),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_132),
.B1(n_162),
.B2(n_163),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_161),
.B(n_147),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_182),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_168),
.B1(n_135),
.B2(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_171),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_172),
.B(n_194),
.C(n_181),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_154),
.C(n_161),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_184),
.C(n_196),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_154),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_145),
.B1(n_133),
.B2(n_159),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_191),
.B1(n_194),
.B2(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_135),
.B1(n_138),
.B2(n_167),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_158),
.C(n_166),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_149),
.B1(n_145),
.B2(n_133),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_186),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_213),
.C(n_180),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_197),
.B(n_178),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_209),
.B(n_198),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_203),
.A2(n_212),
.B1(n_181),
.B2(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_182),
.B(n_196),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_216),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_195),
.B(n_193),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_189),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_171),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_185),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_187),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_177),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_225),
.B(n_201),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_210),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_175),
.B1(n_198),
.B2(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_227),
.C(n_214),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_193),
.B(n_183),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_231),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_223),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_236),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_202),
.C(n_200),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_237),
.C(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_202),
.C(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_239),
.A2(n_230),
.B1(n_201),
.B2(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_228),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_239),
.B1(n_232),
.B2(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_208),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_244),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_229),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_235),
.B(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_225),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_223),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_245),
.C(n_247),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_230),
.B(n_246),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_257),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_256),
.B(n_252),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_258),
.Y(n_261)
);


endmodule