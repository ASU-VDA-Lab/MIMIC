module fake_jpeg_995_n_677 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_677);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_677;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_17),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_58),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_59),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_60),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_61),
.Y(n_228)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_66),
.Y(n_200)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_11),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_69),
.A2(n_78),
.B(n_84),
.Y(n_197)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_72),
.Y(n_212)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_74),
.Y(n_227)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_11),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_11),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_98),
.Y(n_156)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_11),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_12),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_101),
.B(n_108),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_102),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_10),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

BUFx12f_ASAP7_75t_SL g114 ( 
.A(n_40),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_114),
.B(n_21),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_24),
.B(n_55),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_116),
.B(n_50),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_118),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_42),
.Y(n_119)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_50),
.B(n_10),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_120),
.B(n_13),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_35),
.Y(n_123)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_37),
.Y(n_129)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_54),
.Y(n_157)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_45),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_133),
.B(n_147),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_128),
.B1(n_127),
.B2(n_121),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_135),
.A2(n_148),
.B1(n_160),
.B2(n_166),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_45),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_84),
.A2(n_54),
.B1(n_49),
.B2(n_53),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_25),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_151),
.B(n_199),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_157),
.B(n_230),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_53),
.B1(n_54),
.B2(n_28),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_53),
.B1(n_41),
.B2(n_28),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_101),
.A2(n_30),
.B1(n_22),
.B2(n_41),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_174),
.A2(n_179),
.B1(n_205),
.B2(n_210),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_73),
.B(n_52),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_178),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_85),
.A2(n_22),
.B1(n_30),
.B2(n_52),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_185),
.B(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_190),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_59),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_193),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_194),
.A2(n_221),
.B(n_191),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_92),
.B(n_51),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_202),
.Y(n_290)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_60),
.Y(n_203)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_203),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_106),
.B(n_51),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_204),
.B(n_206),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_87),
.A2(n_55),
.B1(n_21),
.B2(n_39),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_61),
.B(n_15),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_119),
.B(n_15),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_217),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_100),
.A2(n_21),
.B1(n_39),
.B2(n_56),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_63),
.B(n_14),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_64),
.B(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_65),
.Y(n_218)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_218),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_58),
.B(n_13),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_222),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_89),
.B(n_13),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_71),
.Y(n_225)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_102),
.Y(n_226)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_103),
.A2(n_21),
.B1(n_37),
.B2(n_1),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_229),
.A2(n_19),
.B1(n_175),
.B2(n_169),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_115),
.B(n_56),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_230),
.B(n_176),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_105),
.A2(n_56),
.B1(n_42),
.B2(n_3),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_107),
.B1(n_112),
.B2(n_42),
.Y(n_243)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_234),
.Y(n_330)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

INVx4_ASAP7_75t_SL g382 ( 
.A(n_235),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_236),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_238),
.B(n_247),
.Y(n_334)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_240),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_178),
.B(n_117),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_241),
.Y(n_361)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_242),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_243),
.A2(n_294),
.B1(n_298),
.B2(n_308),
.Y(n_367)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_244),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_134),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_245),
.Y(n_369)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_174),
.A2(n_140),
.B(n_196),
.C(n_148),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g355 ( 
.A1(n_246),
.A2(n_296),
.B1(n_251),
.B2(n_247),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_155),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_156),
.A2(n_9),
.B1(n_2),
.B2(n_5),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_248),
.A2(n_252),
.B1(n_257),
.B2(n_283),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_250),
.B(n_258),
.Y(n_327)
);

BUFx8_ASAP7_75t_L g251 ( 
.A(n_140),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_157),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_254),
.Y(n_323)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_146),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_259),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_138),
.B(n_1),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_260),
.Y(n_376)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_261),
.Y(n_359)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_263),
.Y(n_373)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

AOI32xp33_ASAP7_75t_L g265 ( 
.A1(n_197),
.A2(n_7),
.A3(n_9),
.B1(n_16),
.B2(n_17),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_265),
.B(n_291),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_141),
.B(n_7),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_267),
.B(n_278),
.C(n_309),
.Y(n_339)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_143),
.Y(n_269)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_269),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_135),
.A2(n_7),
.B1(n_17),
.B2(n_18),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_270),
.A2(n_276),
.B1(n_282),
.B2(n_289),
.Y(n_354)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_163),
.Y(n_273)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_273),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_179),
.A2(n_18),
.B1(n_19),
.B2(n_229),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_277),
.B(n_284),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_145),
.B(n_18),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_139),
.Y(n_280)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_280),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_146),
.A2(n_19),
.B1(n_227),
.B2(n_132),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_182),
.Y(n_284)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_143),
.Y(n_285)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_144),
.Y(n_286)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_286),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_197),
.A2(n_136),
.B(n_181),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_315),
.Y(n_321)
);

INVx5_ASAP7_75t_SL g288 ( 
.A(n_182),
.Y(n_288)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_171),
.A2(n_19),
.B1(n_186),
.B2(n_168),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_215),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_293),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_212),
.A2(n_167),
.B1(n_172),
.B2(n_214),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_295),
.B(n_300),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_219),
.A2(n_223),
.B1(n_187),
.B2(n_198),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_299),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_212),
.A2(n_169),
.B1(n_219),
.B2(n_165),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_175),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_143),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_301),
.B(n_307),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_158),
.B(n_164),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_302),
.B(n_253),
.Y(n_341)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_176),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_305),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_142),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_306),
.B(n_312),
.Y(n_380)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_142),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_173),
.A2(n_213),
.B1(n_184),
.B2(n_161),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_180),
.B(n_183),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_137),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_215),
.B(n_228),
.C(n_180),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_228),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_316),
.Y(n_338)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_137),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_317),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_150),
.B(n_153),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_150),
.B(n_153),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_241),
.Y(n_347)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_154),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_320),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_287),
.A2(n_154),
.B1(n_246),
.B2(n_243),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_326),
.A2(n_349),
.B1(n_362),
.B2(n_289),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_262),
.B(n_311),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_365),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_260),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_335),
.B(n_346),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_341),
.B(n_372),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_260),
.B(n_267),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_235),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_249),
.A2(n_241),
.B1(n_313),
.B2(n_271),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_267),
.B(n_278),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_357),
.Y(n_391)
);

OAI21xp33_ASAP7_75t_SL g405 ( 
.A1(n_355),
.A2(n_301),
.B(n_288),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_278),
.B(n_281),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_238),
.A2(n_276),
.B1(n_308),
.B2(n_275),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_239),
.B(n_238),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_379),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_272),
.B(n_295),
.Y(n_365)
);

MAJx2_ASAP7_75t_L g366 ( 
.A(n_274),
.B(n_290),
.C(n_251),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_371),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_266),
.B(n_314),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_305),
.B(n_268),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_233),
.B(n_292),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_376),
.B(n_310),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_385),
.B(n_410),
.Y(n_449)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_382),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_364),
.B(n_309),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_388),
.B(n_425),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_327),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_399),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_390),
.B(n_393),
.Y(n_464)
);

NAND2x1p5_ASAP7_75t_L g393 ( 
.A(n_321),
.B(n_303),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_349),
.A2(n_309),
.B1(n_319),
.B2(n_318),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_394),
.A2(n_395),
.B1(n_405),
.B2(n_416),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_354),
.A2(n_319),
.B1(n_318),
.B2(n_270),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_326),
.A2(n_317),
.B1(n_316),
.B2(n_304),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_396),
.A2(n_403),
.B1(n_415),
.B2(n_423),
.Y(n_459)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_321),
.A2(n_250),
.B(n_258),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_398),
.A2(n_407),
.B(n_343),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_379),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_400),
.B(n_413),
.Y(n_453)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_381),
.Y(n_401)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_401),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_362),
.A2(n_315),
.B1(n_320),
.B2(n_306),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_261),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_404),
.Y(n_470)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_381),
.Y(n_406)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_369),
.A2(n_285),
.B1(n_236),
.B2(n_279),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_264),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_357),
.B(n_244),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_412),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_263),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_332),
.B(n_240),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_421),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_354),
.A2(n_237),
.B1(n_293),
.B2(n_307),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_335),
.A2(n_242),
.B1(n_269),
.B2(n_361),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_417),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_325),
.B(n_346),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_422),
.Y(n_462)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_419),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_336),
.A2(n_375),
.B1(n_355),
.B2(n_325),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_420),
.A2(n_331),
.B1(n_348),
.B2(n_373),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_380),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_330),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_365),
.A2(n_347),
.B1(n_367),
.B2(n_339),
.Y(n_423)
);

O2A1O1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_355),
.A2(n_369),
.B(n_366),
.C(n_370),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_424),
.A2(n_432),
.B(n_398),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_334),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_355),
.A2(n_324),
.B1(n_338),
.B2(n_360),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_426),
.A2(n_430),
.B1(n_329),
.B2(n_359),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_352),
.B(n_339),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_427),
.B(n_431),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_334),
.B(n_358),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_340),
.C(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_323),
.Y(n_429)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_368),
.A2(n_328),
.B1(n_337),
.B2(n_359),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_330),
.B(n_337),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_333),
.A2(n_356),
.B(n_370),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_456),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_441),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_377),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_443),
.B(n_454),
.C(n_455),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_428),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_409),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_447),
.B(n_448),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_431),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_378),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_452),
.B(n_461),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_374),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_383),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_410),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_402),
.B(n_351),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_458),
.B(n_466),
.C(n_468),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_460),
.Y(n_477)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_401),
.Y(n_463)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_463),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_422),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_467),
.Y(n_478)
);

MAJx2_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_351),
.C(n_344),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_404),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_423),
.B(n_344),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_420),
.A2(n_373),
.B1(n_353),
.B2(n_348),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_471),
.A2(n_424),
.B(n_432),
.Y(n_479)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_417),
.Y(n_472)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_390),
.A2(n_342),
.B1(n_322),
.B2(n_343),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_474),
.A2(n_387),
.B1(n_386),
.B2(n_419),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_404),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_425),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_446),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_480),
.B(n_482),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_439),
.Y(n_481)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_481),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_446),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_489),
.C(n_505),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_427),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_445),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_436),
.A2(n_395),
.B1(n_399),
.B2(n_424),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_485),
.A2(n_503),
.B1(n_459),
.B2(n_461),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_L g487 ( 
.A1(n_444),
.A2(n_393),
.B(n_384),
.Y(n_487)
);

BUFx5_ASAP7_75t_L g551 ( 
.A(n_487),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_418),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_490),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_434),
.A2(n_396),
.B1(n_415),
.B2(n_403),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_493),
.A2(n_499),
.B1(n_504),
.B2(n_509),
.Y(n_521)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_495),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_470),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_434),
.A2(n_392),
.B1(n_412),
.B2(n_384),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_438),
.A2(n_393),
.B(n_394),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_500),
.A2(n_514),
.B(n_495),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_465),
.B(n_473),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_501),
.B(n_507),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_464),
.A2(n_392),
.B1(n_400),
.B2(n_391),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_454),
.B(n_400),
.C(n_391),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_468),
.B(n_458),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_506),
.B(n_508),
.C(n_510),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_457),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_453),
.B(n_385),
.C(n_411),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_464),
.A2(n_388),
.B1(n_416),
.B2(n_429),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_453),
.B(n_397),
.C(n_345),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_457),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_511),
.B(n_513),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_466),
.B(n_345),
.C(n_353),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_512),
.B(n_440),
.C(n_450),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_462),
.B(n_449),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_464),
.A2(n_460),
.B(n_456),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_462),
.B(n_342),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g533 ( 
.A(n_515),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_516),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_492),
.Y(n_517)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_517),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_449),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_518),
.B(n_529),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_527),
.B1(n_534),
.B2(n_540),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_522),
.B(n_510),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_478),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_546),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_509),
.A2(n_459),
.B1(n_474),
.B2(n_451),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_528),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_451),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_500),
.A2(n_475),
.B1(n_467),
.B2(n_435),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_530),
.A2(n_535),
.B1(n_541),
.B2(n_549),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_506),
.B(n_502),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_531),
.B(n_508),
.Y(n_557)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_492),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_514),
.A2(n_469),
.B1(n_433),
.B2(n_435),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_486),
.B(n_470),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_537),
.B(n_512),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_477),
.A2(n_433),
.B1(n_463),
.B2(n_437),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_539),
.A2(n_543),
.B(n_498),
.Y(n_569)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_492),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_477),
.A2(n_437),
.B1(n_440),
.B2(n_450),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_547),
.C(n_548),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_479),
.A2(n_472),
.B1(n_442),
.B2(n_322),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_544),
.A2(n_476),
.B1(n_497),
.B2(n_539),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_480),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_486),
.B(n_483),
.C(n_489),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_502),
.B(n_484),
.C(n_505),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_496),
.A2(n_499),
.B1(n_494),
.B2(n_476),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_482),
.B(n_511),
.Y(n_552)
);

CKINVDCx14_ASAP7_75t_R g567 ( 
.A(n_552),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_532),
.Y(n_553)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_553),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_557),
.B(n_570),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_550),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_561),
.B(n_565),
.Y(n_604)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_552),
.Y(n_564)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_564),
.Y(n_595)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_550),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_526),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_566),
.B(n_568),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_528),
.B(n_507),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_569),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_571),
.B(n_573),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_537),
.B(n_504),
.C(n_498),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_576),
.C(n_579),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_SL g573 ( 
.A(n_531),
.B(n_493),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_521),
.A2(n_527),
.B1(n_525),
.B2(n_536),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_574),
.A2(n_578),
.B1(n_580),
.B2(n_581),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_525),
.B(n_488),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_575),
.B(n_577),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_538),
.B(n_547),
.C(n_524),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_545),
.B(n_488),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_545),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_538),
.B(n_497),
.C(n_503),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_519),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_519),
.B(n_523),
.C(n_551),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_582),
.B(n_566),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_556),
.A2(n_521),
.B1(n_536),
.B2(n_543),
.Y(n_587)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_580),
.A2(n_578),
.B1(n_555),
.B2(n_567),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_590),
.A2(n_597),
.B1(n_605),
.B2(n_604),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_558),
.B(n_542),
.C(n_524),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_591),
.B(n_593),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_556),
.A2(n_517),
.B1(n_544),
.B2(n_533),
.Y(n_592)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_592),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_558),
.B(n_548),
.C(n_522),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_564),
.Y(n_594)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_594),
.Y(n_613)
);

FAx1_ASAP7_75t_SL g596 ( 
.A(n_573),
.B(n_530),
.CI(n_535),
.CON(n_596),
.SN(n_596)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_596),
.B(n_600),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_559),
.A2(n_577),
.B1(n_561),
.B2(n_565),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_563),
.A2(n_520),
.B1(n_523),
.B2(n_549),
.Y(n_598)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_598),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_579),
.B(n_541),
.C(n_532),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_602),
.C(n_603),
.Y(n_615)
);

FAx1_ASAP7_75t_SL g600 ( 
.A(n_574),
.B(n_572),
.CI(n_551),
.CON(n_600),
.SN(n_600)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_576),
.B(n_570),
.C(n_571),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_557),
.B(n_554),
.C(n_559),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_569),
.B(n_563),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_605),
.B(n_562),
.Y(n_609)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_606),
.Y(n_608)
);

MAJx2_ASAP7_75t_L g630 ( 
.A(n_609),
.B(n_626),
.C(n_601),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_599),
.B(n_560),
.Y(n_610)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_610),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_589),
.B(n_568),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_583),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_591),
.B(n_554),
.C(n_560),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_617),
.B(n_620),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_585),
.B(n_575),
.Y(n_619)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_619),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_584),
.B(n_603),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_607),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_621),
.A2(n_627),
.B(n_628),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_607),
.A2(n_595),
.B1(n_586),
.B2(n_604),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_622),
.A2(n_625),
.B1(n_621),
.B2(n_616),
.Y(n_633)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_594),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_623),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_SL g626 ( 
.A(n_601),
.B(n_588),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_SL g627 ( 
.A1(n_600),
.A2(n_596),
.B(n_587),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_592),
.A2(n_598),
.B(n_585),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_628),
.A2(n_627),
.B(n_618),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_624),
.B(n_602),
.C(n_584),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_629),
.B(n_635),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_630),
.B(n_631),
.Y(n_647)
);

NOR2x1p5_ASAP7_75t_L g632 ( 
.A(n_611),
.B(n_596),
.Y(n_632)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_632),
.Y(n_646)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_633),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_615),
.B(n_593),
.C(n_588),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_637),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_615),
.B(n_600),
.C(n_620),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_638),
.B(n_639),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_617),
.B(n_609),
.C(n_611),
.Y(n_639)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_640),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_626),
.B(n_622),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_642),
.B(n_645),
.Y(n_652)
);

NOR2x1_ASAP7_75t_L g643 ( 
.A(n_619),
.B(n_618),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_643),
.A2(n_614),
.B(n_612),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_612),
.A2(n_614),
.B1(n_608),
.B2(n_613),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_629),
.B(n_636),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_648),
.B(n_649),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_634),
.B(n_613),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_650),
.B(n_655),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_639),
.B(n_641),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_654),
.B(n_643),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_658),
.B(n_659),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_SL g659 ( 
.A1(n_657),
.A2(n_637),
.B(n_632),
.Y(n_659)
);

BUFx24_ASAP7_75t_SL g660 ( 
.A(n_653),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_660),
.B(n_665),
.Y(n_666)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_652),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_661),
.A2(n_651),
.B1(n_631),
.B2(n_646),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_SL g663 ( 
.A1(n_656),
.A2(n_644),
.B1(n_638),
.B2(n_642),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_663),
.B(n_647),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_656),
.B(n_633),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_662),
.B(n_652),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_668),
.B(n_669),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_670),
.B(n_668),
.Y(n_672)
);

NOR3xp33_ASAP7_75t_L g673 ( 
.A(n_672),
.B(n_664),
.C(n_667),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_673),
.A2(n_671),
.B(n_666),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_674),
.A2(n_649),
.B(n_645),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_675),
.A2(n_632),
.B(n_647),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_676),
.A2(n_635),
.B(n_630),
.Y(n_677)
);


endmodule