module fake_jpeg_22582_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_4),
.B(n_13),
.Y(n_19)
);

CKINVDCx11_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_44),
.Y(n_58)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_45),
.Y(n_70)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_1),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_1),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_55),
.B1(n_74),
.B2(n_33),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_26),
.B1(n_37),
.B2(n_36),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_57),
.B(n_61),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_85),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_24),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_36),
.B1(n_37),
.B2(n_17),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_18),
.B1(n_31),
.B2(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_18),
.B1(n_31),
.B2(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_67),
.Y(n_96)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_21),
.B1(n_48),
.B2(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_82),
.B1(n_27),
.B2(n_32),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_30),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_22),
.B1(n_23),
.B2(n_20),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_77),
.Y(n_105)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_27),
.B1(n_32),
.B2(n_28),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_87),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_92),
.A2(n_67),
.B(n_56),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_54),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_88),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_50),
.B1(n_56),
.B2(n_83),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_102),
.Y(n_131)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_109),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_52),
.A2(n_33),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_70),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_55),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_8),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_30),
.C(n_24),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_85),
.C(n_87),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_50),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_52),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_5),
.C(n_6),
.Y(n_142)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_16),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_53),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_135),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_126),
.Y(n_159)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_128),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_90),
.B1(n_95),
.B2(n_102),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_103),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_64),
.C(n_65),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_86),
.C(n_59),
.Y(n_177)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_62),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_24),
.B(n_59),
.C(n_66),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_143),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_117),
.B1(n_100),
.B2(n_112),
.Y(n_156)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_84),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_24),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_149),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_24),
.Y(n_174)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_76),
.B1(n_86),
.B2(n_24),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_98),
.B1(n_91),
.B2(n_89),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_101),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_151),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_99),
.B1(n_108),
.B2(n_90),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_94),
.B(n_113),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_170),
.B(n_146),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_178),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_171),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_172),
.B1(n_127),
.B2(n_128),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_179),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_130),
.A2(n_100),
.B1(n_112),
.B2(n_118),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_180),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_110),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_182),
.C(n_135),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_108),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_95),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_184),
.B(n_191),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_190),
.C(n_178),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_199),
.B(n_200),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_174),
.C(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_196),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_155),
.A2(n_130),
.B1(n_136),
.B2(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2x1_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_149),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_141),
.B(n_133),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_164),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_203),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_132),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_158),
.Y(n_226)
);

AOI22x1_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_140),
.B1(n_134),
.B2(n_123),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_90),
.B1(n_145),
.B2(n_124),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_160),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_212),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_217),
.A2(n_223),
.B1(n_124),
.B2(n_196),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_199),
.B(n_159),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_222),
.C(n_227),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_195),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_192),
.B(n_191),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_226),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_199),
.B(n_198),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_226),
.B(n_220),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_201),
.B1(n_194),
.B2(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_193),
.B1(n_189),
.B2(n_201),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_237),
.B1(n_238),
.B2(n_208),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_190),
.C(n_187),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_242),
.C(n_209),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_240),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_189),
.B1(n_205),
.B2(n_171),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_205),
.B1(n_172),
.B2(n_184),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_238),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_195),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_156),
.B1(n_217),
.B2(n_213),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_176),
.C(n_204),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_224),
.B1(n_218),
.B2(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_181),
.B1(n_233),
.B2(n_148),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_230),
.C(n_242),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_240),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_213),
.B(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_223),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_99),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_181),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_263),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_230),
.C(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_252),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_256),
.B(n_251),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_271),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_248),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_245),
.B(n_247),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_261),
.B(n_263),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_258),
.C(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_260),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_8),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_282),
.B1(n_14),
.B2(n_10),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_283),
.C(n_276),
.Y(n_285)
);

OAI321xp33_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_264),
.A3(n_262),
.B1(n_16),
.B2(n_15),
.C(n_143),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.C(n_9),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_287),
.A2(n_284),
.B(n_10),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_288),
.Y(n_290)
);


endmodule