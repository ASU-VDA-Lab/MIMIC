module fake_jpeg_1269_n_165 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_49),
.B1(n_19),
.B2(n_21),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_23),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_50),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_51),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_15),
.A2(n_27),
.B1(n_17),
.B2(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_25),
.B(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_15),
.Y(n_65)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_46),
.Y(n_75)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_78),
.B1(n_81),
.B2(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_7),
.B1(n_35),
.B2(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_32),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_9),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_10),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_88),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_37),
.A2(n_34),
.B1(n_43),
.B2(n_54),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_40),
.A2(n_10),
.B(n_6),
.C(n_7),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_5),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_96),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_7),
.B1(n_77),
.B2(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_103),
.Y(n_122)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_93),
.Y(n_111)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_64),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_86),
.A3(n_58),
.B1(n_70),
.B2(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_77),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_79),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_70),
.B1(n_89),
.B2(n_73),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_87),
.B(n_63),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_87),
.A3(n_73),
.B1(n_61),
.B2(n_71),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_79),
.B(n_83),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_60),
.B(n_80),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_119),
.B(n_116),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_83),
.B(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_91),
.B1(n_103),
.B2(n_108),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_122),
.B1(n_118),
.B2(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_111),
.C(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_107),
.C(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.C(n_132),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_109),
.C(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_133),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_142),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_132),
.C(n_131),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_126),
.C(n_111),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_91),
.B1(n_121),
.B2(n_90),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_102),
.B1(n_105),
.B2(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_145),
.C(n_146),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_106),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_106),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_148),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_99),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_149),
.B(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_152),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_137),
.A3(n_143),
.B1(n_139),
.B2(n_97),
.C1(n_93),
.C2(n_114),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_154),
.B(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_144),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_146),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_159),
.B(n_139),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_162),
.C(n_99),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_114),
.B(n_94),
.Y(n_165)
);


endmodule