module fake_jpeg_30670_n_527 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_68),
.Y(n_112)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_32),
.B(n_7),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_76),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_8),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_22),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_81),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_32),
.B(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_99),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_33),
.B(n_8),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_33),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_104),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_37),
.B(n_8),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_22),
.B(n_50),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_111),
.B(n_144),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_52),
.B1(n_41),
.B2(n_36),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_113),
.A2(n_116),
.B1(n_125),
.B2(n_28),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_70),
.A2(n_52),
.B1(n_31),
.B2(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_55),
.B(n_44),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_120),
.B(n_129),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_67),
.A2(n_39),
.B1(n_38),
.B2(n_47),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_65),
.A2(n_34),
.B(n_50),
.C(n_24),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_52),
.B1(n_36),
.B2(n_31),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_134),
.A2(n_163),
.B1(n_45),
.B2(n_61),
.Y(n_214)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_39),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_137),
.B(n_66),
.Y(n_193)
);

BUFx4f_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_138),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_78),
.A2(n_51),
.B1(n_42),
.B2(n_24),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_43),
.B1(n_28),
.B2(n_74),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_73),
.A2(n_31),
.B1(n_51),
.B2(n_43),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_96),
.B(n_47),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_44),
.Y(n_170)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_174),
.Y(n_221)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_171),
.Y(n_258)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_71),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_37),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_179),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_178),
.B(n_181),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_113),
.A2(n_58),
.B1(n_80),
.B2(n_88),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_183),
.B1(n_214),
.B2(n_217),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_102),
.B1(n_103),
.B2(n_53),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_156),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_193),
.Y(n_225)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_195),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_196),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_152),
.A2(n_54),
.B1(n_77),
.B2(n_100),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_198),
.B1(n_203),
.B2(n_209),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_149),
.A2(n_150),
.B1(n_133),
.B2(n_145),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_200),
.Y(n_239)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_131),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_202),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_205),
.Y(n_249)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

BUFx16f_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_105),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_218),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_215),
.Y(n_235)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_149),
.A2(n_56),
.B1(n_59),
.B2(n_90),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_213),
.B(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_112),
.A2(n_98),
.B1(n_95),
.B2(n_91),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_147),
.B(n_42),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_159),
.B1(n_153),
.B2(n_165),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_219),
.A2(n_245),
.B1(n_260),
.B2(n_134),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_112),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_227),
.B(n_216),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_148),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_136),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_248),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_179),
.B(n_136),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_188),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_155),
.B1(n_161),
.B2(n_154),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_197),
.A2(n_143),
.B1(n_57),
.B2(n_82),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_173),
.B1(n_189),
.B2(n_184),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_171),
.B(n_83),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_149),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_257),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_150),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_183),
.A2(n_150),
.B1(n_163),
.B2(n_141),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_212),
.B1(n_198),
.B2(n_204),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_267),
.B1(n_273),
.B2(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_272),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_229),
.A2(n_194),
.B1(n_172),
.B2(n_180),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_265),
.A2(n_250),
.B(n_224),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_242),
.A2(n_160),
.B1(n_168),
.B2(n_190),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_268),
.A2(n_292),
.B(n_232),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_259),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_231),
.A2(n_187),
.B1(n_203),
.B2(n_176),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_296),
.B1(n_224),
.B2(n_252),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_245),
.A2(n_242),
.B1(n_239),
.B2(n_222),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_127),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_259),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_279),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_244),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_239),
.B1(n_222),
.B2(n_221),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_280),
.A2(n_283),
.B1(n_284),
.B2(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_221),
.A2(n_162),
.B1(n_139),
.B2(n_84),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_235),
.A2(n_209),
.B1(n_127),
.B2(n_45),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_230),
.B(n_46),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_294),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_227),
.B(n_127),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_244),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_246),
.A2(n_189),
.B1(n_209),
.B2(n_46),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_223),
.B(n_29),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_258),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_230),
.A2(n_45),
.B1(n_46),
.B2(n_29),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_261),
.A2(n_254),
.B1(n_225),
.B2(n_243),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_306),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_225),
.B1(n_232),
.B2(n_228),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_300),
.A2(n_315),
.B1(n_326),
.B2(n_263),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_305),
.A2(n_310),
.B(n_285),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_275),
.A2(n_254),
.B1(n_226),
.B2(n_223),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_287),
.C(n_266),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_307),
.B(n_324),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_234),
.B(n_244),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_312),
.A2(n_317),
.B1(n_319),
.B2(n_292),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_273),
.A2(n_247),
.B1(n_228),
.B2(n_226),
.Y(n_317)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_280),
.A2(n_247),
.B1(n_226),
.B2(n_255),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_236),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_277),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_262),
.A2(n_290),
.B1(n_281),
.B2(n_268),
.Y(n_326)
);

AO22x1_ASAP7_75t_SL g328 ( 
.A1(n_267),
.A2(n_251),
.B1(n_258),
.B2(n_252),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_286),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_284),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_279),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_347),
.Y(n_371)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_289),
.Y(n_335)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_291),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_297),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_339),
.A2(n_313),
.B(n_325),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_314),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_340),
.B(n_346),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_327),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_342),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_271),
.B(n_274),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_343),
.A2(n_358),
.B(n_325),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_299),
.A2(n_264),
.B(n_282),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_344),
.A2(n_345),
.B(n_29),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_301),
.A2(n_306),
.B(n_310),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_314),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_302),
.A2(n_288),
.B1(n_283),
.B2(n_270),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_348),
.A2(n_319),
.B1(n_312),
.B2(n_317),
.Y(n_364)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_350),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_326),
.A2(n_269),
.B1(n_278),
.B2(n_286),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_351),
.A2(n_355),
.B1(n_362),
.B2(n_329),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_302),
.A2(n_255),
.B1(n_251),
.B2(n_295),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_357),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_318),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_353),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_237),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_354),
.B(n_359),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_320),
.A2(n_251),
.B1(n_294),
.B2(n_236),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_324),
.Y(n_366)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_304),
.A2(n_236),
.B(n_237),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_316),
.B(n_12),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_308),
.B(n_12),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_360),
.B(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_304),
.A2(n_237),
.B1(n_1),
.B2(n_2),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_363),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_364),
.A2(n_374),
.B1(n_347),
.B2(n_331),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_323),
.C(n_298),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_366),
.C(n_372),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_384),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_307),
.C(n_297),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_356),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_375),
.C(n_386),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_358),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_383),
.B(n_395),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_328),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_343),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_380),
.B(n_360),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_311),
.B(n_303),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_341),
.A2(n_329),
.B(n_328),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_311),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_342),
.B(n_46),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_387),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_336),
.B(n_46),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_390),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_335),
.C(n_345),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_359),
.B(n_6),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_394),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_29),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_393),
.A2(n_333),
.B1(n_353),
.B2(n_341),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_397),
.A2(n_409),
.B1(n_416),
.B2(n_410),
.Y(n_444)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_385),
.Y(n_400)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_401),
.Y(n_434)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_402),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_406),
.Y(n_426)
);

BUFx12_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_408),
.B(n_410),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_371),
.A2(n_337),
.B1(n_351),
.B2(n_343),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_337),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_422),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_393),
.A2(n_352),
.B1(n_340),
.B2(n_346),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_414),
.A2(n_415),
.B1(n_418),
.B2(n_423),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_371),
.A2(n_355),
.B1(n_349),
.B2(n_361),
.Y(n_416)
);

BUFx12f_ASAP7_75t_SL g417 ( 
.A(n_390),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_419),
.B(n_379),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_374),
.A2(n_357),
.B1(n_334),
.B2(n_363),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_358),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_377),
.B(n_362),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_403),
.B(n_375),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_436),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_365),
.C(n_366),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_430),
.C(n_432),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_372),
.C(n_373),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_386),
.C(n_383),
.Y(n_432)
);

XOR2x2_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_395),
.Y(n_436)
);

XOR2x2_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_378),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_437),
.B(n_440),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_411),
.A2(n_388),
.B(n_391),
.Y(n_438)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_438),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_394),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_444),
.Y(n_457)
);

XOR2x2_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_379),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_391),
.C(n_389),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_443),
.C(n_445),
.Y(n_458)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_442),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_370),
.C(n_381),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_398),
.B(n_400),
.C(n_401),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_424),
.B(n_408),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_450),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_432),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_452),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_397),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_433),
.A2(n_420),
.B1(n_409),
.B2(n_406),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_455),
.A2(n_422),
.B1(n_405),
.B2(n_421),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_415),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_425),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_418),
.C(n_416),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_460),
.C(n_439),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_404),
.C(n_419),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_434),
.B(n_423),
.Y(n_461)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_462),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_443),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_464),
.A2(n_437),
.B1(n_436),
.B2(n_440),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_370),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_465),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_431),
.B(n_426),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_476),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_460),
.A2(n_444),
.B1(n_464),
.B2(n_449),
.Y(n_470)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_458),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_457),
.A2(n_425),
.B1(n_446),
.B2(n_379),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_474),
.A2(n_463),
.B1(n_13),
.B2(n_14),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_478),
.B(n_480),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_405),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_471),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_459),
.A2(n_405),
.B1(n_11),
.B2(n_13),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_456),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_481),
.B(n_482),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_453),
.A2(n_6),
.B(n_16),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_447),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_487),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_493),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_458),
.C(n_447),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_489),
.B(n_495),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_451),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_494),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_463),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_4),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_29),
.Y(n_496)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_496),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_470),
.B(n_4),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_497),
.B(n_474),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_490),
.A2(n_477),
.B1(n_475),
.B2(n_468),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_498),
.B(n_497),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_505),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_484),
.A2(n_467),
.B(n_469),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_501),
.A2(n_507),
.B(n_488),
.Y(n_509)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_491),
.A2(n_4),
.B(n_15),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_485),
.A2(n_5),
.B1(n_16),
.B2(n_2),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_493),
.C(n_5),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_489),
.A2(n_5),
.B(n_1),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_511),
.Y(n_518)
);

AOI21xp33_ASAP7_75t_L g510 ( 
.A1(n_502),
.A2(n_486),
.B(n_495),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_515),
.B(n_503),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_500),
.B(n_508),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_514),
.Y(n_519)
);

AOI21x1_ASAP7_75t_SL g515 ( 
.A1(n_505),
.A2(n_5),
.B(n_2),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_516),
.B(n_517),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_498),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_505),
.B(n_499),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_519),
.C(n_515),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_521),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_504),
.B(n_2),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_0),
.B(n_3),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_0),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_0),
.B(n_3),
.Y(n_527)
);


endmodule