module fake_jpeg_16265_n_59 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_43;
wire n_29;
wire n_37;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

AO22x1_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_5),
.B1(n_10),
.B2(n_0),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_2),
.C(n_29),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_27),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_45),
.C(n_44),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_38),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_48),
.B(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_46),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_50),
.B(n_24),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_21),
.Y(n_59)
);


endmodule