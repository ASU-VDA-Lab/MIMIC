module fake_jpeg_30583_n_553 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_553);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_553;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_10),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_4),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_55),
.B(n_56),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_60),
.B(n_61),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_62),
.B(n_63),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_67),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_71),
.B(n_77),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_39),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_25),
.B(n_15),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_81),
.B(n_86),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_87),
.B(n_100),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_12),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_91),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_29),
.B(n_12),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

CKINVDCx10_ASAP7_75t_R g99 ( 
.A(n_44),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_41),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_107),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_20),
.B1(n_23),
.B2(n_42),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_109),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_138),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_137),
.B(n_146),
.Y(n_211)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_78),
.B(n_48),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_148),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_84),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_144),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_65),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_86),
.B(n_48),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_95),
.A2(n_32),
.B1(n_29),
.B2(n_42),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_96),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_85),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_150),
.B(n_93),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_93),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_166),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_64),
.A2(n_42),
.B1(n_32),
.B2(n_27),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_35),
.B1(n_37),
.B2(n_43),
.Y(n_193)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_122),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_174),
.Y(n_278)
);

OAI22x1_ASAP7_75t_L g242 ( 
.A1(n_175),
.A2(n_120),
.B1(n_75),
.B2(n_58),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_176),
.B(n_201),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_178),
.A2(n_70),
.B1(n_134),
.B2(n_117),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_45),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_187),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_53),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_181),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_53),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_183),
.Y(n_269)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_27),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_45),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_188),
.B(n_192),
.Y(n_277)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_154),
.A2(n_33),
.B(n_28),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_43),
.B(n_37),
.C(n_30),
.Y(n_241)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_24),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_193),
.A2(n_215),
.B1(n_178),
.B2(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_96),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_200),
.Y(n_239)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_125),
.A2(n_35),
.B1(n_20),
.B2(n_106),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_202),
.A2(n_219),
.B1(n_158),
.B2(n_120),
.Y(n_233)
);

BUFx4f_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_203),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_125),
.B(n_28),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_214),
.Y(n_243)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_130),
.B(n_35),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_63),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_36),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_115),
.A2(n_105),
.B1(n_103),
.B2(n_101),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_33),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_217),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_121),
.B(n_36),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_221),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_115),
.A2(n_54),
.B1(n_75),
.B2(n_23),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_142),
.B(n_63),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_225),
.B(n_165),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_124),
.B(n_30),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_227),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_180),
.A2(n_121),
.B1(n_119),
.B2(n_126),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_235),
.B(n_241),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_242),
.A2(n_205),
.B1(n_213),
.B2(n_182),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_244),
.A2(n_256),
.B1(n_265),
.B2(n_165),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_126),
.B1(n_119),
.B2(n_117),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_246),
.A2(n_182),
.B1(n_198),
.B2(n_194),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_193),
.A2(n_79),
.B1(n_90),
.B2(n_89),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_172),
.A2(n_82),
.B1(n_80),
.B2(n_76),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_110),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_272),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_173),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_280),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_171),
.B(n_58),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_224),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_273),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_281),
.B(n_298),
.Y(n_325)
);

O2A1O1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_242),
.A2(n_204),
.B(n_217),
.C(n_216),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_283),
.A2(n_307),
.B(n_311),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_201),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_284),
.B(n_286),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_285),
.A2(n_276),
.B1(n_240),
.B2(n_189),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_190),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_287),
.A2(n_319),
.B1(n_283),
.B2(n_324),
.Y(n_329)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_289),
.Y(n_339)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_212),
.C(n_209),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_260),
.C(n_237),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_297),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_296),
.A2(n_274),
.B1(n_235),
.B2(n_265),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_214),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_196),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_308),
.Y(n_349)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

BUFx12_ASAP7_75t_L g301 ( 
.A(n_232),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_301),
.B(n_320),
.Y(n_341)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

BUFx12_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_185),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_304),
.B(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_258),
.Y(n_305)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_256),
.A2(n_225),
.B1(n_134),
.B2(n_196),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_306),
.A2(n_236),
.B1(n_230),
.B2(n_231),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_199),
.B(n_139),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_207),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_238),
.B(n_224),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_312),
.B(n_313),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_223),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_280),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_315),
.B(n_316),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_248),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_278),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_317),
.Y(n_360)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_323),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_238),
.A2(n_112),
.B1(n_127),
.B2(n_114),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_222),
.Y(n_320)
);

INVx13_ASAP7_75t_L g321 ( 
.A(n_237),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_251),
.Y(n_363)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g324 ( 
.A(n_274),
.B(n_207),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_324),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_308),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_350),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_327),
.A2(n_342),
.B1(n_354),
.B2(n_271),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_274),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_356),
.C(n_319),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_329),
.A2(n_294),
.B1(n_282),
.B2(n_315),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_286),
.A2(n_241),
.B(n_240),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_331),
.A2(n_314),
.B(n_317),
.Y(n_376)
);

AO21x1_ASAP7_75t_L g372 ( 
.A1(n_332),
.A2(n_294),
.B(n_297),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_324),
.A2(n_252),
.B1(n_247),
.B2(n_206),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_345),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_324),
.A2(n_252),
.B1(n_247),
.B2(n_127),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_294),
.A2(n_114),
.B1(n_236),
.B2(n_267),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_291),
.A2(n_253),
.B1(n_267),
.B2(n_258),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_203),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_318),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_296),
.A2(n_59),
.B1(n_72),
.B2(n_57),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_286),
.B(n_260),
.C(n_197),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_253),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_282),
.Y(n_365)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_365),
.Y(n_418)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_355),
.Y(n_366)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_366),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_351),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_386),
.Y(n_401)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_370),
.A2(n_373),
.B1(n_390),
.B2(n_394),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_281),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_374),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_372),
.A2(n_381),
.B(n_388),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_329),
.A2(n_283),
.B1(n_284),
.B2(n_306),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_284),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_314),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_380),
.C(n_392),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_335),
.B(n_343),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_377),
.B(n_378),
.Y(n_419)
);

OAI32xp33_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_310),
.A3(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_379)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_379),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_323),
.C(n_302),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_332),
.A2(n_305),
.B(n_285),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_309),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_385),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_384),
.A2(n_345),
.B1(n_364),
.B2(n_340),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_292),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_360),
.B(n_301),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_301),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_387),
.B(n_391),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_362),
.A2(n_301),
.B(n_261),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_331),
.A2(n_322),
.B1(n_271),
.B2(n_249),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_325),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_321),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_398),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_362),
.A2(n_249),
.B1(n_322),
.B2(n_177),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_335),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_336),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_337),
.Y(n_412)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_355),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_344),
.B(n_184),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_346),
.Y(n_402)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_404),
.C(n_423),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_356),
.C(n_328),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_353),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_303),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_373),
.A2(n_354),
.B1(n_364),
.B2(n_342),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_408),
.A2(n_361),
.B1(n_369),
.B2(n_220),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_388),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_415),
.Y(n_436)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_383),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_333),
.Y(n_416)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_351),
.Y(n_420)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_420),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_385),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_421),
.B(n_430),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_375),
.C(n_377),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_368),
.B1(n_397),
.B2(n_412),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_372),
.B(n_321),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_426),
.B(n_381),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_376),
.B(n_339),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_427),
.B(n_431),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_357),
.C(n_334),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_26),
.C(n_1),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_382),
.B(n_357),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_432),
.A2(n_26),
.B(n_2),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_433),
.A2(n_439),
.B1(n_440),
.B2(n_438),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_365),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_441),
.C(n_458),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_405),
.A2(n_384),
.B1(n_396),
.B2(n_382),
.Y(n_437)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_412),
.A2(n_368),
.B1(n_396),
.B2(n_379),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_424),
.A2(n_394),
.B1(n_395),
.B2(n_389),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_361),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_445),
.A2(n_425),
.B1(n_410),
.B2(n_411),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_405),
.A2(n_191),
.B1(n_261),
.B2(n_203),
.Y(n_446)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_446),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_408),
.A2(n_229),
.B1(n_34),
.B2(n_346),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_448),
.B(n_455),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_452),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_414),
.A2(n_34),
.B1(n_346),
.B2(n_38),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_303),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_419),
.B(n_300),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_429),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_418),
.A2(n_34),
.B1(n_38),
.B2(n_139),
.Y(n_455)
);

OAI22x1_ASAP7_75t_SL g456 ( 
.A1(n_406),
.A2(n_300),
.B1(n_228),
.B2(n_2),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_456),
.A2(n_410),
.B1(n_428),
.B2(n_431),
.Y(n_463)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_401),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_457),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_26),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_409),
.C(n_427),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_463),
.A2(n_478),
.B1(n_479),
.B2(n_469),
.Y(n_494)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_454),
.A2(n_409),
.B(n_418),
.C(n_420),
.Y(n_465)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_466),
.B(n_473),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_444),
.A2(n_426),
.B1(n_406),
.B2(n_407),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_474),
.Y(n_485)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_468),
.B(n_453),
.CI(n_441),
.CON(n_484),
.SN(n_484)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_413),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_461),
.C(n_468),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_447),
.B(n_435),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_436),
.A2(n_450),
.B1(n_445),
.B2(n_456),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_400),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_477),
.Y(n_499)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_433),
.A2(n_439),
.B1(n_432),
.B2(n_413),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_442),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_481),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_459),
.A2(n_422),
.B1(n_417),
.B2(n_428),
.Y(n_481)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_482),
.A2(n_3),
.B(n_4),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_490),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_442),
.B(n_449),
.Y(n_486)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_479),
.A2(n_458),
.B(n_443),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_487),
.B(n_493),
.Y(n_509)
);

BUFx12_ASAP7_75t_L g488 ( 
.A(n_482),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_492),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_477),
.A2(n_443),
.B(n_2),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_461),
.Y(n_504)
);

BUFx12_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_478),
.A2(n_0),
.B(n_3),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_494),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_3),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_495),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_5),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_474),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_5),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_462),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_501),
.B(n_506),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_510),
.C(n_512),
.Y(n_519)
);

OAI321xp33_ASAP7_75t_L g505 ( 
.A1(n_499),
.A2(n_465),
.A3(n_464),
.B1(n_472),
.B2(n_475),
.C(n_470),
.Y(n_505)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_505),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_462),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_471),
.C(n_466),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_497),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_492),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_480),
.C(n_26),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_496),
.B1(n_488),
.B2(n_8),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_498),
.A2(n_483),
.B1(n_493),
.B2(n_486),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_514),
.A2(n_494),
.B1(n_484),
.B2(n_9),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_515),
.B(n_516),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_503),
.B(n_489),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_520),
.B(n_523),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_499),
.B(n_490),
.Y(n_521)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_521),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_528),
.Y(n_536)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_525),
.Y(n_531)
);

MAJx2_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_500),
.C(n_484),
.Y(n_526)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_526),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_510),
.A2(n_500),
.B(n_488),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_527),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_492),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_516),
.C(n_502),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_534),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_504),
.C(n_501),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_506),
.C(n_502),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_523),
.C(n_526),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_535),
.A2(n_518),
.B(n_519),
.Y(n_539)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_539),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_541),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_532),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_517),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_542),
.B(n_538),
.Y(n_545)
);

AOI322xp5_ASAP7_75t_L g547 ( 
.A1(n_545),
.A2(n_531),
.A3(n_530),
.B1(n_537),
.B2(n_543),
.C1(n_536),
.C2(n_541),
.Y(n_547)
);

A2O1A1Ixp33_ASAP7_75t_L g549 ( 
.A1(n_547),
.A2(n_548),
.B(n_544),
.C(n_7),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_546),
.B(n_517),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_11),
.B1(n_7),
.B2(n_9),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_SL g551 ( 
.A(n_550),
.B(n_6),
.C(n_9),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_10),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_10),
.Y(n_553)
);


endmodule