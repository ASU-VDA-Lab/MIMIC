module fake_ariane_695_n_1809 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1809);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1809;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_31),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_30),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_145),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_81),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_62),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_26),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_10),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_100),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_42),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_60),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_89),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_50),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_59),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_40),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_18),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_21),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_24),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_131),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_0),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_63),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_35),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_18),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_85),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_41),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_143),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_56),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_74),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_45),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_68),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_41),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_43),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_108),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_99),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_21),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_147),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_142),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_37),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_46),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_49),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_66),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_121),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_11),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_154),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_45),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_124),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_87),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_40),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_153),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_101),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_130),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_93),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_78),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_103),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_69),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_104),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_106),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_118),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_29),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_96),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_125),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_20),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_10),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_44),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_32),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_29),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_149),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_37),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_77),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_58),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_152),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_25),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_6),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_42),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_2),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_30),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_39),
.Y(n_257)
);

CKINVDCx11_ASAP7_75t_R g258 ( 
.A(n_97),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_119),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_48),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_127),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_141),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_48),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_57),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_73),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_4),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_83),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_98),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_12),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

BUFx2_ASAP7_75t_SL g273 ( 
.A(n_72),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_49),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_137),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_7),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_43),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_7),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_107),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_148),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_33),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_111),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_65),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_34),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_22),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_114),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_44),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_17),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_88),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_14),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_64),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_146),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_12),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_53),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_26),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_91),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_32),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_8),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_13),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_95),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_36),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_34),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_22),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_112),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_138),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_6),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_90),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_258),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_304),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_219),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_190),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_194),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_206),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_161),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_191),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_191),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_191),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_210),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_191),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_157),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_230),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_191),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_167),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_191),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_191),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_185),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_230),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_195),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_264),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_156),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_287),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_156),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_186),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_305),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_165),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_212),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_225),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_204),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_165),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_204),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_204),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_208),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_187),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_208),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_284),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_222),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_277),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_189),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_222),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_192),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_287),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_200),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_297),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_172),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_170),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_166),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_202),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_247),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_272),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_205),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_218),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_272),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_197),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_197),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_199),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_199),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_290),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_238),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_170),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_226),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_242),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_327),
.A2(n_299),
.B1(n_308),
.B2(n_300),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_280),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_334),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_216),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_314),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_216),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_292),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_177),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_338),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_173),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

BUFx8_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

NAND2x1_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_158),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g412 ( 
.A1(n_376),
.A2(n_307),
.B(n_226),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_371),
.B(n_168),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_321),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_333),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_321),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_333),
.B(n_207),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_271),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_316),
.B(n_307),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_326),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_377),
.B(n_271),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_329),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_315),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_358),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_331),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_332),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_332),
.Y(n_435)
);

CKINVDCx6p67_ASAP7_75t_R g436 ( 
.A(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_341),
.B(n_171),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_378),
.B(n_207),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_378),
.A2(n_183),
.B(n_174),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_343),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_345),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_379),
.B(n_207),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_345),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_313),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_310),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_348),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_440),
.B(n_335),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_407),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

NOR2x1p5_ASAP7_75t_L g461 ( 
.A(n_397),
.B(n_324),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_339),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_418),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_403),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_368),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_353),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_409),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_R g471 ( 
.A(n_431),
.B(n_322),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_409),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_406),
.B(n_342),
.C(n_330),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_406),
.A2(n_311),
.B1(n_344),
.B2(n_350),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

OAI22x1_ASAP7_75t_L g478 ( 
.A1(n_401),
.A2(n_365),
.B1(n_369),
.B2(n_382),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_423),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_420),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_446),
.A2(n_356),
.B1(n_380),
.B2(n_368),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_368),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_418),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_449),
.Y(n_486)
);

NOR2x1p5_ASAP7_75t_L g487 ( 
.A(n_436),
.B(n_354),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_417),
.A2(n_292),
.B1(n_308),
.B2(n_300),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_415),
.B(n_359),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_420),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_420),
.B(n_363),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_418),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_362),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_423),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_408),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_424),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_448),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_408),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_453),
.Y(n_506)
);

BUFx6f_ASAP7_75t_SL g507 ( 
.A(n_415),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_408),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_408),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_385),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_415),
.B(n_364),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_422),
.B(n_370),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_430),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_419),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_408),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_417),
.A2(n_384),
.B1(n_381),
.B2(n_374),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_R g522 ( 
.A(n_449),
.B(n_373),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_430),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_419),
.B(n_368),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_430),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_391),
.B(n_367),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_415),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_410),
.B(n_353),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_391),
.A2(n_248),
.B1(n_255),
.B2(n_246),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_R g540 ( 
.A(n_415),
.B(n_312),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_436),
.B(n_299),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_453),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_442),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_438),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_391),
.B(n_368),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_398),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_419),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_448),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_442),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_398),
.B(n_368),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_419),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_445),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_387),
.B(n_245),
.C(n_243),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_451),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_436),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_445),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_445),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_398),
.A2(n_211),
.B1(n_278),
.B2(n_256),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_387),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_403),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_387),
.Y(n_564)
);

OA22x2_ASAP7_75t_L g565 ( 
.A1(n_421),
.A2(n_375),
.B1(n_372),
.B2(n_361),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_394),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_398),
.B(n_159),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_414),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_410),
.A2(n_281),
.B1(n_260),
.B2(n_254),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_394),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_394),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_398),
.B(n_383),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_394),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_414),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_396),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_396),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_396),
.B(n_247),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_393),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_398),
.B(n_159),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_396),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_400),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_437),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_451),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_400),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_437),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_402),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_400),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_441),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_441),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_400),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_400),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_402),
.B(n_368),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_399),
.B(n_368),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_451),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_421),
.B(n_355),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_421),
.B(n_160),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_451),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_441),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_410),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_403),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_562),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_565),
.A2(n_547),
.B1(n_573),
.B2(n_597),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_454),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_462),
.B(n_416),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_399),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_405),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_494),
.B(n_416),
.Y(n_610)
);

INVxp67_ASAP7_75t_SL g611 ( 
.A(n_547),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_476),
.B(n_426),
.C(n_439),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_566),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_562),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_405),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_482),
.B(n_429),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_482),
.B(n_490),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_462),
.B(n_426),
.Y(n_618)
);

OAI221xp5_ASAP7_75t_L g619 ( 
.A1(n_483),
.A2(n_276),
.B1(n_182),
.B2(n_265),
.C(n_268),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_517),
.B(n_429),
.Y(n_620)
);

BUFx5_ASAP7_75t_L g621 ( 
.A(n_470),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_470),
.Y(n_623)
);

INVx8_ASAP7_75t_L g624 ( 
.A(n_468),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_532),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_564),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_491),
.B(n_486),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_467),
.B(n_444),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_484),
.B(n_444),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_490),
.B(n_435),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_566),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_L g632 ( 
.A(n_510),
.B(n_498),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_468),
.B(n_435),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_468),
.B(n_447),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_468),
.B(n_447),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_491),
.Y(n_636)
);

BUFx6f_ASAP7_75t_SL g637 ( 
.A(n_597),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_557),
.B(n_444),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_SL g639 ( 
.A(n_558),
.B(n_388),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_602),
.B(n_450),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_602),
.A2(n_439),
.B(n_450),
.C(n_428),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_571),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_585),
.B(n_450),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_597),
.B(n_421),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_564),
.Y(n_645)
);

NOR2xp67_ASAP7_75t_L g646 ( 
.A(n_521),
.B(n_413),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_473),
.B(n_531),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_454),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_527),
.B(n_421),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_531),
.B(n_421),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_510),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_580),
.B(n_401),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_527),
.B(n_428),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_572),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_546),
.A2(n_193),
.B1(n_213),
.B2(n_241),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_568),
.A2(n_301),
.B1(n_253),
.B2(n_274),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_471),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_465),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_557),
.B(n_533),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_557),
.B(n_428),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_533),
.B(n_568),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_466),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_551),
.B(n_419),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_570),
.B(n_428),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_570),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_575),
.B(n_428),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_456),
.B(n_413),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_531),
.B(n_428),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_575),
.B(n_395),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_576),
.B(n_395),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_576),
.B(n_395),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_584),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_584),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_489),
.B(n_419),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_587),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_464),
.B(n_419),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_466),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_561),
.B(n_160),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_466),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_587),
.B(n_425),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_574),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_590),
.B(n_425),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_590),
.B(n_425),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_591),
.B(n_425),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_465),
.B(n_539),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_461),
.B(n_393),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_591),
.B(n_425),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_SL g690 ( 
.A1(n_569),
.A2(n_388),
.B1(n_287),
.B2(n_303),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_601),
.B(n_464),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_601),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_488),
.B(n_404),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_506),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_538),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_577),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_577),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_542),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_567),
.A2(n_368),
.B1(n_443),
.B2(n_178),
.Y(n_699)
);

BUFx6f_ASAP7_75t_SL g700 ( 
.A(n_501),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_464),
.B(n_425),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_549),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_549),
.B(n_404),
.Y(n_703)
);

BUFx8_ASAP7_75t_L g704 ( 
.A(n_507),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_596),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_598),
.Y(n_706)
);

AOI221xp5_ASAP7_75t_L g707 ( 
.A1(n_478),
.A2(n_285),
.B1(n_295),
.B2(n_252),
.C(n_257),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_498),
.B(n_162),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_478),
.B(n_432),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_503),
.B(n_162),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_487),
.B(n_541),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_598),
.A2(n_288),
.B(n_279),
.C(n_309),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_581),
.A2(n_443),
.B1(n_158),
.B2(n_178),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_600),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_503),
.B(n_163),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_536),
.A2(n_443),
.B1(n_163),
.B2(n_164),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_578),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_600),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_L g719 ( 
.A(n_481),
.B(n_425),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_582),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_481),
.B(n_425),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_457),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_558),
.B(n_432),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_556),
.B(n_452),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_507),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_536),
.B(n_355),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_459),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_582),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_512),
.B(n_244),
.C(n_184),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_SL g730 ( 
.A(n_508),
.B(n_223),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_466),
.B(n_433),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_536),
.A2(n_443),
.B1(n_164),
.B2(n_175),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_481),
.B(n_433),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_485),
.B(n_493),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_485),
.B(n_433),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_455),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_485),
.B(n_433),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_599),
.B(n_433),
.Y(n_738)
);

BUFx8_ASAP7_75t_L g739 ( 
.A(n_507),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_493),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_455),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_536),
.A2(n_443),
.B1(n_175),
.B2(n_176),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_493),
.B(n_433),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_565),
.A2(n_443),
.B1(n_412),
.B2(n_452),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_504),
.B(n_433),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_466),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_504),
.B(n_433),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_504),
.B(n_403),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_513),
.B(n_537),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_513),
.B(n_403),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_459),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_563),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_458),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_474),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_458),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_460),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_565),
.Y(n_757)
);

NOR2x1p5_ASAP7_75t_L g758 ( 
.A(n_522),
.B(n_357),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_540),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_563),
.B(n_403),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_460),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_563),
.B(n_403),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_509),
.B(n_357),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_463),
.A2(n_412),
.B1(n_452),
.B2(n_296),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_508),
.B(n_361),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_513),
.B(n_403),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_545),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_563),
.B(n_452),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_474),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_537),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_620),
.B(n_475),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_606),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_613),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_620),
.B(n_537),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_610),
.B(n_475),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_610),
.B(n_519),
.Y(n_776)
);

AOI21xp33_ASAP7_75t_L g777 ( 
.A1(n_619),
.A2(n_495),
.B(n_479),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_648),
.B(n_520),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_604),
.B(n_479),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_SL g780 ( 
.A1(n_690),
.A2(n_176),
.B1(n_233),
.B2(n_286),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_614),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_615),
.A2(n_595),
.B(n_525),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_703),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_648),
.B(n_520),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_658),
.B(n_563),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_658),
.B(n_496),
.C(n_495),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_626),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_646),
.B(n_603),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_645),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_666),
.B(n_496),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_622),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_673),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_674),
.Y(n_793)
);

CKINVDCx11_ASAP7_75t_R g794 ( 
.A(n_711),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_631),
.Y(n_795)
);

AND2x2_ASAP7_75t_SL g796 ( 
.A(n_639),
.B(n_412),
.Y(n_796)
);

INVx5_ASAP7_75t_L g797 ( 
.A(n_726),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_676),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_622),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_623),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_692),
.B(n_497),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_652),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_625),
.B(n_603),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_723),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_625),
.B(n_702),
.C(n_682),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_668),
.B(n_497),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_687),
.B(n_636),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_624),
.B(n_603),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_630),
.A2(n_524),
.B(n_500),
.C(n_514),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_611),
.A2(n_500),
.B1(n_499),
.B2(n_502),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_763),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_694),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_611),
.A2(n_524),
.B1(n_499),
.B2(n_502),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_624),
.B(n_603),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_642),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_627),
.A2(n_534),
.B1(n_514),
.B2(n_515),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_654),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_695),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_668),
.A2(n_515),
.B1(n_530),
.B2(n_534),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_624),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_608),
.B(n_518),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_682),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_707),
.A2(n_469),
.B1(n_526),
.B2(n_535),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_607),
.B(n_372),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_726),
.B(n_583),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_660),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_637),
.A2(n_518),
.B1(n_530),
.B2(n_529),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_698),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_683),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_760),
.A2(n_529),
.B(n_528),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_609),
.B(n_630),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_605),
.B(n_528),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_605),
.B(n_550),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_657),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_722),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_618),
.B(n_519),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_727),
.B(n_550),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_751),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_633),
.B(n_603),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_754),
.B(n_554),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_769),
.B(n_554),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_670),
.B(n_555),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_623),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_671),
.B(n_555),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_672),
.B(n_559),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_SL g846 ( 
.A(n_690),
.B(n_181),
.C(n_180),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_637),
.A2(n_559),
.B1(n_523),
.B2(n_548),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_705),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_758),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_649),
.B(n_463),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_696),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_706),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_697),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_623),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_653),
.B(n_469),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_757),
.B(n_472),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_SL g857 ( 
.A(n_612),
.B(n_294),
.C(n_180),
.Y(n_857)
);

BUFx6f_ASAP7_75t_SL g858 ( 
.A(n_711),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_749),
.B(n_472),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_726),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_704),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_714),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_693),
.B(n_519),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_759),
.B(n_375),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_718),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_623),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_749),
.B(n_643),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_634),
.B(n_635),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_688),
.B(n_583),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_651),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_675),
.A2(n_593),
.B(n_592),
.C(n_589),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_700),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_651),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_651),
.Y(n_874)
);

BUFx8_ASAP7_75t_L g875 ( 
.A(n_700),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_717),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_651),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_725),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_704),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_663),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_691),
.B(n_477),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_617),
.B(n_523),
.Y(n_882)
);

INVxp33_ASAP7_75t_L g883 ( 
.A(n_709),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_720),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_616),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_730),
.B(n_523),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_711),
.B(n_586),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_644),
.B(n_765),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_662),
.A2(n_480),
.B1(n_505),
.B2(n_516),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_767),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_765),
.B(n_586),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_663),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_767),
.Y(n_893)
);

AND2x6_ASAP7_75t_L g894 ( 
.A(n_740),
.B(n_477),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_736),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_728),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_741),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_L g898 ( 
.A(n_729),
.B(n_525),
.C(n_592),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_753),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_640),
.B(n_589),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_755),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_756),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_729),
.B(n_548),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_647),
.B(n_548),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_663),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_739),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_716),
.A2(n_516),
.B1(n_480),
.B2(n_560),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_761),
.Y(n_908)
);

AND2x4_ASAP7_75t_SL g909 ( 
.A(n_725),
.B(n_223),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_661),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_638),
.A2(n_593),
.B(n_560),
.C(n_552),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_638),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_740),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_665),
.B(n_492),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_650),
.A2(n_553),
.B1(n_492),
.B2(n_552),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_681),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_684),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_667),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_SL g919 ( 
.A(n_679),
.B(n_233),
.C(n_227),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_659),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_732),
.B(n_553),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_770),
.B(n_505),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_669),
.A2(n_553),
.B1(n_544),
.B2(n_543),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_739),
.B(n_526),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_770),
.B(n_535),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_663),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_678),
.B(n_543),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_675),
.A2(n_544),
.B1(n_579),
.B2(n_181),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_742),
.B(n_227),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_708),
.B(n_179),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_678),
.Y(n_931)
);

NOR2x2_ASAP7_75t_L g932 ( 
.A(n_656),
.B(n_0),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_641),
.B(n_412),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_678),
.Y(n_934)
);

AO21x1_ASAP7_75t_L g935 ( 
.A1(n_738),
.A2(n_221),
.B(n_234),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_678),
.B(n_286),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_685),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_686),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_680),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_734),
.B(n_412),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_655),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_743),
.B(n_412),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_689),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_712),
.B(n_452),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_701),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_743),
.B(n_452),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_680),
.B(n_291),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_721),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_680),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_724),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_744),
.B(n_452),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_710),
.A2(n_579),
.B1(n_291),
.B2(n_294),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_680),
.B(n_579),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_746),
.Y(n_954)
);

BUFx5_ASAP7_75t_L g955 ( 
.A(n_621),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_748),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_802),
.B(n_715),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_811),
.B(n_452),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_773),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_863),
.B(n_746),
.Y(n_960)
);

O2A1O1Ixp5_ASAP7_75t_L g961 ( 
.A1(n_921),
.A2(n_760),
.B(n_762),
.C(n_664),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_822),
.B(n_738),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_776),
.A2(n_713),
.B1(n_747),
.B2(n_745),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_772),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_795),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_794),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_774),
.A2(n_771),
.B(n_831),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_831),
.B(n_764),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_775),
.A2(n_629),
.B(n_628),
.C(n_664),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_771),
.A2(n_677),
.B(n_719),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_811),
.B(n_764),
.Y(n_971)
);

NOR2x1_ASAP7_75t_L g972 ( 
.A(n_879),
.B(n_731),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_885),
.B(n_747),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_867),
.A2(n_782),
.B(n_942),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_812),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_783),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_836),
.B(n_746),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_818),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_802),
.B(n_744),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_797),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_918),
.A2(n_733),
.B1(n_735),
.B2(n_737),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_820),
.B(n_797),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_791),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_797),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_799),
.B(n_731),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_797),
.B(n_746),
.Y(n_986)
);

O2A1O1Ixp5_ASAP7_75t_L g987 ( 
.A1(n_904),
.A2(n_762),
.B(n_768),
.C(n_766),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_834),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_860),
.B(n_752),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_860),
.B(n_752),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_867),
.A2(n_750),
.B(n_768),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_860),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_824),
.B(n_752),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_815),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_942),
.A2(n_752),
.B(n_699),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_890),
.B(n_893),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_806),
.A2(n_269),
.B(n_250),
.C(n_259),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_820),
.B(n_579),
.Y(n_998)
);

BUFx2_ASAP7_75t_SL g999 ( 
.A(n_858),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_860),
.B(n_621),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_807),
.B(n_632),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_859),
.A2(n_632),
.B(n_511),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_R g1003 ( 
.A(n_872),
.B(n_621),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_941),
.B(n_621),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_828),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_878),
.B(n_263),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_L g1007 ( 
.A(n_846),
.B(n_249),
.C(n_262),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_809),
.A2(n_579),
.B(n_511),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_878),
.B(n_306),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_875),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_817),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_874),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_804),
.B(n_869),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_826),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_864),
.B(n_621),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_781),
.B(n_621),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_829),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_888),
.A2(n_302),
.B1(n_298),
.B2(n_273),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_787),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_858),
.B(n_579),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_780),
.B(n_298),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_868),
.B(n_302),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_930),
.B(n_223),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_789),
.B(n_579),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_919),
.B(n_293),
.C(n_261),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_792),
.B(n_1),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_880),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_875),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_859),
.A2(n_511),
.B(n_386),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_810),
.A2(n_289),
.B(n_267),
.C(n_386),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_910),
.B(n_188),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_946),
.A2(n_511),
.B(n_390),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_946),
.A2(n_511),
.B(n_390),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_842),
.A2(n_390),
.B(n_389),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_874),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_842),
.A2(n_390),
.B(n_389),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_793),
.B(n_1),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_798),
.B(n_2),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_851),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_861),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_906),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_887),
.B(n_386),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_883),
.A2(n_796),
.B1(n_929),
.B2(n_853),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_816),
.A2(n_283),
.B1(n_217),
.B2(n_215),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_810),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_805),
.B(n_251),
.Y(n_1046)
);

BUFx2_ASAP7_75t_SL g1047 ( 
.A(n_874),
.Y(n_1047)
);

BUFx2_ASAP7_75t_SL g1048 ( 
.A(n_874),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_844),
.A2(n_386),
.B(n_389),
.C(n_5),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_876),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_857),
.A2(n_825),
.B1(n_786),
.B2(n_849),
.Y(n_1051)
);

OA21x2_ASAP7_75t_L g1052 ( 
.A1(n_933),
.A2(n_389),
.B(n_235),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_835),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_887),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_920),
.B(n_838),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_924),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_825),
.B(n_251),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_777),
.A2(n_282),
.B1(n_203),
.B2(n_201),
.C(n_198),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_844),
.A2(n_845),
.B(n_940),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_924),
.B(n_232),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_845),
.A2(n_3),
.B(n_4),
.C(n_9),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_940),
.A2(n_392),
.B(n_385),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_884),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_832),
.B(n_833),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_913),
.B(n_296),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_832),
.B(n_9),
.Y(n_1066)
);

BUFx8_ASAP7_75t_L g1067 ( 
.A(n_843),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_913),
.B(n_296),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_881),
.A2(n_392),
.B(n_385),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_850),
.A2(n_855),
.B(n_821),
.C(n_779),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_909),
.B(n_912),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_L g1072 ( 
.A1(n_935),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_870),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_833),
.B(n_15),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_937),
.B(n_16),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_953),
.B(n_161),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_880),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_SL g1078 ( 
.A1(n_779),
.A2(n_16),
.B(n_17),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_830),
.A2(n_232),
.B(n_161),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_881),
.A2(n_392),
.B(n_385),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_933),
.A2(n_392),
.B(n_385),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_850),
.A2(n_19),
.B(n_23),
.C(n_24),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_777),
.A2(n_196),
.B(n_209),
.C(n_275),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_896),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_938),
.B(n_19),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_813),
.A2(n_266),
.B1(n_214),
.B2(n_220),
.Y(n_1086)
);

OR2x6_ASAP7_75t_SL g1087 ( 
.A(n_932),
.B(n_887),
.Y(n_1087)
);

INVx5_ASAP7_75t_L g1088 ( 
.A(n_894),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_924),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_897),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_901),
.A2(n_251),
.B1(n_224),
.B2(n_270),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_914),
.A2(n_392),
.B(n_385),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_778),
.B(n_228),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_827),
.B(n_236),
.Y(n_1094)
);

NOR2xp67_ASAP7_75t_SL g1095 ( 
.A(n_880),
.B(n_926),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_855),
.A2(n_229),
.B(n_231),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_784),
.B(n_237),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_837),
.A2(n_392),
.B(n_385),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_848),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_843),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_926),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_908),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_1023),
.A2(n_944),
.B(n_788),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1045),
.B(n_916),
.Y(n_1104)
);

AOI221x1_ASAP7_75t_L g1105 ( 
.A1(n_1007),
.A2(n_871),
.B1(n_889),
.B2(n_898),
.C(n_852),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1079),
.A2(n_889),
.B(n_911),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_R g1107 ( 
.A(n_1028),
.B(n_843),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_967),
.A2(n_790),
.B(n_801),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_1100),
.Y(n_1109)
);

NOR4xp25_ASAP7_75t_L g1110 ( 
.A(n_1061),
.B(n_862),
.C(n_865),
.D(n_785),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_975),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1059),
.A2(n_956),
.A3(n_948),
.B(n_945),
.Y(n_1112)
);

AND2x6_ASAP7_75t_L g1113 ( 
.A(n_980),
.B(n_953),
.Y(n_1113)
);

O2A1O1Ixp5_ASAP7_75t_L g1114 ( 
.A1(n_974),
.A2(n_886),
.B(n_936),
.C(n_947),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1021),
.A2(n_903),
.B(n_803),
.C(n_882),
.Y(n_1115)
);

AO22x2_ASAP7_75t_L g1116 ( 
.A1(n_1045),
.A2(n_902),
.B1(n_895),
.B2(n_899),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1081),
.A2(n_839),
.B(n_837),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1059),
.A2(n_819),
.B(n_900),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_974),
.A2(n_917),
.A3(n_943),
.B(n_840),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1064),
.B(n_790),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_978),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_SL g1122 ( 
.A(n_1047),
.B(n_808),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1062),
.A2(n_841),
.B(n_840),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_SL g1124 ( 
.A1(n_1070),
.A2(n_801),
.B(n_841),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_997),
.A2(n_847),
.B(n_928),
.C(n_952),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1005),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_959),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_967),
.A2(n_925),
.B1(n_891),
.B2(n_922),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_965),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1070),
.A2(n_925),
.B(n_934),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_997),
.A2(n_800),
.B(n_854),
.C(n_873),
.Y(n_1131)
);

AO21x1_ASAP7_75t_L g1132 ( 
.A1(n_1030),
.A2(n_870),
.B(n_814),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1007),
.A2(n_800),
.B(n_854),
.C(n_873),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1087),
.B(n_877),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1012),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_966),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_968),
.B(n_934),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_983),
.B(n_823),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_964),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_979),
.B(n_954),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_963),
.A2(n_970),
.B(n_981),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1025),
.A2(n_894),
.B1(n_856),
.B2(n_927),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1019),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_973),
.B(n_954),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_1076),
.B(n_905),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_976),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_962),
.B(n_877),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_970),
.A2(n_949),
.B(n_927),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_L g1149 ( 
.A(n_1003),
.B(n_955),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1062),
.A2(n_1080),
.B(n_1069),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_977),
.A2(n_926),
.B(n_939),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1013),
.B(n_856),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1055),
.B(n_931),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_969),
.A2(n_995),
.B(n_991),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1069),
.A2(n_907),
.B(n_951),
.Y(n_1155)
);

NOR4xp25_ASAP7_75t_L g1156 ( 
.A(n_1061),
.B(n_23),
.C(n_25),
.D(n_27),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1080),
.A2(n_915),
.B(n_923),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1025),
.B(n_892),
.C(n_905),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_993),
.B(n_939),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_957),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1092),
.A2(n_892),
.A3(n_950),
.B(n_955),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1092),
.A2(n_955),
.B(n_894),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_969),
.A2(n_939),
.B(n_931),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1098),
.A2(n_955),
.A3(n_894),
.B(n_866),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1098),
.A2(n_955),
.B(n_931),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1015),
.B(n_866),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1032),
.A2(n_866),
.B(n_392),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_995),
.A2(n_232),
.B(n_161),
.Y(n_1168)
);

AND2x2_ASAP7_75t_SL g1169 ( 
.A(n_980),
.B(n_161),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_999),
.B(n_232),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1030),
.A2(n_232),
.B(n_240),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1053),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1032),
.A2(n_392),
.B(n_385),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_961),
.A2(n_239),
.B(n_28),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_SL g1175 ( 
.A(n_1082),
.B(n_27),
.C(n_28),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1066),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_L g1177 ( 
.A1(n_960),
.A2(n_110),
.B(n_150),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_991),
.A2(n_105),
.B(n_144),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_SL g1179 ( 
.A1(n_1046),
.A2(n_38),
.B(n_39),
.C(n_46),
.Y(n_1179)
);

AND2x6_ASAP7_75t_L g1180 ( 
.A(n_980),
.B(n_113),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1033),
.A2(n_115),
.B(n_139),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1004),
.A2(n_70),
.B(n_129),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_988),
.B(n_38),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1099),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1096),
.A2(n_47),
.B(n_52),
.C(n_55),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1001),
.B(n_47),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1006),
.B(n_61),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_996),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1033),
.A2(n_67),
.B(n_117),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1022),
.A2(n_123),
.B(n_126),
.C(n_151),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_994),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_961),
.A2(n_987),
.B(n_1029),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1011),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1002),
.A2(n_1008),
.B(n_1029),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1002),
.A2(n_1034),
.B(n_1036),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_1074),
.A2(n_1075),
.B(n_1085),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_982),
.B(n_1054),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1014),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1009),
.B(n_985),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1067),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1017),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1071),
.B(n_1051),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_987),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1065),
.B(n_1068),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_958),
.B(n_982),
.Y(n_1205)
);

OAI22x1_ASAP7_75t_L g1206 ( 
.A1(n_1089),
.A2(n_1057),
.B1(n_972),
.B2(n_1097),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_1010),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1083),
.A2(n_1082),
.B(n_1072),
.C(n_1018),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1039),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1016),
.A2(n_1088),
.B(n_1052),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1072),
.C(n_1093),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1049),
.A2(n_1026),
.B(n_1038),
.C(n_1037),
.Y(n_1212)
);

BUFx12f_ASAP7_75t_L g1213 ( 
.A(n_1040),
.Y(n_1213)
);

OR2x6_ASAP7_75t_L g1214 ( 
.A(n_1060),
.B(n_1056),
.Y(n_1214)
);

OA22x2_ASAP7_75t_L g1215 ( 
.A1(n_1060),
.A2(n_1094),
.B1(n_971),
.B2(n_1078),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1067),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1060),
.B(n_1042),
.Y(n_1217)
);

INVx6_ASAP7_75t_L g1218 ( 
.A(n_1041),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1042),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1088),
.A2(n_1044),
.B1(n_1058),
.B2(n_1086),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1024),
.A2(n_986),
.B(n_989),
.C(n_990),
.Y(n_1221)
);

AOI221x1_ASAP7_75t_L g1222 ( 
.A1(n_984),
.A2(n_992),
.B1(n_1073),
.B2(n_1102),
.C(n_1063),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1027),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1052),
.A2(n_1000),
.B(n_992),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_984),
.A2(n_1073),
.B(n_1043),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1091),
.A2(n_1088),
.B(n_998),
.C(n_1095),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_SL g1227 ( 
.A1(n_998),
.A2(n_1048),
.B(n_1088),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1012),
.A2(n_1035),
.B(n_1027),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1035),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1050),
.A2(n_1084),
.A3(n_1090),
.B(n_1020),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1027),
.A2(n_1077),
.B(n_1101),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1077),
.A2(n_1059),
.B(n_967),
.Y(n_1232)
);

AO21x2_ASAP7_75t_L g1233 ( 
.A1(n_1077),
.A2(n_1081),
.B(n_1062),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1101),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1101),
.B(n_607),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1012),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_975),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1070),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1070),
.A2(n_771),
.B(n_831),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1021),
.A2(n_639),
.B1(n_610),
.B2(n_846),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_982),
.B(n_820),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1021),
.B(n_501),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1079),
.A2(n_1081),
.B(n_1062),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_983),
.B(n_607),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_SL g1245 ( 
.A1(n_960),
.A2(n_1046),
.B(n_1057),
.C(n_377),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1070),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_975),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1079),
.A2(n_1081),
.B(n_1062),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_993),
.Y(n_1249)
);

BUFx2_ASAP7_75t_SL g1250 ( 
.A(n_1200),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1194),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1199),
.B(n_1188),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1217),
.B(n_1231),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1218),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1111),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1240),
.A2(n_1175),
.B1(n_1242),
.B2(n_1176),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1154),
.A2(n_1150),
.B(n_1195),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1140),
.Y(n_1258)
);

AO21x1_ASAP7_75t_L g1259 ( 
.A1(n_1212),
.A2(n_1174),
.B(n_1204),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_1141),
.A2(n_1246),
.B(n_1238),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1211),
.A2(n_1239),
.B(n_1174),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1149),
.A2(n_1108),
.B(n_1118),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1203),
.A2(n_1168),
.B(n_1173),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_L g1264 ( 
.A(n_1109),
.B(n_1202),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1147),
.A2(n_1186),
.B1(n_1220),
.B2(n_1120),
.Y(n_1265)
);

AO22x2_ASAP7_75t_L g1266 ( 
.A1(n_1196),
.A2(n_1124),
.B1(n_1222),
.B2(n_1249),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1106),
.A2(n_1167),
.B(n_1162),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1208),
.A2(n_1125),
.B(n_1185),
.C(n_1118),
.Y(n_1268)
);

OR2x6_ASAP7_75t_L g1269 ( 
.A(n_1116),
.B(n_1214),
.Y(n_1269)
);

AND2x6_ASAP7_75t_SL g1270 ( 
.A(n_1183),
.B(n_1136),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1232),
.A2(n_1123),
.B(n_1210),
.Y(n_1271)
);

AOI21xp33_ASAP7_75t_L g1272 ( 
.A1(n_1206),
.A2(n_1115),
.B(n_1103),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_1140),
.Y(n_1273)
);

CKINVDCx12_ASAP7_75t_R g1274 ( 
.A(n_1170),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1169),
.B(n_1241),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1235),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1120),
.A2(n_1232),
.B(n_1128),
.Y(n_1277)
);

O2A1O1Ixp5_ASAP7_75t_L g1278 ( 
.A1(n_1132),
.A2(n_1178),
.B(n_1114),
.C(n_1131),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1121),
.Y(n_1279)
);

OAI211xp5_ASAP7_75t_SL g1280 ( 
.A1(n_1186),
.A2(n_1176),
.B(n_1187),
.C(n_1247),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1165),
.A2(n_1157),
.B(n_1155),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1218),
.Y(n_1282)
);

AOI221x1_ASAP7_75t_L g1283 ( 
.A1(n_1171),
.A2(n_1116),
.B1(n_1103),
.B2(n_1190),
.C(n_1163),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1224),
.A2(n_1117),
.B(n_1148),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1107),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1181),
.A2(n_1189),
.B(n_1192),
.Y(n_1286)
);

OAI221xp5_ASAP7_75t_L g1287 ( 
.A1(n_1156),
.A2(n_1110),
.B1(n_1142),
.B2(n_1133),
.C(n_1134),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1146),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1126),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1145),
.A2(n_1142),
.B(n_1130),
.C(n_1104),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_L g1291 ( 
.A(n_1156),
.B(n_1179),
.C(n_1245),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1128),
.A2(n_1105),
.A3(n_1137),
.B(n_1104),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1110),
.A2(n_1233),
.B(n_1137),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1143),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1112),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1233),
.A2(n_1226),
.B(n_1225),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1136),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1158),
.A2(n_1144),
.B(n_1151),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_SL g1299 ( 
.A1(n_1144),
.A2(n_1122),
.B(n_1221),
.Y(n_1299)
);

AND2x2_ASAP7_75t_SL g1300 ( 
.A(n_1145),
.B(n_1216),
.Y(n_1300)
);

INVxp67_ASAP7_75t_SL g1301 ( 
.A(n_1153),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1166),
.A2(n_1182),
.B(n_1159),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1119),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1215),
.B(n_1158),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1153),
.A2(n_1159),
.B(n_1138),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1119),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1119),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1172),
.A2(n_1184),
.B(n_1237),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1244),
.B(n_1152),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1160),
.A2(n_1193),
.B1(n_1198),
.B2(n_1191),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1177),
.A2(n_1231),
.B(n_1201),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1170),
.A2(n_1229),
.B(n_1236),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1205),
.B(n_1139),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1223),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1219),
.B(n_1214),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1161),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1113),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1192),
.A2(n_1227),
.B(n_1228),
.Y(n_1318)
);

OAI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1170),
.A2(n_1214),
.B1(n_1234),
.B2(n_1229),
.C(n_1135),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1135),
.A2(n_1236),
.B1(n_1241),
.B2(n_1213),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1164),
.A2(n_1161),
.B(n_1127),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1180),
.A2(n_1113),
.B(n_1197),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1129),
.Y(n_1323)
);

INVx3_ASAP7_75t_SL g1324 ( 
.A(n_1207),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1209),
.A2(n_1180),
.B1(n_1113),
.B2(n_1197),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1230),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1180),
.A2(n_1113),
.B1(n_1207),
.B2(n_1230),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1180),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1164),
.A2(n_1248),
.B(n_1243),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1161),
.A2(n_1248),
.B(n_1243),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1199),
.B(n_1188),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1111),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1112),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1223),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1211),
.A2(n_620),
.B(n_1045),
.C(n_1208),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1235),
.Y(n_1336)
);

CKINVDCx14_ASAP7_75t_R g1337 ( 
.A(n_1107),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1240),
.A2(n_780),
.B1(n_846),
.B2(n_707),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1169),
.B(n_797),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1199),
.B(n_1188),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1235),
.Y(n_1341)
);

INVx4_ASAP7_75t_SL g1342 ( 
.A(n_1180),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1204),
.A2(n_610),
.B(n_776),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1164),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1194),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1210),
.A2(n_1194),
.B(n_1110),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1204),
.A2(n_610),
.B(n_776),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1240),
.A2(n_1045),
.B1(n_610),
.B2(n_1242),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1164),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1204),
.A2(n_610),
.B(n_776),
.Y(n_1350)
);

BUFx4f_ASAP7_75t_SL g1351 ( 
.A(n_1136),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1235),
.B(n_1244),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1141),
.A2(n_1239),
.B(n_967),
.Y(n_1353)
);

NOR3xp33_ASAP7_75t_L g1354 ( 
.A(n_1240),
.B(n_1242),
.C(n_465),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1136),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1194),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1217),
.B(n_1231),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1235),
.B(n_1244),
.Y(n_1358)
);

OR2x6_ASAP7_75t_L g1359 ( 
.A(n_1116),
.B(n_1239),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1112),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1238),
.A2(n_1246),
.A3(n_1194),
.B(n_1210),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1150),
.A2(n_1195),
.B(n_1141),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1204),
.A2(n_610),
.B(n_776),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1200),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1240),
.B(n_1204),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1240),
.A2(n_780),
.B1(n_846),
.B2(n_707),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1141),
.A2(n_1239),
.B(n_967),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1199),
.B(n_1188),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1240),
.A2(n_610),
.B1(n_1156),
.B2(n_1021),
.C(n_780),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1204),
.A2(n_610),
.B(n_776),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1199),
.B(n_1188),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1111),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1111),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1204),
.A2(n_610),
.B(n_776),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1241),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1235),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1210),
.A2(n_1081),
.B(n_1168),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1194),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1140),
.B(n_1116),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1194),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1210),
.A2(n_1194),
.B(n_1110),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1194),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1309),
.B(n_1252),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1328),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1331),
.B(n_1340),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1368),
.B(n_1371),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1254),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1256),
.A2(n_1348),
.B1(n_1369),
.B2(n_1374),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1341),
.B(n_1376),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1265),
.B(n_1352),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1354),
.A2(n_1363),
.B(n_1350),
.C(n_1347),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1343),
.A2(n_1370),
.B(n_1280),
.C(n_1256),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1358),
.B(n_1313),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1254),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1308),
.Y(n_1395)
);

O2A1O1Ixp5_ASAP7_75t_L g1396 ( 
.A1(n_1261),
.A2(n_1259),
.B(n_1268),
.C(n_1353),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1258),
.B(n_1273),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1367),
.A2(n_1262),
.B(n_1268),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1257),
.A2(n_1382),
.B(n_1251),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1308),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1255),
.B(n_1279),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1308),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1342),
.B(n_1328),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1253),
.B(n_1357),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1253),
.B(n_1357),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1282),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1289),
.B(n_1294),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1332),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1338),
.A2(n_1366),
.B1(n_1335),
.B2(n_1287),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1338),
.A2(n_1366),
.B1(n_1359),
.B2(n_1337),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1290),
.A2(n_1359),
.B(n_1322),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1372),
.B(n_1373),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1300),
.B(n_1314),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1301),
.B(n_1264),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1359),
.A2(n_1337),
.B1(n_1288),
.B2(n_1290),
.Y(n_1415)
);

BUFx8_ASAP7_75t_L g1416 ( 
.A(n_1355),
.Y(n_1416)
);

O2A1O1Ixp5_ASAP7_75t_L g1417 ( 
.A1(n_1278),
.A2(n_1277),
.B(n_1304),
.C(n_1298),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1272),
.A2(n_1359),
.B(n_1304),
.C(n_1299),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1282),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1300),
.B(n_1314),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1260),
.A2(n_1266),
.B(n_1346),
.Y(n_1421)
);

O2A1O1Ixp5_ASAP7_75t_L g1422 ( 
.A1(n_1291),
.A2(n_1349),
.B(n_1344),
.C(n_1377),
.Y(n_1422)
);

AND2x6_ASAP7_75t_L g1423 ( 
.A(n_1342),
.B(n_1379),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1323),
.Y(n_1424)
);

O2A1O1Ixp5_ASAP7_75t_L g1425 ( 
.A1(n_1344),
.A2(n_1349),
.B(n_1305),
.C(n_1316),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1375),
.B(n_1334),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1275),
.A2(n_1334),
.B1(n_1364),
.B2(n_1320),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1342),
.B(n_1269),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1375),
.B(n_1334),
.Y(n_1429)
);

NOR2xp67_ASAP7_75t_L g1430 ( 
.A(n_1312),
.B(n_1319),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1260),
.A2(n_1266),
.B(n_1381),
.Y(n_1431)
);

INVx3_ASAP7_75t_SL g1432 ( 
.A(n_1364),
.Y(n_1432)
);

O2A1O1Ixp5_ASAP7_75t_L g1433 ( 
.A1(n_1344),
.A2(n_1349),
.B(n_1316),
.C(n_1303),
.Y(n_1433)
);

AOI221x1_ASAP7_75t_SL g1434 ( 
.A1(n_1351),
.A2(n_1355),
.B1(n_1270),
.B2(n_1297),
.C(n_1324),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1269),
.B(n_1315),
.Y(n_1435)
);

O2A1O1Ixp5_ASAP7_75t_L g1436 ( 
.A1(n_1303),
.A2(n_1307),
.B(n_1306),
.C(n_1333),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1269),
.B(n_1266),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1285),
.B(n_1310),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1250),
.B(n_1327),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1327),
.B(n_1325),
.Y(n_1440)
);

O2A1O1Ixp5_ASAP7_75t_L g1441 ( 
.A1(n_1306),
.A2(n_1307),
.B(n_1333),
.C(n_1295),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1339),
.A2(n_1317),
.B1(n_1297),
.B2(n_1260),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1317),
.A2(n_1302),
.B1(n_1271),
.B2(n_1362),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1257),
.A2(n_1251),
.B(n_1380),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1302),
.A2(n_1271),
.B1(n_1362),
.B2(n_1274),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1345),
.A2(n_1382),
.B(n_1380),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1293),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1302),
.A2(n_1271),
.B1(n_1362),
.B2(n_1274),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1292),
.B(n_1321),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1292),
.B(n_1311),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1346),
.A2(n_1381),
.B(n_1283),
.Y(n_1451)
);

AOI221x1_ASAP7_75t_SL g1452 ( 
.A1(n_1292),
.A2(n_1361),
.B1(n_1295),
.B2(n_1360),
.C(n_1326),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1311),
.B(n_1296),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1311),
.B(n_1296),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1360),
.A2(n_1361),
.B1(n_1318),
.B2(n_1286),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1330),
.A2(n_1286),
.B(n_1329),
.C(n_1284),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1321),
.A2(n_1281),
.B(n_1284),
.C(n_1263),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1361),
.B(n_1281),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1361),
.A2(n_1329),
.B(n_1267),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1263),
.A2(n_1330),
.B(n_1356),
.C(n_1378),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1267),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1276),
.B(n_1336),
.Y(n_1462)
);

NOR2xp67_ASAP7_75t_L g1463 ( 
.A(n_1334),
.B(n_1264),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1297),
.A2(n_1256),
.B1(n_1242),
.B2(n_1337),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1256),
.A2(n_1348),
.B1(n_1369),
.B2(n_1343),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1257),
.A2(n_1367),
.B(n_1353),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1328),
.A2(n_1261),
.B(n_1290),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1256),
.A2(n_1348),
.B1(n_1369),
.B2(n_1343),
.Y(n_1468)
);

AOI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1348),
.A2(n_1240),
.B(n_1365),
.C(n_1354),
.Y(n_1469)
);

AOI21x1_ASAP7_75t_SL g1470 ( 
.A1(n_1259),
.A2(n_1204),
.B(n_1186),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1276),
.B(n_1336),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1395),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1400),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1450),
.B(n_1437),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1402),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1397),
.B(n_1398),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1447),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1408),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1428),
.B(n_1411),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1401),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1424),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1451),
.A2(n_1421),
.B(n_1431),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1466),
.B(n_1458),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1412),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1396),
.A2(n_1467),
.B(n_1466),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1407),
.Y(n_1486)
);

BUFx2_ASAP7_75t_SL g1487 ( 
.A(n_1463),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1416),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1457),
.A2(n_1453),
.B(n_1454),
.Y(n_1490)
);

AOI21xp33_ASAP7_75t_L g1491 ( 
.A1(n_1409),
.A2(n_1469),
.B(n_1465),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1449),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1416),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1414),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1443),
.B(n_1445),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1452),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1448),
.B(n_1461),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1404),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1457),
.A2(n_1459),
.B(n_1455),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1405),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1387),
.B(n_1394),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1389),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1436),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1441),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1459),
.B(n_1471),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1462),
.B(n_1396),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1391),
.B(n_1383),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1433),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1428),
.B(n_1403),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1435),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1464),
.A2(n_1468),
.B1(n_1388),
.B2(n_1410),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1399),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1425),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1446),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1433),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1392),
.A2(n_1417),
.B(n_1467),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1425),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1422),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1387),
.B(n_1394),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1512),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1476),
.B(n_1390),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1483),
.B(n_1446),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1512),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1497),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1483),
.B(n_1446),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1475),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1483),
.B(n_1444),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1477),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1512),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1476),
.B(n_1393),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1475),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1505),
.B(n_1444),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1472),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1506),
.B(n_1430),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1506),
.B(n_1415),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1479),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1506),
.B(n_1442),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1505),
.B(n_1456),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1512),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1509),
.B(n_1423),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1473),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1514),
.Y(n_1542)
);

OAI322xp33_ASAP7_75t_L g1543 ( 
.A1(n_1511),
.A2(n_1418),
.A3(n_1427),
.B1(n_1470),
.B2(n_1406),
.C1(n_1419),
.C2(n_1432),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1477),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1511),
.A2(n_1440),
.B1(n_1438),
.B2(n_1423),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1514),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1496),
.B(n_1413),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1505),
.B(n_1490),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1496),
.B(n_1420),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1490),
.B(n_1460),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1439),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1528),
.Y(n_1552)
);

NOR5xp2_ASAP7_75t_SL g1553 ( 
.A(n_1543),
.B(n_1491),
.C(n_1470),
.D(n_1516),
.E(n_1434),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1526),
.Y(n_1554)
);

OAI21xp33_ASAP7_75t_L g1555 ( 
.A1(n_1550),
.A2(n_1491),
.B(n_1516),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1541),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1545),
.A2(n_1494),
.B1(n_1507),
.B2(n_1517),
.C(n_1513),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1526),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1521),
.B(n_1507),
.Y(n_1559)
);

CKINVDCx8_ASAP7_75t_R g1560 ( 
.A(n_1540),
.Y(n_1560)
);

OAI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1535),
.A2(n_1479),
.B1(n_1485),
.B2(n_1513),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1541),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1524),
.B(n_1502),
.Y(n_1564)
);

AOI31xp33_ASAP7_75t_L g1565 ( 
.A1(n_1545),
.A2(n_1495),
.A3(n_1488),
.B(n_1519),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1531),
.Y(n_1566)
);

OAI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1537),
.A2(n_1494),
.B1(n_1517),
.B2(n_1518),
.C(n_1492),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1523),
.A2(n_1515),
.B(n_1508),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1534),
.A2(n_1518),
.B1(n_1495),
.B2(n_1479),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_R g1570 ( 
.A(n_1524),
.B(n_1479),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1524),
.B(n_1495),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1533),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1548),
.A2(n_1423),
.B1(n_1474),
.B2(n_1510),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1528),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1548),
.A2(n_1423),
.B1(n_1490),
.B2(n_1499),
.Y(n_1575)
);

AOI331xp33_ASAP7_75t_L g1576 ( 
.A1(n_1521),
.A2(n_1484),
.A3(n_1478),
.B1(n_1486),
.B2(n_1480),
.B3(n_1481),
.C1(n_1504),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1534),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1548),
.B(n_1484),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_R g1579 ( 
.A(n_1550),
.B(n_1537),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1544),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1490),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1535),
.A2(n_1487),
.B1(n_1498),
.B2(n_1500),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1530),
.B(n_1432),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1530),
.B(n_1493),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1541),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1544),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1547),
.A2(n_1492),
.B1(n_1480),
.B2(n_1503),
.C(n_1504),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1538),
.B(n_1498),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1543),
.A2(n_1499),
.B(n_1482),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1550),
.A2(n_1515),
.B(n_1508),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1538),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1530),
.B(n_1416),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1532),
.B(n_1500),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1591),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1589),
.A2(n_1523),
.B(n_1539),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1590),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1554),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1555),
.A2(n_1565),
.B(n_1591),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1590),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1554),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1560),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1574),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1558),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1571),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1571),
.B(n_1532),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1558),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1564),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1555),
.A2(n_1549),
.B(n_1547),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1590),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1581),
.B(n_1536),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1590),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1584),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1563),
.Y(n_1613)
);

OA21x2_ASAP7_75t_L g1614 ( 
.A1(n_1568),
.A2(n_1520),
.B(n_1529),
.Y(n_1614)
);

INVx11_ASAP7_75t_L g1615 ( 
.A(n_1592),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1581),
.A2(n_1520),
.B(n_1529),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1559),
.B(n_1522),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1556),
.Y(n_1618)
);

NAND2x1_ASAP7_75t_SL g1619 ( 
.A(n_1564),
.B(n_1540),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1532),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1563),
.Y(n_1621)
);

NOR2x1_ASAP7_75t_L g1622 ( 
.A(n_1587),
.B(n_1547),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1566),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1560),
.B(n_1540),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1576),
.B(n_1522),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1566),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1583),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1586),
.B(n_1549),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1572),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1552),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1565),
.A2(n_1561),
.B(n_1575),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1627),
.Y(n_1632)
);

AOI31xp33_ASAP7_75t_L g1633 ( 
.A1(n_1631),
.A2(n_1579),
.A3(n_1569),
.B(n_1557),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_SL g1634 ( 
.A(n_1598),
.B(n_1567),
.C(n_1553),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1612),
.B(n_1552),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1612),
.B(n_1588),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1540),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1597),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1625),
.B(n_1549),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1608),
.B(n_1578),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1597),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1604),
.B(n_1588),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1600),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1594),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1600),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1625),
.B(n_1580),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1603),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1603),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1606),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1606),
.Y(n_1651)
);

AND2x4_ASAP7_75t_SL g1652 ( 
.A(n_1601),
.B(n_1540),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1604),
.B(n_1593),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1601),
.B(n_1593),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1608),
.B(n_1578),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1613),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1601),
.B(n_1522),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1628),
.B(n_1551),
.Y(n_1658)
);

AND2x4_ASAP7_75t_SL g1659 ( 
.A(n_1602),
.B(n_1540),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1628),
.B(n_1551),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1627),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1627),
.Y(n_1662)
);

CKINVDCx16_ASAP7_75t_R g1663 ( 
.A(n_1594),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1613),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1605),
.B(n_1525),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1617),
.B(n_1551),
.Y(n_1666)
);

NAND2x1_ASAP7_75t_L g1667 ( 
.A(n_1607),
.B(n_1610),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1630),
.B(n_1556),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1622),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1621),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1621),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1630),
.B(n_1562),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1623),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1632),
.B(n_1605),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1632),
.B(n_1607),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1643),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1662),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1647),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_SL g1680 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1633),
.A2(n_1669),
.B1(n_1634),
.B2(n_1598),
.C(n_1631),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1647),
.Y(n_1682)
);

NAND2x1p5_ASAP7_75t_L g1683 ( 
.A(n_1661),
.B(n_1630),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1661),
.B(n_1622),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1638),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1641),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1663),
.A2(n_1609),
.B1(n_1570),
.B2(n_1596),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1645),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1642),
.B(n_1609),
.C(n_1630),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1636),
.B(n_1620),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1636),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1642),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1694)
);

CKINVDCx16_ASAP7_75t_R g1695 ( 
.A(n_1637),
.Y(n_1695)
);

NAND2x1_ASAP7_75t_SL g1696 ( 
.A(n_1637),
.B(n_1654),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1653),
.B(n_1617),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1654),
.Y(n_1699)
);

NOR2x1p5_ASAP7_75t_SL g1700 ( 
.A(n_1644),
.B(n_1596),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1646),
.B(n_1609),
.C(n_1630),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1658),
.B(n_1660),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1653),
.B(n_1624),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1658),
.B(n_1623),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1648),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1649),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1637),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1650),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1678),
.B(n_1657),
.Y(n_1709)
);

CKINVDCx16_ASAP7_75t_R g1710 ( 
.A(n_1695),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1705),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1688),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1659),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1692),
.B(n_1615),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1675),
.B(n_1659),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1696),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1675),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1681),
.A2(n_1609),
.B1(n_1599),
.B2(n_1596),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1676),
.B(n_1667),
.Y(n_1719)
);

NAND2x1p5_ASAP7_75t_L g1720 ( 
.A(n_1694),
.B(n_1609),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1685),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1684),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1686),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1702),
.B(n_1660),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1702),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1706),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1708),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1679),
.B(n_1666),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1699),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1677),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1699),
.Y(n_1731)
);

OAI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1687),
.A2(n_1655),
.B1(n_1640),
.B2(n_1610),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1677),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1717),
.B(n_1691),
.Y(n_1734)
);

OAI21xp33_ASAP7_75t_L g1735 ( 
.A1(n_1709),
.A2(n_1682),
.B(n_1679),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1712),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1718),
.A2(n_1611),
.B1(n_1599),
.B2(n_1680),
.Y(n_1737)
);

OR2x6_ASAP7_75t_L g1738 ( 
.A(n_1717),
.B(n_1683),
.Y(n_1738)
);

OAI222xp33_ASAP7_75t_L g1739 ( 
.A1(n_1710),
.A2(n_1682),
.B1(n_1611),
.B2(n_1599),
.C1(n_1707),
.C2(n_1610),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1722),
.A2(n_1674),
.B1(n_1680),
.B2(n_1611),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1725),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1725),
.B(n_1691),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1716),
.A2(n_1690),
.B1(n_1703),
.B2(n_1701),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1732),
.A2(n_1674),
.B1(n_1693),
.B2(n_1689),
.C(n_1700),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1714),
.B(n_1615),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1716),
.A2(n_1595),
.B(n_1683),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1729),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1724),
.Y(n_1748)
);

NOR4xp25_ASAP7_75t_SL g1749 ( 
.A(n_1730),
.B(n_1700),
.C(n_1664),
.D(n_1673),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1724),
.A2(n_1703),
.B1(n_1697),
.B2(n_1694),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1731),
.A2(n_1693),
.B1(n_1657),
.B2(n_1610),
.Y(n_1751)
);

AOI322xp5_ASAP7_75t_L g1752 ( 
.A1(n_1711),
.A2(n_1665),
.A3(n_1525),
.B1(n_1527),
.B2(n_1573),
.C1(n_1698),
.C2(n_1553),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1749),
.B(n_1715),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1748),
.B(n_1715),
.Y(n_1754)
);

INVxp67_ASAP7_75t_SL g1755 ( 
.A(n_1745),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1741),
.B(n_1735),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1742),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1738),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1734),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1736),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1750),
.B(n_1714),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1747),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1743),
.B(n_1731),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_SL g1764 ( 
.A(n_1753),
.B(n_1740),
.C(n_1744),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1756),
.A2(n_1753),
.B1(n_1737),
.B2(n_1763),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1759),
.B(n_1733),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1758),
.A2(n_1752),
.B1(n_1746),
.B2(n_1751),
.C(n_1720),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1761),
.B(n_1719),
.Y(n_1768)
);

AOI322xp5_ASAP7_75t_L g1769 ( 
.A1(n_1762),
.A2(n_1721),
.A3(n_1723),
.B1(n_1727),
.B2(n_1726),
.C1(n_1739),
.C2(n_1719),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1757),
.A2(n_1728),
.B1(n_1758),
.B2(n_1738),
.Y(n_1770)
);

NAND2x1_ASAP7_75t_L g1771 ( 
.A(n_1754),
.B(n_1719),
.Y(n_1771)
);

AOI322xp5_ASAP7_75t_L g1772 ( 
.A1(n_1762),
.A2(n_1713),
.A3(n_1665),
.B1(n_1553),
.B2(n_1698),
.C1(n_1728),
.C2(n_1694),
.Y(n_1772)
);

AOI221x1_ASAP7_75t_L g1773 ( 
.A1(n_1760),
.A2(n_1713),
.B1(n_1671),
.B2(n_1651),
.C(n_1656),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1765),
.A2(n_1754),
.B1(n_1713),
.B2(n_1755),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1764),
.A2(n_1720),
.B(n_1670),
.Y(n_1775)
);

OAI21xp33_ASAP7_75t_L g1776 ( 
.A1(n_1772),
.A2(n_1720),
.B(n_1704),
.Y(n_1776)
);

O2A1O1Ixp5_ASAP7_75t_L g1777 ( 
.A1(n_1771),
.A2(n_1704),
.B(n_1672),
.C(n_1668),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1770),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1767),
.A2(n_1618),
.B1(n_1542),
.B2(n_1546),
.C(n_1582),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1778),
.B(n_1774),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1777),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1776),
.B(n_1768),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1775),
.Y(n_1783)
);

NOR3xp33_ASAP7_75t_L g1784 ( 
.A(n_1779),
.B(n_1766),
.C(n_1769),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1778),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1778),
.B(n_1773),
.C(n_1595),
.Y(n_1786)
);

AOI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1783),
.A2(n_1785),
.B(n_1781),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1786),
.A2(n_1610),
.B1(n_1618),
.B2(n_1666),
.C(n_1616),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1782),
.A2(n_1595),
.B(n_1618),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_R g1790 ( 
.A(n_1780),
.B(n_1668),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1784),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1785),
.Y(n_1792)
);

AND3x4_ASAP7_75t_L g1793 ( 
.A(n_1790),
.B(n_1672),
.C(n_1668),
.Y(n_1793)
);

AO22x2_ASAP7_75t_L g1794 ( 
.A1(n_1791),
.A2(n_1672),
.B1(n_1626),
.B2(n_1629),
.Y(n_1794)
);

NOR3xp33_ASAP7_75t_L g1795 ( 
.A(n_1787),
.B(n_1489),
.C(n_1501),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1795),
.B(n_1792),
.Y(n_1796)
);

NOR2x1_ASAP7_75t_L g1797 ( 
.A(n_1796),
.B(n_1793),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1797),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1797),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1798),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1799),
.B(n_1794),
.Y(n_1801)
);

AND2x2_ASAP7_75t_SL g1802 ( 
.A(n_1800),
.B(n_1788),
.Y(n_1802)
);

OAI22x1_ASAP7_75t_L g1803 ( 
.A1(n_1801),
.A2(n_1789),
.B1(n_1626),
.B2(n_1629),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_L g1804 ( 
.A(n_1802),
.B(n_1616),
.C(n_1489),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1803),
.B1(n_1616),
.B2(n_1614),
.Y(n_1805)
);

OAI21xp33_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1562),
.B(n_1585),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1806),
.B(n_1616),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1614),
.B1(n_1585),
.B2(n_1546),
.Y(n_1808)
);

AOI211xp5_ASAP7_75t_L g1809 ( 
.A1(n_1808),
.A2(n_1426),
.B(n_1429),
.C(n_1384),
.Y(n_1809)
);


endmodule