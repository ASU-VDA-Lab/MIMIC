module fake_jpeg_27387_n_36 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_36);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_36;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_15),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_5),
.Y(n_25)
);

OAI22x1_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_20),
.B1(n_18),
.B2(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_21),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.C(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_20),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_7),
.B(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_4),
.B1(n_11),
.B2(n_3),
.Y(n_35)
);

NAND5xp2_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_1),
.C(n_2),
.D(n_3),
.E(n_30),
.Y(n_36)
);


endmodule