module real_aes_15491_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_839, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_839;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g110 ( .A(n_0), .B(n_111), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_1), .A2(n_3), .B1(n_137), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_2), .A2(n_42), .B1(n_144), .B2(n_250), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_4), .A2(n_23), .B1(n_215), .B2(n_250), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_5), .A2(n_15), .B1(n_134), .B2(n_183), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_6), .A2(n_58), .B1(n_162), .B2(n_217), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_7), .A2(n_16), .B1(n_144), .B2(n_166), .Y(n_527) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_9), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_10), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_11), .A2(n_18), .B1(n_161), .B2(n_164), .Y(n_160) );
BUFx2_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
OR2x2_ASAP7_75t_L g799 ( .A(n_12), .B(n_38), .Y(n_799) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_13), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_14), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g815 ( .A1(n_17), .A2(n_71), .B1(n_816), .B2(n_817), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_17), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_19), .A2(n_99), .B1(n_134), .B2(n_137), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_20), .A2(n_39), .B1(n_178), .B2(n_180), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_21), .B(n_135), .Y(n_228) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_22), .A2(n_56), .B(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_24), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_25), .Y(n_622) );
INVx4_ASAP7_75t_R g539 ( .A(n_26), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_27), .B(n_141), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_28), .A2(n_46), .B1(n_194), .B2(n_196), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_29), .A2(n_65), .B1(n_794), .B2(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_29), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_30), .A2(n_52), .B1(n_134), .B2(n_196), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_31), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_32), .B(n_178), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_33), .Y(n_241) );
INVx1_ASAP7_75t_L g552 ( .A(n_34), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_35), .B(n_250), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_SL g488 ( .A1(n_36), .A2(n_140), .B(n_144), .C(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_37), .A2(n_53), .B1(n_144), .B2(n_196), .Y(n_620) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_40), .A2(n_86), .B1(n_144), .B2(n_214), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_41), .A2(n_45), .B1(n_144), .B2(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_43), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_44), .A2(n_57), .B1(n_134), .B2(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g574 ( .A(n_47), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_48), .B(n_144), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_49), .Y(n_514) );
INVx2_ASAP7_75t_L g809 ( .A(n_50), .Y(n_809) );
BUFx3_ASAP7_75t_L g114 ( .A(n_51), .Y(n_114) );
INVx1_ASAP7_75t_L g826 ( .A(n_51), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_54), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_55), .A2(n_87), .B1(n_144), .B2(n_196), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_59), .A2(n_74), .B1(n_143), .B2(n_194), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_60), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_61), .A2(n_76), .B1(n_144), .B2(n_166), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_62), .A2(n_98), .B1(n_134), .B2(n_164), .Y(n_238) );
AND2x4_ASAP7_75t_L g130 ( .A(n_63), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g153 ( .A(n_64), .Y(n_153) );
INVx1_ASAP7_75t_L g794 ( .A(n_65), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_66), .A2(n_102), .B1(n_115), .B2(n_834), .Y(n_101) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_67), .A2(n_90), .B1(n_194), .B2(n_196), .Y(n_548) );
AO22x1_ASAP7_75t_L g505 ( .A1(n_68), .A2(n_75), .B1(n_180), .B2(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g131 ( .A(n_69), .Y(n_131) );
AND2x2_ASAP7_75t_L g492 ( .A(n_70), .B(n_234), .Y(n_492) );
INVx1_ASAP7_75t_L g816 ( .A(n_71), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_72), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_73), .B(n_217), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_77), .B(n_250), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_78), .Y(n_803) );
INVx2_ASAP7_75t_L g141 ( .A(n_79), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_80), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_81), .B(n_234), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_82), .A2(n_97), .B1(n_196), .B2(n_217), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_83), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_84), .B(n_151), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_85), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_88), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_89), .B(n_234), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_91), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_92), .B(n_234), .Y(n_511) );
INVx1_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_93), .B(n_825), .Y(n_824) );
NAND2xp33_ASAP7_75t_L g231 ( .A(n_94), .B(n_135), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_95), .A2(n_168), .B(n_217), .C(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g541 ( .A(n_96), .B(n_542), .Y(n_541) );
NAND2xp33_ASAP7_75t_L g519 ( .A(n_100), .B(n_179), .Y(n_519) );
BUFx12f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_SL g837 ( .A(n_103), .Y(n_837) );
AND2x6_ASAP7_75t_L g103 ( .A(n_104), .B(n_108), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
NOR3x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .C(n_114), .Y(n_108) );
INVx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_112), .Y(n_472) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g791 ( .A(n_113), .Y(n_791) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_114), .B(n_799), .Y(n_798) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_805), .B(n_810), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_792), .B(n_800), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_117), .A2(n_801), .B1(n_802), .B2(n_804), .Y(n_800) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_471), .B1(n_473), .B2(n_790), .Y(n_118) );
INVx2_ASAP7_75t_L g818 ( .A(n_119), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_119), .B(n_820), .Y(n_819) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_380), .Y(n_119) );
NOR2x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_319), .Y(n_120) );
NAND4xp25_ASAP7_75t_L g121 ( .A(n_122), .B(n_270), .C(n_289), .D(n_300), .Y(n_121) );
O2A1O1Ixp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_201), .B(n_208), .C(n_242), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_173), .Y(n_123) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_124), .B(n_335), .C(n_336), .Y(n_334) );
AND2x2_ASAP7_75t_L g416 ( .A(n_124), .B(n_298), .Y(n_416) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_157), .Y(n_124) );
AND2x2_ASAP7_75t_L g260 ( .A(n_125), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g278 ( .A(n_125), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g295 ( .A(n_125), .Y(n_295) );
AND2x2_ASAP7_75t_L g340 ( .A(n_125), .B(n_175), .Y(n_340) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
AND2x4_ASAP7_75t_L g288 ( .A(n_126), .B(n_279), .Y(n_288) );
AO31x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_132), .A3(n_148), .B(n_154), .Y(n_126) );
AO31x2_ASAP7_75t_L g236 ( .A1(n_127), .A2(n_169), .A3(n_237), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_128), .A2(n_534), .B(n_537), .Y(n_533) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AO31x2_ASAP7_75t_L g158 ( .A1(n_129), .A2(n_159), .A3(n_169), .B(n_171), .Y(n_158) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_129), .A2(n_176), .A3(n_185), .B(n_187), .Y(n_175) );
AO31x2_ASAP7_75t_L g247 ( .A1(n_129), .A2(n_248), .A3(n_252), .B(n_253), .Y(n_247) );
AO31x2_ASAP7_75t_L g525 ( .A1(n_129), .A2(n_156), .A3(n_526), .B(n_529), .Y(n_525) );
BUFx10_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g198 ( .A(n_130), .Y(n_198) );
INVx1_ASAP7_75t_L g491 ( .A(n_130), .Y(n_491) );
BUFx10_ASAP7_75t_L g523 ( .A(n_130), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B1(n_142), .B2(n_145), .Y(n_132) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_135), .Y(n_506) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
INVx3_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
INVx2_ASAP7_75t_L g215 ( .A(n_136), .Y(n_215) );
INVx1_ASAP7_75t_L g217 ( .A(n_136), .Y(n_217) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_136), .Y(n_250) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_138), .B(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_139), .A2(n_160), .B1(n_165), .B2(n_167), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_139), .A2(n_145), .B1(n_177), .B2(n_182), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_139), .A2(n_145), .B1(n_193), .B2(n_195), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_139), .A2(n_213), .B1(n_216), .B2(n_218), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_139), .A2(n_230), .B(n_231), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_139), .A2(n_167), .B1(n_238), .B2(n_239), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_139), .A2(n_145), .B1(n_249), .B2(n_251), .Y(n_248) );
OAI22x1_ASAP7_75t_L g526 ( .A1(n_139), .A2(n_218), .B1(n_527), .B2(n_528), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_139), .A2(n_218), .B1(n_548), .B2(n_549), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_139), .A2(n_501), .B1(n_619), .B2(n_620), .Y(n_618) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_L g226 ( .A1(n_140), .A2(n_166), .B(n_227), .C(n_228), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_140), .B(n_505), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_140), .A2(n_519), .B(n_520), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_140), .A2(n_500), .B(n_505), .C(n_508), .Y(n_560) );
BUFx8_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
INVx1_ASAP7_75t_L g487 ( .A(n_141), .Y(n_487) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g164 ( .A(n_144), .Y(n_164) );
INVx4_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g501 ( .A(n_146), .Y(n_501) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g517 ( .A(n_147), .Y(n_517) );
AO31x2_ASAP7_75t_L g191 ( .A1(n_148), .A2(n_192), .A3(n_197), .B(n_199), .Y(n_191) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_148), .A2(n_533), .B(n_541), .Y(n_532) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_SL g171 ( .A(n_150), .B(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_150), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g156 ( .A(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
OAI21xp33_ASAP7_75t_L g508 ( .A1(n_151), .A2(n_491), .B(n_503), .Y(n_508) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_156), .B(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g206 ( .A(n_157), .B(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g263 ( .A(n_157), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_157), .Y(n_286) );
INVx1_ASAP7_75t_L g297 ( .A(n_157), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_157), .B(n_189), .Y(n_306) );
INVx2_ASAP7_75t_L g313 ( .A(n_157), .Y(n_313) );
INVx4_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g258 ( .A(n_158), .B(n_175), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_158), .B(n_265), .Y(n_331) );
AND2x2_ASAP7_75t_L g339 ( .A(n_158), .B(n_191), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_158), .B(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g392 ( .A(n_158), .Y(n_392) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_163), .B(n_536), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_166), .A2(n_514), .B(n_515), .C(n_516), .Y(n_513) );
INVx1_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
AOI21x1_ASAP7_75t_L g479 ( .A1(n_169), .A2(n_480), .B(n_492), .Y(n_479) );
AO31x2_ASAP7_75t_L g546 ( .A1(n_169), .A2(n_197), .A3(n_547), .B(n_551), .Y(n_546) );
BUFx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_170), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g542 ( .A(n_170), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_170), .B(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_170), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g408 ( .A(n_174), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_189), .Y(n_174) );
INVx1_ASAP7_75t_L g207 ( .A(n_175), .Y(n_207) );
INVx1_ASAP7_75t_L g265 ( .A(n_175), .Y(n_265) );
INVx2_ASAP7_75t_L g299 ( .A(n_175), .Y(n_299) );
OR2x2_ASAP7_75t_L g303 ( .A(n_175), .B(n_191), .Y(n_303) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_175), .Y(n_352) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_179), .A2(n_184), .B1(n_539), .B2(n_540), .Y(n_538) );
OAI21xp33_ASAP7_75t_SL g570 ( .A1(n_180), .A2(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AO31x2_ASAP7_75t_L g211 ( .A1(n_185), .A2(n_197), .A3(n_212), .B(n_219), .Y(n_211) );
BUFx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_186), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_SL g224 ( .A(n_186), .Y(n_224) );
INVx4_ASAP7_75t_L g234 ( .A(n_186), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_186), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_186), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g578 ( .A(n_186), .B(n_523), .Y(n_578) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g325 ( .A(n_190), .B(n_205), .Y(n_325) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_191), .Y(n_261) );
INVx2_ASAP7_75t_L g279 ( .A(n_191), .Y(n_279) );
AND2x4_ASAP7_75t_L g298 ( .A(n_191), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g386 ( .A(n_191), .Y(n_386) );
INVx2_ASAP7_75t_L g550 ( .A(n_196), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_196), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_SL g232 ( .A(n_198), .Y(n_232) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_206), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g304 ( .A(n_204), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_204), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g367 ( .A(n_205), .Y(n_367) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2x1_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_210), .B(n_222), .Y(n_317) );
INVx1_ASAP7_75t_L g415 ( .A(n_210), .Y(n_415) );
BUFx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g255 ( .A(n_211), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g269 ( .A(n_211), .B(n_247), .Y(n_269) );
AND2x4_ASAP7_75t_L g292 ( .A(n_211), .B(n_235), .Y(n_292) );
INVx2_ASAP7_75t_L g309 ( .A(n_211), .Y(n_309) );
AND2x2_ASAP7_75t_L g335 ( .A(n_211), .B(n_236), .Y(n_335) );
INVx1_ASAP7_75t_L g400 ( .A(n_211), .Y(n_400) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_215), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_218), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g360 ( .A(n_221), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_235), .Y(n_221) );
AND2x2_ASAP7_75t_L g326 ( .A(n_222), .B(n_283), .Y(n_326) );
AND2x4_ASAP7_75t_L g342 ( .A(n_222), .B(n_309), .Y(n_342) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx2_ASAP7_75t_L g336 ( .A(n_223), .Y(n_336) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_233), .Y(n_223) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_224), .A2(n_225), .B(n_233), .Y(n_257) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_229), .B(n_232), .Y(n_225) );
INVx2_ASAP7_75t_L g252 ( .A(n_234), .Y(n_252) );
NOR2x1_ASAP7_75t_L g521 ( .A(n_234), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g268 ( .A(n_235), .Y(n_268) );
INVx3_ASAP7_75t_L g274 ( .A(n_235), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_235), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_235), .B(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g308 ( .A(n_236), .B(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g432 ( .A(n_236), .Y(n_432) );
OAI33xp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_258), .A3(n_259), .B1(n_260), .B2(n_262), .B3(n_266), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2x1_ASAP7_75t_L g244 ( .A(n_245), .B(n_255), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g366 ( .A(n_246), .B(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g275 ( .A(n_247), .B(n_257), .Y(n_275) );
INVx2_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
INVx1_ASAP7_75t_L g291 ( .A(n_247), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_250), .B(n_483), .Y(n_482) );
AO31x2_ASAP7_75t_L g617 ( .A1(n_252), .A2(n_523), .A3(n_618), .B(n_621), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_255), .A2(n_311), .B1(n_314), .B2(n_318), .Y(n_310) );
OR2x2_ASAP7_75t_L g450 ( .A(n_255), .B(n_268), .Y(n_450) );
AND2x4_ASAP7_75t_L g354 ( .A(n_256), .B(n_316), .Y(n_354) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_257), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_258), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g318 ( .A(n_258), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_258), .B(n_294), .Y(n_396) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g369 ( .A(n_260), .Y(n_369) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g427 ( .A(n_263), .B(n_295), .Y(n_427) );
NAND2x1_ASAP7_75t_L g445 ( .A(n_263), .B(n_294), .Y(n_445) );
AND2x2_ASAP7_75t_L g469 ( .A(n_263), .B(n_288), .Y(n_469) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g459 ( .A(n_267), .B(n_336), .Y(n_459) );
NOR2x1p5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g393 ( .A(n_268), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g361 ( .A(n_269), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_276), .B1(n_280), .B2(n_284), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
AND2x2_ASAP7_75t_L g368 ( .A(n_273), .B(n_336), .Y(n_368) );
AND2x2_ASAP7_75t_L g405 ( .A(n_273), .B(n_354), .Y(n_405) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g280 ( .A(n_274), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_274), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g446 ( .A(n_274), .B(n_275), .Y(n_446) );
AND2x2_ASAP7_75t_L g307 ( .A(n_275), .B(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g426 ( .A(n_275), .B(n_292), .Y(n_426) );
AND2x2_ASAP7_75t_L g470 ( .A(n_275), .B(n_335), .Y(n_470) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI222xp33_ASAP7_75t_L g404 ( .A1(n_280), .A2(n_405), .B1(n_406), .B2(n_409), .C1(n_411), .C2(n_412), .Y(n_404) );
AND2x2_ASAP7_75t_L g327 ( .A(n_281), .B(n_295), .Y(n_327) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g358 ( .A(n_282), .Y(n_358) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_282), .Y(n_403) );
INVx2_ASAP7_75t_L g316 ( .A(n_283), .Y(n_316) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g373 ( .A(n_286), .Y(n_373) );
INVx2_ASAP7_75t_L g379 ( .A(n_287), .Y(n_379) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g363 ( .A(n_288), .B(n_352), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x4_ASAP7_75t_L g394 ( .A(n_291), .B(n_342), .Y(n_394) );
INVx2_ASAP7_75t_L g441 ( .A(n_291), .Y(n_441) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g384 ( .A(n_295), .B(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g418 ( .A(n_295), .B(n_303), .Y(n_418) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_298), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g430 ( .A(n_298), .B(n_346), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_305), .B(n_307), .C(n_310), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
OR2x2_ASAP7_75t_L g311 ( .A(n_303), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_304), .B(n_339), .Y(n_443) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g419 ( .A(n_306), .B(n_388), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_308), .B(n_358), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_308), .A2(n_324), .B1(n_366), .B2(n_368), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_308), .B(n_336), .Y(n_371) );
AND2x2_ASAP7_75t_L g440 ( .A(n_308), .B(n_441), .Y(n_440) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_311), .A2(n_413), .B(n_434), .C(n_437), .Y(n_433) );
INVx2_ASAP7_75t_L g346 ( .A(n_313), .Y(n_346) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g424 ( .A(n_316), .Y(n_424) );
INVx1_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_318), .A2(n_365), .B1(n_369), .B2(n_370), .Y(n_364) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_332), .C(n_355), .Y(n_319) );
AO22x1_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_326), .B1(n_327), .B2(n_328), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_325), .Y(n_458) );
OR2x2_ASAP7_75t_L g465 ( .A(n_325), .B(n_346), .Y(n_465) );
AND2x2_ASAP7_75t_L g377 ( .A(n_326), .B(n_335), .Y(n_377) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g453 ( .A(n_331), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_337), .C(n_343), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
AND2x4_ASAP7_75t_SL g411 ( .A(n_335), .B(n_354), .Y(n_411) );
INVx1_ASAP7_75t_SL g422 ( .A(n_335), .Y(n_422) );
OR2x2_ASAP7_75t_L g374 ( .A(n_336), .B(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x4_ASAP7_75t_L g351 ( .A(n_339), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g409 ( .A(n_340), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g431 ( .A(n_342), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g456 ( .A(n_342), .B(n_436), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B1(n_350), .B2(n_353), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AND2x4_ASAP7_75t_L g391 ( .A(n_347), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g413 ( .A(n_347), .Y(n_413) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g468 ( .A(n_351), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR3xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_364), .C(n_372), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_362), .Y(n_356) );
INVx1_ASAP7_75t_L g437 ( .A(n_358), .Y(n_437) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_363), .A2(n_461), .B1(n_464), .B2(n_466), .C1(n_468), .C2(n_470), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_366), .B(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g389 ( .A(n_367), .Y(n_389) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B(n_376), .C(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_438), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_404), .C(n_414), .D(n_425), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_393), .B1(n_395), .B2(n_397), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .C(n_390), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_384), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_388), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g435 ( .A(n_400), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g449 ( .A(n_401), .Y(n_449) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_402), .Y(n_467) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx3_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B(n_417), .C(n_423), .Y(n_414) );
AOI21xp33_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_419), .B(n_420), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_418), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_428), .B2(n_431), .C(n_433), .Y(n_425) );
INVx1_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
AOI31xp33_ASAP7_75t_L g447 ( .A1(n_429), .A2(n_448), .A3(n_449), .B(n_450), .Y(n_447) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_432), .Y(n_436) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_451), .C(n_460), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B1(n_444), .B2(n_446), .C(n_447), .Y(n_439) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g448 ( .A(n_446), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B1(n_457), .B2(n_459), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_690), .Y(n_474) );
NAND3xp33_ASAP7_75t_SL g475 ( .A(n_476), .B(n_593), .C(n_652), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_493), .B1(n_580), .B2(n_586), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g649 ( .A(n_478), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_478), .B(n_567), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_478), .B(n_613), .Y(n_760) );
AND2x2_ASAP7_75t_L g766 ( .A(n_478), .B(n_592), .Y(n_766) );
INVxp67_ASAP7_75t_L g771 ( .A(n_478), .Y(n_771) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g584 ( .A(n_479), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_488), .B(n_491), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B(n_486), .Y(n_481) );
BUFx4f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_487), .B(n_574), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_543), .B(n_553), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_524), .Y(n_495) );
INVx1_ASAP7_75t_L g687 ( .A(n_496), .Y(n_687) );
AND2x2_ASAP7_75t_L g716 ( .A(n_496), .B(n_678), .Y(n_716) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_509), .Y(n_496) );
AND2x2_ASAP7_75t_L g610 ( .A(n_497), .B(n_532), .Y(n_610) );
INVx1_ASAP7_75t_L g665 ( .A(n_497), .Y(n_665) );
AND2x2_ASAP7_75t_L g715 ( .A(n_497), .B(n_531), .Y(n_715) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g590 ( .A(n_498), .B(n_531), .Y(n_590) );
AND2x4_ASAP7_75t_L g734 ( .A(n_498), .B(n_532), .Y(n_734) );
AOI21x1_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_504), .B(n_507), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI21x1_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_503), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_501), .A2(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g659 ( .A(n_509), .Y(n_659) );
AND2x2_ASAP7_75t_L g728 ( .A(n_509), .B(n_532), .Y(n_728) );
AND2x2_ASAP7_75t_L g735 ( .A(n_509), .B(n_561), .Y(n_735) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g557 ( .A(n_510), .Y(n_557) );
BUFx3_ASAP7_75t_L g592 ( .A(n_510), .Y(n_592) );
AND2x2_ASAP7_75t_L g603 ( .A(n_510), .B(n_589), .Y(n_603) );
AND2x2_ASAP7_75t_L g666 ( .A(n_510), .B(n_525), .Y(n_666) );
AND2x2_ASAP7_75t_L g671 ( .A(n_510), .B(n_532), .Y(n_671) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_518), .B(n_521), .Y(n_512) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_524), .B(n_677), .Y(n_779) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
INVx2_ASAP7_75t_L g561 ( .A(n_525), .Y(n_561) );
OR2x2_ASAP7_75t_L g564 ( .A(n_525), .B(n_532), .Y(n_564) );
INVx2_ASAP7_75t_L g589 ( .A(n_525), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_525), .B(n_559), .Y(n_605) );
AND2x2_ASAP7_75t_L g678 ( .A(n_525), .B(n_532), .Y(n_678) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g606 ( .A(n_532), .Y(n_606) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_544), .B(n_641), .Y(n_787) );
BUFx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g599 ( .A(n_545), .Y(n_599) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g579 ( .A(n_546), .Y(n_579) );
AND2x2_ASAP7_75t_L g585 ( .A(n_546), .B(n_567), .Y(n_585) );
INVx1_ASAP7_75t_L g633 ( .A(n_546), .Y(n_633) );
OR2x2_ASAP7_75t_L g638 ( .A(n_546), .B(n_617), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_546), .B(n_617), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_546), .B(n_616), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_546), .B(n_584), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_562), .B(n_565), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
OR2x2_ASAP7_75t_L g563 ( .A(n_556), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g714 ( .A(n_556), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g744 ( .A(n_556), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_557), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g712 ( .A(n_557), .Y(n_712) );
OR2x2_ASAP7_75t_L g625 ( .A(n_558), .B(n_626), .Y(n_625) );
INVxp33_ASAP7_75t_L g743 ( .A(n_558), .Y(n_743) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx2_ASAP7_75t_L g647 ( .A(n_559), .Y(n_647) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g601 ( .A(n_561), .Y(n_601) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI221xp5_ASAP7_75t_SL g709 ( .A1(n_563), .A2(n_634), .B1(n_639), .B2(n_710), .C(n_713), .Y(n_709) );
OR2x2_ASAP7_75t_L g696 ( .A(n_564), .B(n_647), .Y(n_696) );
INVx2_ASAP7_75t_L g745 ( .A(n_564), .Y(n_745) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g645 ( .A(n_566), .Y(n_645) );
OR2x2_ASAP7_75t_L g648 ( .A(n_566), .B(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_566), .Y(n_689) );
OR2x2_ASAP7_75t_L g702 ( .A(n_566), .B(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_579), .Y(n_566) );
NAND2x1p5_ASAP7_75t_SL g598 ( .A(n_567), .B(n_583), .Y(n_598) );
INVx3_ASAP7_75t_L g613 ( .A(n_567), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_567), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
AND2x2_ASAP7_75t_L g717 ( .A(n_567), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g724 ( .A(n_567), .B(n_631), .Y(n_724) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_575), .B(n_578), .Y(n_569) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_585), .Y(n_580) );
AND2x2_ASAP7_75t_L g776 ( .A(n_581), .B(n_635), .Y(n_776) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g680 ( .A(n_583), .B(n_650), .Y(n_680) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g615 ( .A(n_584), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g641 ( .A(n_584), .B(n_617), .Y(n_641) );
AND2x4_ASAP7_75t_L g738 ( .A(n_585), .B(n_708), .Y(n_738) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_591), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g657 ( .A(n_590), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_591), .B(n_678), .Y(n_762) );
AND2x2_ASAP7_75t_L g769 ( .A(n_591), .B(n_729), .Y(n_769) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g694 ( .A(n_592), .Y(n_694) );
AOI321xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_607), .A3(n_623), .B1(n_624), .B2(n_627), .C(n_642), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_595), .B(n_604), .Y(n_594) );
AOI21xp33_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_600), .B(n_602), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_597), .A2(n_608), .B(n_611), .Y(n_607) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
OR2x2_ASAP7_75t_L g706 ( .A(n_598), .B(n_638), .Y(n_706) );
INVx1_ASAP7_75t_L g698 ( .A(n_599), .Y(n_698) );
INVx2_ASAP7_75t_L g683 ( .A(n_600), .Y(n_683) );
OAI32xp33_ASAP7_75t_L g786 ( .A1(n_600), .A2(n_748), .A3(n_759), .B1(n_787), .B2(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g701 ( .A(n_601), .Y(n_701) );
INVx1_ASAP7_75t_L g651 ( .A(n_602), .Y(n_651) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_SL g739 ( .A(n_603), .B(n_646), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_604), .B(n_608), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_604), .A2(n_680), .B1(n_741), .B2(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g729 ( .A(n_605), .Y(n_729) );
INVx1_ASAP7_75t_L g626 ( .A(n_606), .Y(n_626) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g711 ( .A(n_610), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_611), .B(n_628), .C(n_634), .D(n_639), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVxp67_ASAP7_75t_L g653 ( .A(n_612), .Y(n_653) );
AND2x2_ASAP7_75t_L g732 ( .A(n_612), .B(n_641), .Y(n_732) );
OR2x2_ASAP7_75t_L g741 ( .A(n_612), .B(n_615), .Y(n_741) );
AND2x2_ASAP7_75t_L g765 ( .A(n_612), .B(n_637), .Y(n_765) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g679 ( .A(n_613), .B(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g686 ( .A(n_613), .B(n_633), .Y(n_686) );
INVx1_ASAP7_75t_L g750 ( .A(n_614), .Y(n_750) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g658 ( .A(n_615), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g708 ( .A(n_615), .Y(n_708) );
INVx1_ASAP7_75t_L g650 ( .A(n_616), .Y(n_650) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g631 ( .A(n_617), .Y(n_631) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AND2x4_ASAP7_75t_L g644 ( .A(n_630), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g685 ( .A(n_630), .Y(n_685) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_632), .Y(n_749) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x2_ASAP7_75t_L g640 ( .A(n_636), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g726 ( .A(n_638), .Y(n_726) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g703 ( .A(n_641), .Y(n_703) );
AND2x2_ASAP7_75t_L g746 ( .A(n_641), .B(n_686), .Y(n_746) );
O2A1O1Ixp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_646), .B(n_648), .C(n_651), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g757 ( .A(n_646), .B(n_735), .Y(n_757) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g661 ( .A(n_649), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_667), .C(n_681), .Y(n_652) );
OAI21xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B(n_660), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_656), .A2(n_764), .B(n_767), .Y(n_763) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g677 ( .A(n_659), .Y(n_677) );
AND2x2_ASAP7_75t_L g737 ( .A(n_659), .B(n_734), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g756 ( .A(n_664), .Y(n_756) );
AND2x2_ASAP7_75t_L g782 ( .A(n_664), .B(n_745), .Y(n_782) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g670 ( .A(n_665), .Y(n_670) );
INVx2_ASAP7_75t_L g721 ( .A(n_666), .Y(n_721) );
NAND2x1_ASAP7_75t_L g755 ( .A(n_666), .B(n_756), .Y(n_755) );
AOI33xp33_ASAP7_75t_L g773 ( .A1(n_666), .A2(n_686), .A3(n_724), .B1(n_734), .B2(n_766), .B3(n_839), .Y(n_773) );
OAI22xp33_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_672), .B1(n_675), .B2(n_679), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
AND2x2_ASAP7_75t_L g700 ( .A(n_671), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_672), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
OR2x2_ASAP7_75t_L g785 ( .A(n_674), .B(n_719), .Y(n_785) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
OAI22xp33_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_684), .B1(n_687), .B2(n_688), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_685), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_685), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g707 ( .A(n_686), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g772 ( .A(n_686), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_751), .Y(n_690) );
NOR4xp25_ASAP7_75t_L g691 ( .A(n_692), .B(n_709), .C(n_730), .D(n_747), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_697), .B1(n_699), .B2(n_702), .C(n_704), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_SL g747 ( .A1(n_693), .A2(n_748), .B(n_749), .C(n_750), .Y(n_747) );
NAND2x1_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g780 ( .A(n_696), .Y(n_780) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_700), .A2(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OR2x6_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B(n_717), .C(n_720), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g759 ( .A(n_719), .B(n_760), .Y(n_759) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_719), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_725), .B2(n_727), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
OAI211xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .B(n_736), .C(n_742), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g781 ( .A1(n_734), .A2(n_782), .B1(n_783), .B2(n_784), .C(n_786), .Y(n_781) );
INVx3_ASAP7_75t_L g789 ( .A(n_734), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_736) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g748 ( .A(n_745), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_774), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_763), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_757), .B(n_758), .C(n_761), .Y(n_753) );
INVx2_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NOR3xp33_ASAP7_75t_L g777 ( .A(n_757), .B(n_778), .C(n_780), .Y(n_777) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_770), .B(n_773), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_777), .B(n_781), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g804 ( .A(n_791), .B(n_798), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_796), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_793), .B(n_797), .Y(n_801) );
INVxp67_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g827 ( .A(n_799), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g812 ( .A(n_809), .Y(n_812) );
OAI21x1_ASAP7_75t_SL g810 ( .A1(n_811), .A2(n_813), .B(n_828), .Y(n_810) );
BUFx3_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_821), .Y(n_813) );
AOI21x1_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_818), .B(n_819), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_815), .Y(n_820) );
INVx5_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
CKINVDCx8_ASAP7_75t_R g832 ( .A(n_823), .Y(n_832) );
AND2x6_ASAP7_75t_SL g823 ( .A(n_824), .B(n_827), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
INVx4_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
INVx8_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
endmodule