module fake_jpeg_13377_n_34 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_34);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_4),
.A2(n_2),
.B1(n_3),
.B2(n_1),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_10),
.A2(n_11),
.B1(n_9),
.B2(n_8),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_3),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

OAI32xp33_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_7),
.A3(n_19),
.B1(n_12),
.B2(n_14),
.Y(n_22)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_20),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_24),
.B(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_16),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_14),
.B(n_13),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_28),
.B1(n_18),
.B2(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_31),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_29),
.C(n_32),
.Y(n_34)
);


endmodule