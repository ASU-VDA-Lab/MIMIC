module real_jpeg_25246_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_2),
.A2(n_25),
.B1(n_35),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_65),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_65),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_24),
.B1(n_68),
.B2(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_3),
.A2(n_25),
.B1(n_35),
.B2(n_71),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_71),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_71),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_4),
.A2(n_25),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_4),
.A2(n_62),
.B1(n_69),
.B2(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_5),
.A2(n_25),
.B1(n_35),
.B2(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_82),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_82),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_9),
.B(n_77),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_33),
.B1(n_56),
.B2(n_57),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_9),
.A2(n_40),
.B(n_87),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_9),
.B(n_99),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_9),
.A2(n_102),
.B1(n_197),
.B2(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_35),
.B(n_212),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_11),
.A2(n_25),
.B1(n_35),
.B2(n_94),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_15),
.Y(n_133)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_15),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_19),
.B(n_113),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_100),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_20),
.A2(n_21),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_22),
.B(n_52),
.C(n_66),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_23),
.A2(n_36),
.B1(n_37),
.B2(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_23),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.A3(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_23)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_35),
.B1(n_55),
.B2(n_59),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_25),
.B(n_33),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_28),
.A2(n_29),
.B1(n_69),
.B2(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_31),
.A2(n_33),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_33),
.A2(n_57),
.B(n_89),
.C(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_33),
.B(n_90),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_33),
.B(n_200),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_35),
.A2(n_55),
.A3(n_57),
.B1(n_213),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_37)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_38),
.B(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_38),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_40),
.B1(n_87),
.B2(n_89),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_39),
.B(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_45),
.A2(n_48),
.B(n_129),
.Y(n_157)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_48),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_66),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_61),
.B(n_63),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_61),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_53),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_53),
.A2(n_98),
.B1(n_99),
.B2(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_54),
.A2(n_123),
.B1(n_154),
.B2(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_54)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_57),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_56),
.B(n_59),
.Y(n_220)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_64),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_83),
.B(n_100),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.C(n_97),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_97),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_91),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_85),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_85),
.A2(n_171),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_85),
.A2(n_179),
.B1(n_180),
.B2(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_110),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_90),
.A2(n_135),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_90),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_91),
.B(n_179),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_109),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_102),
.A2(n_130),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_102),
.A2(n_133),
.B1(n_188),
.B2(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_102),
.A2(n_104),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_127),
.B2(n_137),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_126),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_135),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_161),
.B(n_248),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_158),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_145),
.B(n_158),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_146),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_152),
.B(n_231),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_242),
.B(n_247),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_226),
.B(n_241),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_206),
.B(n_225),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_184),
.B(n_205),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_174),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_174),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_181),
.C(n_182),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_193),
.B(n_204),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_191),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_198),
.B(n_203),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_195),
.B(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_207),
.B(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_218),
.B1(n_223),
.B2(n_224),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_217),
.C(n_223),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_227),
.B(n_228),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_236),
.C(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);


endmodule