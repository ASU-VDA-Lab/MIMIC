module fake_jpeg_10573_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_8),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_21),
.B1(n_16),
.B2(n_18),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_21),
.B1(n_16),
.B2(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_63),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_21),
.B1(n_30),
.B2(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_19),
.B1(n_25),
.B2(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_28),
.B1(n_18),
.B2(n_20),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_55),
.B1(n_54),
.B2(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_19),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_73),
.B(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_31),
.B1(n_22),
.B2(n_27),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_32),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_100),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_88),
.B1(n_98),
.B2(n_103),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_85),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_87),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_90),
.Y(n_130)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_67),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_58),
.B1(n_69),
.B2(n_49),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_59),
.B1(n_50),
.B2(n_61),
.Y(n_104)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_13),
.B(n_1),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_116),
.B1(n_122),
.B2(n_13),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_35),
.B1(n_17),
.B2(n_22),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_29),
.B1(n_27),
.B2(n_2),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_10),
.B(n_1),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_43),
.B1(n_38),
.B2(n_45),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_88),
.B1(n_103),
.B2(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_45),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_100),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_100),
.C(n_102),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_137),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_160),
.B1(n_152),
.B2(n_146),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_135),
.A2(n_140),
.B(n_145),
.Y(n_165)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_143),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_43),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_138),
.B(n_142),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_97),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_117),
.B1(n_109),
.B2(n_104),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_159),
.B1(n_121),
.B2(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_93),
.B1(n_90),
.B2(n_89),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_160),
.B1(n_164),
.B2(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_150),
.B(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_77),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_128),
.B1(n_119),
.B2(n_112),
.Y(n_190)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_46),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_77),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_162),
.B(n_163),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_96),
.B1(n_95),
.B2(n_92),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_26),
.B1(n_34),
.B2(n_91),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_46),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_161),
.Y(n_191)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_112),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_105),
.A2(n_34),
.B1(n_26),
.B2(n_76),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_166),
.A2(n_180),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_118),
.B1(n_107),
.B2(n_113),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_167),
.A2(n_169),
.B1(n_186),
.B2(n_193),
.Y(n_205)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_118),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_144),
.B1(n_162),
.B2(n_159),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_187),
.B1(n_197),
.B2(n_7),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_46),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_179),
.C(n_199),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_113),
.B1(n_131),
.B2(n_111),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_196),
.B1(n_151),
.B2(n_163),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_83),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_135),
.A2(n_131),
.B(n_129),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_189),
.B(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_129),
.B1(n_125),
.B2(n_111),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_138),
.A2(n_125),
.B1(n_128),
.B2(n_119),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_139),
.B1(n_147),
.B2(n_150),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_84),
.B1(n_79),
.B2(n_34),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_7),
.B1(n_1),
.B2(n_3),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_133),
.A2(n_26),
.B1(n_0),
.B2(n_2),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_142),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_7),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_201),
.B(n_222),
.Y(n_233)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_149),
.B(n_136),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_226),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_149),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_212),
.C(n_213),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_215),
.B1(n_218),
.B2(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_216),
.B1(n_197),
.B2(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_0),
.C(n_4),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_4),
.C(n_5),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_184),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_167),
.B1(n_166),
.B2(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_224),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_6),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_9),
.B(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_170),
.B(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_175),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_11),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_175),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_179),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_246),
.C(n_249),
.Y(n_257)
);

NOR2x1p5_ASAP7_75t_SL g239 ( 
.A(n_201),
.B(n_165),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_244),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_165),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_183),
.C(n_185),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_193),
.B1(n_191),
.B2(n_198),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_191),
.C(n_172),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_205),
.C(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_251),
.C(n_204),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_181),
.C(n_196),
.Y(n_251)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_214),
.B1(n_221),
.B2(n_224),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_208),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_259),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_223),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_261),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_227),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_225),
.C(n_207),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_269),
.C(n_271),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_238),
.B1(n_236),
.B2(n_239),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_221),
.B1(n_209),
.B2(n_181),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_211),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_241),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_176),
.C(n_173),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_249),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_274),
.C(n_245),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_233),
.B(n_222),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_243),
.C(n_247),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_243),
.B1(n_252),
.B2(n_253),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_288),
.B1(n_270),
.B2(n_260),
.Y(n_293)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_265),
.B(n_241),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_287),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_188),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_289),
.C(n_292),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_253),
.B1(n_247),
.B2(n_245),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_293),
.A2(n_298),
.B1(n_219),
.B2(n_12),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_263),
.B1(n_218),
.B2(n_215),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_299),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_273),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_257),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_229),
.B1(n_226),
.B2(n_272),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_257),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_258),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_289),
.C(n_279),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_202),
.B(n_173),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_269),
.C(n_276),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_317),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_281),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_311),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_286),
.B(n_290),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_288),
.B(n_277),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_315),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_307),
.A2(n_202),
.B1(n_175),
.B2(n_219),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_305),
.B1(n_297),
.B2(n_306),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_199),
.Y(n_315)
);

INVx11_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_319),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_11),
.B(n_12),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_304),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_295),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_322),
.B(n_324),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_297),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_308),
.A2(n_296),
.B(n_303),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_316),
.B(n_309),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_313),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_331),
.B(n_333),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_322),
.A2(n_317),
.B(n_313),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_325),
.C(n_323),
.Y(n_336)
);

OAI21x1_ASAP7_75t_SL g334 ( 
.A1(n_330),
.A2(n_326),
.B(n_325),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_328),
.C(n_335),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_12),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_13),
.C(n_15),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_15),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_15),
.Y(n_342)
);


endmodule