module fake_jpeg_258_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_38),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_51),
.B1(n_49),
.B2(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_61),
.B1(n_52),
.B2(n_53),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_34),
.B1(n_37),
.B2(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_34),
.B(n_41),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_57),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_58),
.C(n_53),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_54),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_39),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_72),
.B(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_58),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_42),
.A3(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_46),
.Y(n_93)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_85),
.B1(n_10),
.B2(n_9),
.C(n_12),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_68),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_70),
.C(n_58),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_96),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_13),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_0),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_103),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_24),
.B(n_25),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_5),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_110),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_112),
.B1(n_114),
.B2(n_96),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_9),
.A3(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_16),
.B1(n_22),
.B2(n_23),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_95),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_119),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_111),
.C(n_104),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_116),
.B1(n_91),
.B2(n_109),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_108),
.C(n_110),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_124),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_27),
.B(n_28),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_29),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_33),
.Y(n_130)
);


endmodule