module real_jpeg_25286_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_0),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_0),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_0),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_0),
.B(n_35),
.Y(n_117)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_21),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_2),
.B(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_114),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_4),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_4),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_4),
.B(n_21),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx8_ASAP7_75t_SL g116 ( 
.A(n_6),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_46),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_9),
.B(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_13),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_9),
.B(n_25),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_11),
.B(n_13),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_12),
.B(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_12),
.B(n_28),
.Y(n_110)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_96),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_55),
.C(n_68),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_38),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_30),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_18),
.B(n_30),
.C(n_38),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.C(n_26),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_19),
.A2(n_20),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_31),
.B(n_33),
.C(n_34),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_39),
.B(n_49),
.C(n_50),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_52),
.B(n_54),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.C(n_67),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_92),
.C(n_93),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.C(n_82),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_75),
.C(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.C(n_87),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_111),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_107),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_107),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.CI(n_110),
.CON(n_107),
.SN(n_107)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_119),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_112),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_117),
.CI(n_118),
.CON(n_112),
.SN(n_112)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);


endmodule