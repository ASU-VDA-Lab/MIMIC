module fake_netlist_6_1764_n_5364 (n_992, n_1, n_801, n_1234, n_1199, n_741, n_1027, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_212, n_700, n_50, n_1038, n_578, n_1003, n_365, n_168, n_1237, n_1061, n_77, n_783, n_798, n_188, n_509, n_245, n_1209, n_677, n_805, n_1151, n_396, n_350, n_78, n_442, n_480, n_142, n_1009, n_62, n_1160, n_883, n_1238, n_1032, n_1247, n_893, n_1099, n_1192, n_471, n_424, n_369, n_287, n_415, n_830, n_65, n_230, n_461, n_873, n_141, n_383, n_200, n_447, n_1172, n_852, n_71, n_229, n_1078, n_250, n_544, n_1140, n_35, n_836, n_375, n_522, n_945, n_1143, n_1232, n_616, n_658, n_1119, n_428, n_641, n_822, n_693, n_1056, n_758, n_516, n_1163, n_1180, n_943, n_491, n_42, n_772, n_666, n_371, n_940, n_770, n_567, n_405, n_213, n_538, n_1106, n_886, n_343, n_953, n_1094, n_494, n_539, n_493, n_155, n_45, n_454, n_638, n_1211, n_381, n_887, n_112, n_713, n_126, n_58, n_976, n_224, n_48, n_734, n_1088, n_196, n_1231, n_917, n_574, n_9, n_907, n_6, n_14, n_659, n_407, n_913, n_808, n_867, n_1230, n_473, n_1193, n_1054, n_559, n_44, n_163, n_281, n_551, n_699, n_564, n_451, n_824, n_279, n_686, n_757, n_594, n_577, n_166, n_619, n_521, n_572, n_395, n_813, n_323, n_606, n_818, n_1123, n_92, n_513, n_645, n_331, n_916, n_483, n_102, n_608, n_261, n_630, n_32, n_541, n_512, n_121, n_433, n_792, n_476, n_2, n_219, n_264, n_263, n_1162, n_860, n_788, n_939, n_821, n_938, n_1068, n_329, n_982, n_549, n_1075, n_408, n_932, n_61, n_237, n_243, n_979, n_905, n_117, n_175, n_322, n_993, n_689, n_354, n_134, n_547, n_558, n_1064, n_634, n_136, n_966, n_764, n_692, n_733, n_1233, n_487, n_241, n_30, n_1107, n_1014, n_882, n_586, n_423, n_318, n_1111, n_715, n_1251, n_88, n_530, n_277, n_618, n_199, n_1167, n_674, n_871, n_922, n_268, n_210, n_1069, n_5, n_612, n_178, n_247, n_1165, n_355, n_702, n_347, n_1175, n_328, n_429, n_1012, n_195, n_780, n_675, n_903, n_286, n_254, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_816, n_1157, n_1188, n_877, n_604, n_825, n_728, n_1063, n_26, n_55, n_267, n_1124, n_515, n_598, n_696, n_961, n_437, n_1082, n_593, n_514, n_687, n_697, n_890, n_637, n_295, n_701, n_950, n_388, n_190, n_484, n_170, n_891, n_949, n_678, n_283, n_91, n_507, n_968, n_909, n_881, n_1008, n_760, n_590, n_63, n_362, n_148, n_161, n_22, n_462, n_1033, n_1052, n_304, n_694, n_125, n_297, n_595, n_627, n_524, n_342, n_1044, n_449, n_131, n_1208, n_1164, n_1072, n_495, n_815, n_1100, n_585, n_840, n_874, n_1128, n_382, n_673, n_1071, n_1067, n_898, n_255, n_284, n_865, n_925, n_1101, n_15, n_1026, n_38, n_289, n_615, n_1249, n_59, n_1127, n_320, n_108, n_639, n_963, n_794, n_727, n_894, n_685, n_353, n_605, n_826, n_872, n_1139, n_86, n_104, n_718, n_1018, n_542, n_847, n_644, n_682, n_851, n_305, n_72, n_996, n_532, n_173, n_413, n_791, n_510, n_837, n_79, n_948, n_704, n_977, n_1005, n_536, n_622, n_147, n_581, n_765, n_432, n_987, n_631, n_720, n_153, n_842, n_156, n_145, n_843, n_656, n_989, n_797, n_1246, n_899, n_189, n_738, n_1035, n_294, n_499, n_705, n_11, n_1004, n_1176, n_1022, n_614, n_529, n_425, n_684, n_1181, n_37, n_486, n_947, n_1117, n_1087, n_648, n_657, n_1049, n_803, n_290, n_118, n_926, n_927, n_919, n_478, n_929, n_107, n_1228, n_417, n_446, n_89, n_777, n_272, n_526, n_1183, n_69, n_293, n_53, n_458, n_1070, n_998, n_16, n_717, n_18, n_154, n_1178, n_98, n_1073, n_1000, n_796, n_252, n_1195, n_184, n_552, n_216, n_912, n_745, n_1142, n_716, n_623, n_1048, n_1201, n_884, n_731, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_312, n_66, n_958, n_292, n_1250, n_100, n_1137, n_880, n_889, n_150, n_589, n_819, n_767, n_600, n_964, n_831, n_477, n_954, n_864, n_1110, n_399, n_124, n_211, n_231, n_40, n_505, n_319, n_537, n_311, n_10, n_403, n_1080, n_723, n_596, n_123, n_546, n_562, n_1141, n_386, n_1220, n_556, n_162, n_1136, n_128, n_1125, n_970, n_642, n_995, n_276, n_1159, n_1092, n_441, n_221, n_1060, n_444, n_146, n_1252, n_1223, n_303, n_511, n_193, n_1053, n_416, n_520, n_418, n_1093, n_113, n_4, n_266, n_296, n_775, n_651, n_1153, n_439, n_217, n_518, n_1185, n_453, n_215, n_914, n_759, n_426, n_317, n_90, n_54, n_488, n_497, n_773, n_920, n_99, n_13, n_1224, n_1135, n_1169, n_1179, n_401, n_324, n_335, n_463, n_1243, n_848, n_120, n_301, n_274, n_1096, n_1091, n_36, n_983, n_427, n_496, n_906, n_688, n_1077, n_351, n_259, n_177, n_385, n_858, n_613, n_736, n_501, n_956, n_960, n_663, n_856, n_379, n_778, n_1134, n_410, n_1129, n_554, n_602, n_664, n_171, n_169, n_435, n_793, n_326, n_587, n_580, n_762, n_1030, n_1202, n_465, n_1079, n_341, n_828, n_607, n_316, n_419, n_28, n_1103, n_144, n_1203, n_820, n_951, n_106, n_725, n_952, n_999, n_358, n_160, n_186, n_0, n_368, n_575, n_994, n_732, n_974, n_392, n_724, n_1020, n_1042, n_628, n_557, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_485, n_67, n_443, n_892, n_768, n_421, n_238, n_1095, n_202, n_597, n_280, n_1187, n_610, n_1024, n_198, n_179, n_248, n_517, n_667, n_1206, n_621, n_1037, n_1115, n_750, n_901, n_468, n_923, n_504, n_183, n_1015, n_466, n_1057, n_603, n_991, n_235, n_1126, n_340, n_710, n_1108, n_1182, n_39, n_73, n_785, n_746, n_609, n_101, n_167, n_127, n_1168, n_1216, n_133, n_96, n_302, n_380, n_137, n_20, n_1190, n_397, n_122, n_34, n_218, n_1213, n_70, n_172, n_239, n_97, n_782, n_490, n_220, n_809, n_1043, n_986, n_80, n_1081, n_402, n_352, n_800, n_1084, n_1171, n_460, n_662, n_374, n_1152, n_450, n_921, n_711, n_579, n_937, n_370, n_650, n_1046, n_1145, n_330, n_1121, n_1102, n_972, n_258, n_456, n_260, n_313, n_624, n_962, n_1041, n_565, n_356, n_936, n_1186, n_1062, n_885, n_896, n_83, n_654, n_411, n_152, n_1222, n_599, n_776, n_321, n_105, n_227, n_204, n_482, n_934, n_420, n_394, n_164, n_23, n_942, n_543, n_1225, n_325, n_804, n_464, n_533, n_806, n_879, n_959, n_584, n_244, n_76, n_548, n_94, n_282, n_833, n_523, n_707, n_345, n_799, n_1155, n_139, n_41, n_273, n_787, n_1146, n_159, n_1086, n_1066, n_157, n_550, n_275, n_652, n_560, n_1241, n_569, n_737, n_1235, n_1229, n_306, n_21, n_346, n_3, n_1029, n_790, n_138, n_1210, n_49, n_299, n_1248, n_902, n_333, n_1047, n_431, n_24, n_459, n_502, n_672, n_285, n_85, n_655, n_706, n_1045, n_786, n_1236, n_834, n_19, n_29, n_75, n_743, n_766, n_430, n_1002, n_545, n_489, n_251, n_1019, n_636, n_729, n_110, n_151, n_876, n_774, n_660, n_438, n_1200, n_479, n_869, n_1154, n_1113, n_646, n_528, n_391, n_1098, n_817, n_262, n_187, n_897, n_846, n_841, n_1001, n_508, n_1050, n_1177, n_332, n_1150, n_398, n_1191, n_566, n_1023, n_1076, n_1118, n_194, n_57, n_1007, n_855, n_52, n_591, n_256, n_853, n_440, n_695, n_875, n_209, n_367, n_680, n_661, n_278, n_671, n_7, n_933, n_740, n_703, n_978, n_384, n_1217, n_751, n_749, n_310, n_969, n_988, n_1065, n_84, n_568, n_143, n_180, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_739, n_400, n_955, n_337, n_214, n_246, n_1097, n_935, n_781, n_789, n_1130, n_181, n_182, n_573, n_769, n_676, n_327, n_1120, n_832, n_555, n_389, n_814, n_669, n_176, n_114, n_300, n_222, n_747, n_74, n_1105, n_721, n_742, n_535, n_691, n_372, n_111, n_314, n_378, n_1196, n_377, n_863, n_601, n_338, n_918, n_748, n_506, n_1114, n_56, n_763, n_1147, n_360, n_119, n_957, n_895, n_866, n_1227, n_191, n_387, n_452, n_744, n_971, n_946, n_344, n_761, n_1205, n_174, n_1173, n_525, n_1116, n_611, n_1219, n_8, n_1174, n_1016, n_795, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_1083, n_109, n_445, n_930, n_888, n_1112, n_234, n_910, n_911, n_82, n_27, n_236, n_653, n_752, n_908, n_944, n_576, n_1028, n_472, n_270, n_414, n_563, n_1011, n_1215, n_25, n_93, n_839, n_708, n_668, n_626, n_990, n_779, n_1104, n_854, n_1058, n_498, n_1122, n_870, n_904, n_1253, n_709, n_366, n_103, n_1109, n_185, n_712, n_348, n_376, n_390, n_1148, n_31, n_334, n_1161, n_1085, n_232, n_46, n_1239, n_771, n_470, n_475, n_924, n_298, n_492, n_1149, n_265, n_1184, n_228, n_719, n_455, n_363, n_1090, n_592, n_829, n_1156, n_393, n_984, n_503, n_132, n_868, n_570, n_859, n_406, n_735, n_878, n_620, n_130, n_519, n_307, n_469, n_1218, n_500, n_981, n_714, n_291, n_1144, n_357, n_985, n_481, n_997, n_802, n_561, n_33, n_980, n_1198, n_436, n_116, n_409, n_1244, n_240, n_756, n_810, n_1133, n_635, n_95, n_1194, n_1051, n_253, n_583, n_249, n_201, n_1039, n_1034, n_1158, n_754, n_941, n_975, n_1031, n_115, n_553, n_43, n_849, n_753, n_467, n_269, n_359, n_973, n_1055, n_582, n_861, n_857, n_967, n_571, n_271, n_404, n_158, n_206, n_679, n_633, n_1170, n_665, n_588, n_225, n_308, n_309, n_1010, n_149, n_1040, n_915, n_632, n_1166, n_812, n_1131, n_534, n_1006, n_373, n_87, n_257, n_730, n_670, n_203, n_207, n_1089, n_205, n_1242, n_681, n_1226, n_412, n_640, n_81, n_965, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_422, n_722, n_862, n_135, n_165, n_540, n_457, n_364, n_629, n_900, n_531, n_827, n_60, n_361, n_1025, n_336, n_12, n_1013, n_192, n_51, n_649, n_1240, n_5364);

input n_992;
input n_1;
input n_801;
input n_1234;
input n_1199;
input n_741;
input n_1027;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_212;
input n_700;
input n_50;
input n_1038;
input n_578;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_77;
input n_783;
input n_798;
input n_188;
input n_509;
input n_245;
input n_1209;
input n_677;
input n_805;
input n_1151;
input n_396;
input n_350;
input n_78;
input n_442;
input n_480;
input n_142;
input n_1009;
input n_62;
input n_1160;
input n_883;
input n_1238;
input n_1032;
input n_1247;
input n_893;
input n_1099;
input n_1192;
input n_471;
input n_424;
input n_369;
input n_287;
input n_415;
input n_830;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_200;
input n_447;
input n_1172;
input n_852;
input n_71;
input n_229;
input n_1078;
input n_250;
input n_544;
input n_1140;
input n_35;
input n_836;
input n_375;
input n_522;
input n_945;
input n_1143;
input n_1232;
input n_616;
input n_658;
input n_1119;
input n_428;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_758;
input n_516;
input n_1163;
input n_1180;
input n_943;
input n_491;
input n_42;
input n_772;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_405;
input n_213;
input n_538;
input n_1106;
input n_886;
input n_343;
input n_953;
input n_1094;
input n_494;
input n_539;
input n_493;
input n_155;
input n_45;
input n_454;
input n_638;
input n_1211;
input n_381;
input n_887;
input n_112;
input n_713;
input n_126;
input n_58;
input n_976;
input n_224;
input n_48;
input n_734;
input n_1088;
input n_196;
input n_1231;
input n_917;
input n_574;
input n_9;
input n_907;
input n_6;
input n_14;
input n_659;
input n_407;
input n_913;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1054;
input n_559;
input n_44;
input n_163;
input n_281;
input n_551;
input n_699;
input n_564;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_577;
input n_166;
input n_619;
input n_521;
input n_572;
input n_395;
input n_813;
input n_323;
input n_606;
input n_818;
input n_1123;
input n_92;
input n_513;
input n_645;
input n_331;
input n_916;
input n_483;
input n_102;
input n_608;
input n_261;
input n_630;
input n_32;
input n_541;
input n_512;
input n_121;
input n_433;
input n_792;
input n_476;
input n_2;
input n_219;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_788;
input n_939;
input n_821;
input n_938;
input n_1068;
input n_329;
input n_982;
input n_549;
input n_1075;
input n_408;
input n_932;
input n_61;
input n_237;
input n_243;
input n_979;
input n_905;
input n_117;
input n_175;
input n_322;
input n_993;
input n_689;
input n_354;
input n_134;
input n_547;
input n_558;
input n_1064;
input n_634;
input n_136;
input n_966;
input n_764;
input n_692;
input n_733;
input n_1233;
input n_487;
input n_241;
input n_30;
input n_1107;
input n_1014;
input n_882;
input n_586;
input n_423;
input n_318;
input n_1111;
input n_715;
input n_1251;
input n_88;
input n_530;
input n_277;
input n_618;
input n_199;
input n_1167;
input n_674;
input n_871;
input n_922;
input n_268;
input n_210;
input n_1069;
input n_5;
input n_612;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_1175;
input n_328;
input n_429;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_903;
input n_286;
input n_254;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_816;
input n_1157;
input n_1188;
input n_877;
input n_604;
input n_825;
input n_728;
input n_1063;
input n_26;
input n_55;
input n_267;
input n_1124;
input n_515;
input n_598;
input n_696;
input n_961;
input n_437;
input n_1082;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_295;
input n_701;
input n_950;
input n_388;
input n_190;
input n_484;
input n_170;
input n_891;
input n_949;
input n_678;
input n_283;
input n_91;
input n_507;
input n_968;
input n_909;
input n_881;
input n_1008;
input n_760;
input n_590;
input n_63;
input n_362;
input n_148;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_304;
input n_694;
input n_125;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_1044;
input n_449;
input n_131;
input n_1208;
input n_1164;
input n_1072;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_840;
input n_874;
input n_1128;
input n_382;
input n_673;
input n_1071;
input n_1067;
input n_898;
input n_255;
input n_284;
input n_865;
input n_925;
input n_1101;
input n_15;
input n_1026;
input n_38;
input n_289;
input n_615;
input n_1249;
input n_59;
input n_1127;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_605;
input n_826;
input n_872;
input n_1139;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_305;
input n_72;
input n_996;
input n_532;
input n_173;
input n_413;
input n_791;
input n_510;
input n_837;
input n_79;
input n_948;
input n_704;
input n_977;
input n_1005;
input n_536;
input n_622;
input n_147;
input n_581;
input n_765;
input n_432;
input n_987;
input n_631;
input n_720;
input n_153;
input n_842;
input n_156;
input n_145;
input n_843;
input n_656;
input n_989;
input n_797;
input n_1246;
input n_899;
input n_189;
input n_738;
input n_1035;
input n_294;
input n_499;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_1022;
input n_614;
input n_529;
input n_425;
input n_684;
input n_1181;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_1087;
input n_648;
input n_657;
input n_1049;
input n_803;
input n_290;
input n_118;
input n_926;
input n_927;
input n_919;
input n_478;
input n_929;
input n_107;
input n_1228;
input n_417;
input n_446;
input n_89;
input n_777;
input n_272;
input n_526;
input n_1183;
input n_69;
input n_293;
input n_53;
input n_458;
input n_1070;
input n_998;
input n_16;
input n_717;
input n_18;
input n_154;
input n_1178;
input n_98;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_184;
input n_552;
input n_216;
input n_912;
input n_745;
input n_1142;
input n_716;
input n_623;
input n_1048;
input n_1201;
input n_884;
input n_731;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_312;
input n_66;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_880;
input n_889;
input n_150;
input n_589;
input n_819;
input n_767;
input n_600;
input n_964;
input n_831;
input n_477;
input n_954;
input n_864;
input n_1110;
input n_399;
input n_124;
input n_211;
input n_231;
input n_40;
input n_505;
input n_319;
input n_537;
input n_311;
input n_10;
input n_403;
input n_1080;
input n_723;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_386;
input n_1220;
input n_556;
input n_162;
input n_1136;
input n_128;
input n_1125;
input n_970;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_1092;
input n_441;
input n_221;
input n_1060;
input n_444;
input n_146;
input n_1252;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1053;
input n_416;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_4;
input n_266;
input n_296;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_217;
input n_518;
input n_1185;
input n_453;
input n_215;
input n_914;
input n_759;
input n_426;
input n_317;
input n_90;
input n_54;
input n_488;
input n_497;
input n_773;
input n_920;
input n_99;
input n_13;
input n_1224;
input n_1135;
input n_1169;
input n_1179;
input n_401;
input n_324;
input n_335;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_301;
input n_274;
input n_1096;
input n_1091;
input n_36;
input n_983;
input n_427;
input n_496;
input n_906;
input n_688;
input n_1077;
input n_351;
input n_259;
input n_177;
input n_385;
input n_858;
input n_613;
input n_736;
input n_501;
input n_956;
input n_960;
input n_663;
input n_856;
input n_379;
input n_778;
input n_1134;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_664;
input n_171;
input n_169;
input n_435;
input n_793;
input n_326;
input n_587;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_465;
input n_1079;
input n_341;
input n_828;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1103;
input n_144;
input n_1203;
input n_820;
input n_951;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_732;
input n_974;
input n_392;
input n_724;
input n_1020;
input n_1042;
input n_628;
input n_557;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_485;
input n_67;
input n_443;
input n_892;
input n_768;
input n_421;
input n_238;
input n_1095;
input n_202;
input n_597;
input n_280;
input n_1187;
input n_610;
input n_1024;
input n_198;
input n_179;
input n_248;
input n_517;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1115;
input n_750;
input n_901;
input n_468;
input n_923;
input n_504;
input n_183;
input n_1015;
input n_466;
input n_1057;
input n_603;
input n_991;
input n_235;
input n_1126;
input n_340;
input n_710;
input n_1108;
input n_1182;
input n_39;
input n_73;
input n_785;
input n_746;
input n_609;
input n_101;
input n_167;
input n_127;
input n_1168;
input n_1216;
input n_133;
input n_96;
input n_302;
input n_380;
input n_137;
input n_20;
input n_1190;
input n_397;
input n_122;
input n_34;
input n_218;
input n_1213;
input n_70;
input n_172;
input n_239;
input n_97;
input n_782;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_986;
input n_80;
input n_1081;
input n_402;
input n_352;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_662;
input n_374;
input n_1152;
input n_450;
input n_921;
input n_711;
input n_579;
input n_937;
input n_370;
input n_650;
input n_1046;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_972;
input n_258;
input n_456;
input n_260;
input n_313;
input n_624;
input n_962;
input n_1041;
input n_565;
input n_356;
input n_936;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_654;
input n_411;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_105;
input n_227;
input n_204;
input n_482;
input n_934;
input n_420;
input n_394;
input n_164;
input n_23;
input n_942;
input n_543;
input n_1225;
input n_325;
input n_804;
input n_464;
input n_533;
input n_806;
input n_879;
input n_959;
input n_584;
input n_244;
input n_76;
input n_548;
input n_94;
input n_282;
input n_833;
input n_523;
input n_707;
input n_345;
input n_799;
input n_1155;
input n_139;
input n_41;
input n_273;
input n_787;
input n_1146;
input n_159;
input n_1086;
input n_1066;
input n_157;
input n_550;
input n_275;
input n_652;
input n_560;
input n_1241;
input n_569;
input n_737;
input n_1235;
input n_1229;
input n_306;
input n_21;
input n_346;
input n_3;
input n_1029;
input n_790;
input n_138;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_902;
input n_333;
input n_1047;
input n_431;
input n_24;
input n_459;
input n_502;
input n_672;
input n_285;
input n_85;
input n_655;
input n_706;
input n_1045;
input n_786;
input n_1236;
input n_834;
input n_19;
input n_29;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1002;
input n_545;
input n_489;
input n_251;
input n_1019;
input n_636;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_660;
input n_438;
input n_1200;
input n_479;
input n_869;
input n_1154;
input n_1113;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_817;
input n_262;
input n_187;
input n_897;
input n_846;
input n_841;
input n_1001;
input n_508;
input n_1050;
input n_1177;
input n_332;
input n_1150;
input n_398;
input n_1191;
input n_566;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_855;
input n_52;
input n_591;
input n_256;
input n_853;
input n_440;
input n_695;
input n_875;
input n_209;
input n_367;
input n_680;
input n_661;
input n_278;
input n_671;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_384;
input n_1217;
input n_751;
input n_749;
input n_310;
input n_969;
input n_988;
input n_1065;
input n_84;
input n_568;
input n_143;
input n_180;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_739;
input n_400;
input n_955;
input n_337;
input n_214;
input n_246;
input n_1097;
input n_935;
input n_781;
input n_789;
input n_1130;
input n_181;
input n_182;
input n_573;
input n_769;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_555;
input n_389;
input n_814;
input n_669;
input n_176;
input n_114;
input n_300;
input n_222;
input n_747;
input n_74;
input n_1105;
input n_721;
input n_742;
input n_535;
input n_691;
input n_372;
input n_111;
input n_314;
input n_378;
input n_1196;
input n_377;
input n_863;
input n_601;
input n_338;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1147;
input n_360;
input n_119;
input n_957;
input n_895;
input n_866;
input n_1227;
input n_191;
input n_387;
input n_452;
input n_744;
input n_971;
input n_946;
input n_344;
input n_761;
input n_1205;
input n_174;
input n_1173;
input n_525;
input n_1116;
input n_611;
input n_1219;
input n_8;
input n_1174;
input n_1016;
input n_795;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_1083;
input n_109;
input n_445;
input n_930;
input n_888;
input n_1112;
input n_234;
input n_910;
input n_911;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_908;
input n_944;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_414;
input n_563;
input n_1011;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_708;
input n_668;
input n_626;
input n_990;
input n_779;
input n_1104;
input n_854;
input n_1058;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_366;
input n_103;
input n_1109;
input n_185;
input n_712;
input n_348;
input n_376;
input n_390;
input n_1148;
input n_31;
input n_334;
input n_1161;
input n_1085;
input n_232;
input n_46;
input n_1239;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_492;
input n_1149;
input n_265;
input n_1184;
input n_228;
input n_719;
input n_455;
input n_363;
input n_1090;
input n_592;
input n_829;
input n_1156;
input n_393;
input n_984;
input n_503;
input n_132;
input n_868;
input n_570;
input n_859;
input n_406;
input n_735;
input n_878;
input n_620;
input n_130;
input n_519;
input n_307;
input n_469;
input n_1218;
input n_500;
input n_981;
input n_714;
input n_291;
input n_1144;
input n_357;
input n_985;
input n_481;
input n_997;
input n_802;
input n_561;
input n_33;
input n_980;
input n_1198;
input n_436;
input n_116;
input n_409;
input n_1244;
input n_240;
input n_756;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_1051;
input n_253;
input n_583;
input n_249;
input n_201;
input n_1039;
input n_1034;
input n_1158;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_553;
input n_43;
input n_849;
input n_753;
input n_467;
input n_269;
input n_359;
input n_973;
input n_1055;
input n_582;
input n_861;
input n_857;
input n_967;
input n_571;
input n_271;
input n_404;
input n_158;
input n_206;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_588;
input n_225;
input n_308;
input n_309;
input n_1010;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_812;
input n_1131;
input n_534;
input n_1006;
input n_373;
input n_87;
input n_257;
input n_730;
input n_670;
input n_203;
input n_207;
input n_1089;
input n_205;
input n_1242;
input n_681;
input n_1226;
input n_412;
input n_640;
input n_81;
input n_965;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_422;
input n_722;
input n_862;
input n_135;
input n_165;
input n_540;
input n_457;
input n_364;
input n_629;
input n_900;
input n_531;
input n_827;
input n_60;
input n_361;
input n_1025;
input n_336;
input n_12;
input n_1013;
input n_192;
input n_51;
input n_649;
input n_1240;

output n_5364;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_1351;
wire n_5254;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_3089;
wire n_4978;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_4686;
wire n_2317;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1971;
wire n_1781;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_4814;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_2625;
wire n_1400;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_2764;
wire n_2895;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_5183;
wire n_2145;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1512;
wire n_1451;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_3179;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_4345;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_4528;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_5035;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_5359;
wire n_1955;
wire n_1791;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_4189;
wire n_3817;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_4512;
wire n_1378;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_3569;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_3027;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1461;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_4027;
wire n_3154;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1570;
wire n_1702;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_3552;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_5335;
wire n_3444;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_3266;
wire n_3574;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_4504;
wire n_3844;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_5248;
wire n_1708;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_2356;
wire n_1511;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_2739;
wire n_1620;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_4047;
wire n_3413;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_3725;
wire n_3933;
wire n_2311;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_1987;
wire n_2271;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_2954;
wire n_2728;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_3442;
wire n_1880;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_5087;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_3133;
wire n_1959;
wire n_5257;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_3654;
wire n_2848;
wire n_1849;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_2338;
wire n_3324;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_5282;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1951;
wire n_4362;
wire n_3311;
wire n_3913;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_4404;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4844;
wire n_4438;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_3250;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_2598;
wire n_1683;
wire n_1916;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_4016;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4192;
wire n_4109;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_5348;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_2390;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_3381;
wire n_1548;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_4170;
wire n_4143;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_3515;
wire n_2951;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_4910;
wire n_3083;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5203;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_4521;
wire n_1566;
wire n_3204;
wire n_4920;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_4730;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1517;
wire n_1867;
wire n_1393;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_2256;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_2806;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_2593;
wire n_4255;
wire n_4071;
wire n_3568;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1309;
wire n_2961;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1530;
wire n_4745;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_3599;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_3022;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_4800;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_3227;
wire n_3289;
wire n_2733;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_3326;
wire n_2036;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_4097;
wire n_1666;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_4754;
wire n_2993;
wire n_4647;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_3636;
wire n_2327;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_2755;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1692;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_2376;
wire n_1405;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_3307;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_2141;
wire n_5316;
wire n_3930;
wire n_4943;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_2021;
wire n_4942;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_3157;
wire n_4841;
wire n_3221;
wire n_1758;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_2045;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_2566;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_4913;
wire n_2312;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_2042;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_1770;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_4089;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_4865;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_3155;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_2405;
wire n_4050;
wire n_2647;
wire n_2336;
wire n_2521;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_3822;
wire n_4163;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_4372;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_4673;
wire n_2519;
wire n_3415;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_4019;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_2316;
wire n_1771;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1475;
wire n_3103;
wire n_2354;
wire n_1774;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_3144;
wire n_3244;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2357;
wire n_2025;
wire n_4654;
wire n_3640;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_2278;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_2704;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_3377;
wire n_2727;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_1794;
wire n_4493;
wire n_4924;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_2066;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1327;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_2380;
wire n_4786;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_3493;
wire n_3774;
wire n_2910;
wire n_3268;
wire n_1785;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_2287;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_3334;
wire n_5097;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_2600;
wire n_3508;
wire n_4353;
wire n_4787;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_2440;
wire n_3521;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_2909;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_4210;
wire n_4981;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_1557;
wire n_3945;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1019),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_477),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1065),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_479),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_989),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_547),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_99),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1197),
.Y(n_1261)
);

BUFx10_ASAP7_75t_L g1262 ( 
.A(n_698),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_997),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1244),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_587),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_593),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_377),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1055),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1093),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_25),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_753),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_862),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1187),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_943),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1056),
.Y(n_1275)
);

BUFx2_ASAP7_75t_SL g1276 ( 
.A(n_843),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1144),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_446),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_423),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_978),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_604),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1224),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_831),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_839),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1015),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1062),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_858),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_716),
.Y(n_1288)
);

BUFx10_ASAP7_75t_L g1289 ( 
.A(n_968),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1023),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1030),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_771),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_247),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1164),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_922),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_487),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_928),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_947),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1115),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1070),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_314),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_268),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_456),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1236),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_578),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_744),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1026),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_932),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_308),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_374),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_452),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_429),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_535),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1063),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1105),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_404),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_378),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_573),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_595),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_235),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_692),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1018),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_31),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_437),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_864),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1126),
.Y(n_1326)
);

BUFx5_ASAP7_75t_L g1327 ( 
.A(n_1129),
.Y(n_1327)
);

BUFx5_ASAP7_75t_L g1328 ( 
.A(n_261),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_896),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_688),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1190),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1179),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_151),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_956),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_693),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_387),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_868),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1231),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_708),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1232),
.Y(n_1340)
);

BUFx8_ASAP7_75t_SL g1341 ( 
.A(n_873),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_357),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_238),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_411),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1243),
.Y(n_1345)
);

BUFx10_ASAP7_75t_L g1346 ( 
.A(n_444),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_957),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_454),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_897),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_921),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_936),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1205),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_203),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_223),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1079),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_242),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_412),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_720),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_422),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_578),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1180),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_33),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_546),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_976),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_107),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1198),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_951),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1048),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_992),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_349),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1138),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1036),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1068),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_923),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_888),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1117),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_810),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1212),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1082),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_481),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_248),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_771),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1142),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_993),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_309),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_351),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1163),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_585),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_797),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1091),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_415),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1203),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_952),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1149),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1184),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_10),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_39),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_754),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_830),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_122),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1239),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_930),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_528),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1155),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1166),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_902),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_805),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1029),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1216),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_335),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_911),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_510),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1153),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_994),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_933),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_684),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_811),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1151),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_234),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_381),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1033),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_858),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_907),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1037),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1054),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_372),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_728),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_620),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_840),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1175),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_212),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1221),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_758),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_873),
.Y(n_1434)
);

BUFx10_ASAP7_75t_L g1435 ( 
.A(n_926),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_906),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_197),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_313),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_386),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_977),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_200),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_107),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1139),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1195),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_790),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_47),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_569),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_500),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1074),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_239),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1124),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_980),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_173),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_589),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_570),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_375),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_920),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1242),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_809),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_376),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1113),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_176),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1204),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_525),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_970),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_265),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1120),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1021),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1001),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1102),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_547),
.Y(n_1471)
);

BUFx2_ASAP7_75t_SL g1472 ( 
.A(n_835),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1046),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_565),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_974),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1143),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1042),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1218),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1051),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_274),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_522),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_222),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1165),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_50),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1167),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_83),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1215),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_263),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_42),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_673),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1217),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1075),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_544),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_379),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_765),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_991),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_969),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1131),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_971),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_510),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_471),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_934),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_899),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1250),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_358),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_357),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_966),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_136),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_397),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_94),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_607),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_53),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_723),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_813),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1086),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_849),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_498),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1088),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_976),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_560),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_127),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_939),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_864),
.Y(n_1523)
);

BUFx10_ASAP7_75t_L g1524 ( 
.A(n_677),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_836),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_255),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_161),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1177),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1108),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_735),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_506),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_123),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_543),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_532),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_494),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1252),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_857),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1061),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1080),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_656),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_848),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1162),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_245),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_979),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_929),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_611),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_552),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_331),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_945),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_468),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1152),
.Y(n_1551)
);

CKINVDCx16_ASAP7_75t_R g1552 ( 
.A(n_441),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_82),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_197),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_791),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_897),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1160),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_347),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_560),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_173),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1130),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_553),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_683),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1206),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1125),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_540),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1183),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_954),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1034),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_797),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1196),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_589),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1038),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1178),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_743),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_734),
.Y(n_1576)
);

BUFx10_ASAP7_75t_L g1577 ( 
.A(n_759),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_125),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1199),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_676),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_573),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_500),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_867),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_157),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_224),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_234),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1235),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_961),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_651),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_14),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1122),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_64),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1161),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_105),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_714),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_839),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1172),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_418),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_919),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1112),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1238),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1107),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_427),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_486),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_254),
.Y(n_1605)
);

BUFx10_ASAP7_75t_L g1606 ( 
.A(n_613),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_195),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1027),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_636),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_371),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_664),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_536),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_536),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_84),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1118),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1247),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_924),
.Y(n_1617)
);

BUFx10_ASAP7_75t_L g1618 ( 
.A(n_846),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1214),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1032),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_743),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_566),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_598),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_367),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_836),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1192),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1148),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1043),
.Y(n_1628)
);

CKINVDCx16_ASAP7_75t_R g1629 ( 
.A(n_271),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_727),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_93),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_455),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_831),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1223),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_89),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_257),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_678),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_773),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_608),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_27),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_261),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1003),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1092),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1154),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1207),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_722),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_937),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1241),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_100),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_125),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_829),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_942),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1100),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1084),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1085),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1181),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_935),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_838),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_65),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1140),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_813),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_998),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_746),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_226),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_218),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_279),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_867),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1171),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1017),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1186),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_139),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_681),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_666),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_315),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_283),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_120),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_667),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_744),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1111),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_123),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_264),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_257),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_431),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_676),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1189),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_593),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_135),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_18),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1066),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1209),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_555),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_946),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_820),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_962),
.Y(n_1694)
);

INVx4_ASAP7_75t_R g1695 ( 
.A(n_235),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_89),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_450),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1248),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_995),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1194),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1050),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1110),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_458),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1089),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_568),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_936),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_28),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_534),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1002),
.Y(n_1709)
);

CKINVDCx16_ASAP7_75t_R g1710 ( 
.A(n_1169),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1090),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1132),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1185),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1000),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_287),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_810),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_566),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1159),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_715),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1071),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_39),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_101),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_777),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_789),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_965),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_960),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_431),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_624),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_291),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1077),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1067),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_663),
.Y(n_1732)
);

CKINVDCx20_ASAP7_75t_R g1733 ( 
.A(n_622),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_802),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_118),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_612),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_927),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_371),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1246),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_773),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_300),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1053),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1249),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_675),
.Y(n_1744)
);

BUFx8_ASAP7_75t_SL g1745 ( 
.A(n_579),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_594),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_102),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_565),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_747),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1035),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_935),
.Y(n_1751)
);

BUFx5_ASAP7_75t_L g1752 ( 
.A(n_168),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1014),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_351),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1201),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_296),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_238),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_695),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_830),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_131),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_400),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_189),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1011),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_778),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_715),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_328),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_97),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_176),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1007),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1078),
.Y(n_1770)
);

BUFx10_ASAP7_75t_L g1771 ( 
.A(n_636),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_296),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1039),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_48),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_451),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_600),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_192),
.Y(n_1777)
);

CKINVDCx16_ASAP7_75t_R g1778 ( 
.A(n_958),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1098),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_29),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_100),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_506),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_957),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1073),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_940),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_206),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_402),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_249),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_801),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_996),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1237),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1168),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_944),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_260),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1010),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1009),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1049),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_206),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_199),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_104),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_4),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1233),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1087),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_916),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1022),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_478),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_741),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_159),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_134),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1076),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_844),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_205),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_986),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_460),
.Y(n_1814)
);

CKINVDCx14_ASAP7_75t_R g1815 ( 
.A(n_979),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_946),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1060),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1136),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_418),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1004),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1222),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_925),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_923),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_686),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_988),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_252),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_931),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_434),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1157),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_909),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_749),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1141),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_70),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_853),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_228),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_7),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1147),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1230),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_941),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1024),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_424),
.Y(n_1841)
);

BUFx10_ASAP7_75t_L g1842 ( 
.A(n_950),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_937),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_938),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_793),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1123),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_132),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1145),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_949),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1135),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_709),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_227),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1191),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_762),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_724),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1069),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1119),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_768),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_803),
.Y(n_1859)
);

CKINVDCx20_ASAP7_75t_R g1860 ( 
.A(n_1106),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_777),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_49),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1083),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_543),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1188),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_597),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1229),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_55),
.Y(n_1868)
);

CKINVDCx20_ASAP7_75t_R g1869 ( 
.A(n_1044),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_264),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_927),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1005),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_375),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1156),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_218),
.Y(n_1875)
);

CKINVDCx16_ASAP7_75t_R g1876 ( 
.A(n_414),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_350),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_984),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_415),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_553),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_972),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_549),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_725),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_857),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_893),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1210),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1211),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1245),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1006),
.Y(n_1889)
);

BUFx5_ASAP7_75t_L g1890 ( 
.A(n_967),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1096),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_594),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_64),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_546),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_863),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_607),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_513),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1047),
.Y(n_1898)
);

CKINVDCx20_ASAP7_75t_R g1899 ( 
.A(n_192),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_348),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1081),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_515),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_518),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_747),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_666),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_376),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1174),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_165),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_451),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_203),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1208),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_104),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_258),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_904),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1127),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1220),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_11),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_491),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1040),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_508),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_575),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1200),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_955),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_922),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_959),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_381),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1240),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_480),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1173),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_38),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_551),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_815),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_144),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_901),
.Y(n_1934)
);

BUFx10_ASAP7_75t_L g1935 ( 
.A(n_833),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1116),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1170),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1045),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_981),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_719),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_459),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1234),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1016),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_380),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1072),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_990),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_72),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1137),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_148),
.Y(n_1949)
);

CKINVDCx16_ASAP7_75t_R g1950 ( 
.A(n_585),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_60),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1121),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1150),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_609),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_315),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1128),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1094),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1182),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_452),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_150),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_853),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_302),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_1251),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_903),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_978),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_152),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1101),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_406),
.Y(n_1968)
);

INVxp67_ASAP7_75t_SL g1969 ( 
.A(n_18),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1226),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_504),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1012),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_812),
.Y(n_1973)
);

CKINVDCx14_ASAP7_75t_R g1974 ( 
.A(n_331),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_318),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1213),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_848),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1013),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_131),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_952),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1114),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_26),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1020),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1031),
.Y(n_1984)
);

CKINVDCx14_ASAP7_75t_R g1985 ( 
.A(n_1109),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_948),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_959),
.Y(n_1987)
);

INVx1_ASAP7_75t_SL g1988 ( 
.A(n_220),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_217),
.Y(n_1989)
);

INVx2_ASAP7_75t_SL g1990 ( 
.A(n_22),
.Y(n_1990)
);

INVxp67_ASAP7_75t_SL g1991 ( 
.A(n_1103),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_181),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_99),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_532),
.Y(n_1994)
);

INVx2_ASAP7_75t_SL g1995 ( 
.A(n_975),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_779),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_161),
.Y(n_1997)
);

BUFx3_ASAP7_75t_L g1998 ( 
.A(n_498),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_183),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_755),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1058),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1052),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_964),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_733),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_969),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1097),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_953),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1099),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_395),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1225),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_382),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1095),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_933),
.Y(n_2013)
);

CKINVDCx16_ASAP7_75t_R g2014 ( 
.A(n_477),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_166),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1219),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_491),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_185),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_509),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_171),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1057),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_735),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_435),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_549),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_362),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1202),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1146),
.Y(n_2027)
);

CKINVDCx14_ASAP7_75t_R g2028 ( 
.A(n_1059),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_963),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_75),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1041),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1028),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1227),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_495),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_385),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_741),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1008),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1025),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_70),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1064),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_601),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_166),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_737),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_420),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1104),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_799),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_349),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_838),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_433),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_669),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_1176),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_115),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1193),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1158),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_251),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1134),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_445),
.Y(n_2057)
);

CKINVDCx16_ASAP7_75t_R g2058 ( 
.A(n_697),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_461),
.Y(n_2059)
);

BUFx10_ASAP7_75t_L g2060 ( 
.A(n_906),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_25),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_511),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1253),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_999),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_769),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1228),
.Y(n_2066)
);

BUFx2_ASAP7_75t_L g2067 ( 
.A(n_215),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_973),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_815),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_48),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_914),
.Y(n_2071)
);

CKINVDCx20_ASAP7_75t_R g2072 ( 
.A(n_787),
.Y(n_2072)
);

INVx2_ASAP7_75t_SL g2073 ( 
.A(n_202),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1133),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_121),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_103),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_388),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_198),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1341),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1745),
.Y(n_2080)
);

INVxp67_ASAP7_75t_L g2081 ( 
.A(n_1407),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1459),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1328),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1328),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1328),
.Y(n_2085)
);

CKINVDCx16_ASAP7_75t_R g2086 ( 
.A(n_1552),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_1756),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1815),
.B(n_0),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1328),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1328),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1317),
.Y(n_2091)
);

BUFx2_ASAP7_75t_SL g2092 ( 
.A(n_1294),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1752),
.Y(n_2093)
);

CKINVDCx20_ASAP7_75t_R g2094 ( 
.A(n_1299),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1752),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1752),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1254),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1752),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1752),
.Y(n_2099)
);

INVxp67_ASAP7_75t_SL g2100 ( 
.A(n_1424),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1256),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1890),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1890),
.Y(n_2103)
);

INVx1_ASAP7_75t_SL g2104 ( 
.A(n_1808),
.Y(n_2104)
);

INVxp67_ASAP7_75t_SL g2105 ( 
.A(n_1539),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1890),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1890),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1890),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1696),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1696),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_1629),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1934),
.B(n_2067),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1280),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_1263),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1280),
.Y(n_2115)
);

BUFx2_ASAP7_75t_L g2116 ( 
.A(n_1974),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_1350),
.Y(n_2117)
);

CKINVDCx16_ASAP7_75t_R g2118 ( 
.A(n_1778),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_1262),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1280),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_1454),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1370),
.Y(n_2122)
);

INVxp33_ASAP7_75t_L g2123 ( 
.A(n_1259),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_1262),
.Y(n_2124)
);

CKINVDCx14_ASAP7_75t_R g2125 ( 
.A(n_1985),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1269),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1370),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1370),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1445),
.Y(n_2129)
);

INVxp33_ASAP7_75t_SL g2130 ( 
.A(n_1255),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1275),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1445),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1445),
.Y(n_2133)
);

INVxp33_ASAP7_75t_L g2134 ( 
.A(n_1265),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1277),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1578),
.Y(n_2136)
);

CKINVDCx16_ASAP7_75t_R g2137 ( 
.A(n_1876),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1578),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1578),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1604),
.Y(n_2140)
);

BUFx2_ASAP7_75t_L g2141 ( 
.A(n_1480),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1604),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1604),
.Y(n_2143)
);

INVx1_ASAP7_75t_SL g2144 ( 
.A(n_1367),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_1594),
.Y(n_2145)
);

CKINVDCx16_ASAP7_75t_R g2146 ( 
.A(n_1950),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_1605),
.Y(n_2147)
);

NOR2xp67_ASAP7_75t_L g2148 ( 
.A(n_1639),
.B(n_0),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1282),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1605),
.Y(n_2150)
);

CKINVDCx20_ASAP7_75t_R g2151 ( 
.A(n_1322),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_2074),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1605),
.Y(n_2153)
);

CKINVDCx20_ASAP7_75t_R g2154 ( 
.A(n_1352),
.Y(n_2154)
);

CKINVDCx20_ASAP7_75t_R g2155 ( 
.A(n_1515),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1676),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1676),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_1287),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1676),
.Y(n_2159)
);

CKINVDCx16_ASAP7_75t_R g2160 ( 
.A(n_2014),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1680),
.Y(n_2161)
);

CKINVDCx16_ASAP7_75t_R g2162 ( 
.A(n_2058),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1680),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1680),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1715),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1715),
.Y(n_2166)
);

INVx1_ASAP7_75t_SL g2167 ( 
.A(n_1381),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_1550),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1715),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1726),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1726),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1726),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1749),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1749),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1285),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1749),
.Y(n_2176)
);

INVxp33_ASAP7_75t_SL g2177 ( 
.A(n_1266),
.Y(n_2177)
);

INVxp33_ASAP7_75t_L g2178 ( 
.A(n_1278),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1268),
.Y(n_2179)
);

INVxp67_ASAP7_75t_SL g2180 ( 
.A(n_1867),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1762),
.Y(n_2181)
);

INVxp67_ASAP7_75t_SL g2182 ( 
.A(n_1485),
.Y(n_2182)
);

INVxp67_ASAP7_75t_L g2183 ( 
.A(n_1289),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1762),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1286),
.Y(n_2185)
);

INVxp33_ASAP7_75t_L g2186 ( 
.A(n_1279),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1762),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1767),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_1290),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_1601),
.B(n_2),
.Y(n_2190)
);

HB1xp67_ASAP7_75t_L g2191 ( 
.A(n_1517),
.Y(n_2191)
);

INVxp33_ASAP7_75t_L g2192 ( 
.A(n_1281),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1767),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1767),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_1457),
.Y(n_2195)
);

BUFx2_ASAP7_75t_L g2196 ( 
.A(n_1531),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1828),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1828),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1291),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1828),
.Y(n_2200)
);

HB1xp67_ASAP7_75t_L g2201 ( 
.A(n_1692),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1971),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1971),
.Y(n_2203)
);

BUFx5_ASAP7_75t_L g2204 ( 
.A(n_1258),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1971),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_1289),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_1264),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2052),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2052),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2052),
.Y(n_2210)
);

BUFx2_ASAP7_75t_L g2211 ( 
.A(n_1697),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_1300),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1799),
.Y(n_2213)
);

CKINVDCx20_ASAP7_75t_R g2214 ( 
.A(n_1860),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1908),
.Y(n_2215)
);

INVxp33_ASAP7_75t_SL g2216 ( 
.A(n_1270),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1964),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1998),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_1418),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2000),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2069),
.Y(n_2221)
);

CKINVDCx20_ASAP7_75t_R g2222 ( 
.A(n_1869),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2070),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2071),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2077),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2078),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1293),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1327),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1295),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1301),
.Y(n_2230)
);

CKINVDCx14_ASAP7_75t_R g2231 ( 
.A(n_2028),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1306),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2062),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1309),
.Y(n_2234)
);

INVxp67_ASAP7_75t_L g2235 ( 
.A(n_1292),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1310),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1313),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1318),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1329),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1327),
.Y(n_2240)
);

CKINVDCx16_ASAP7_75t_R g2241 ( 
.A(n_1710),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1330),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1336),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_1304),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1528),
.Y(n_2245)
);

INVxp67_ASAP7_75t_SL g2246 ( 
.A(n_1791),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2129),
.Y(n_2247)
);

BUFx3_ASAP7_75t_L g2248 ( 
.A(n_2152),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_L g2249 ( 
.A(n_2130),
.B(n_1261),
.Y(n_2249)
);

INVx5_ASAP7_75t_L g2250 ( 
.A(n_2213),
.Y(n_2250)
);

INVx1_ASAP7_75t_SL g2251 ( 
.A(n_2144),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_2213),
.Y(n_2252)
);

OAI22x1_ASAP7_75t_SL g2253 ( 
.A1(n_2104),
.A2(n_1450),
.B1(n_1460),
.B2(n_1297),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_2147),
.Y(n_2254)
);

INVx5_ASAP7_75t_L g2255 ( 
.A(n_2147),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_2193),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_2193),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2138),
.Y(n_2258)
);

BUFx3_ASAP7_75t_L g2259 ( 
.A(n_2207),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2143),
.Y(n_2260)
);

BUFx3_ASAP7_75t_L g2261 ( 
.A(n_2219),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_2165),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2166),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2116),
.B(n_1394),
.Y(n_2264)
);

INVx5_ASAP7_75t_L g2265 ( 
.A(n_2179),
.Y(n_2265)
);

OAI22x1_ASAP7_75t_SL g2266 ( 
.A1(n_2145),
.A2(n_1566),
.B1(n_1580),
.B2(n_1556),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_2097),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2245),
.B(n_1409),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2174),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_L g2270 ( 
.A1(n_2228),
.A2(n_1390),
.B(n_1376),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_2194),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2113),
.Y(n_2272)
);

INVx5_ASAP7_75t_L g2273 ( 
.A(n_2091),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2125),
.B(n_1463),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2179),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2101),
.B(n_1483),
.Y(n_2276)
);

INVx5_ASAP7_75t_L g2277 ( 
.A(n_2117),
.Y(n_2277)
);

BUFx8_ASAP7_75t_SL g2278 ( 
.A(n_2079),
.Y(n_2278)
);

BUFx12f_ASAP7_75t_L g2279 ( 
.A(n_2080),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2179),
.Y(n_2280)
);

CKINVDCx11_ASAP7_75t_R g2281 ( 
.A(n_2094),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2115),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_2120),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2122),
.Y(n_2284)
);

CKINVDCx8_ASAP7_75t_R g2285 ( 
.A(n_2092),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2114),
.B(n_1564),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2127),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_2126),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_2128),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_2121),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2132),
.Y(n_2291)
);

INVxp67_ASAP7_75t_L g2292 ( 
.A(n_2082),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_2133),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2136),
.Y(n_2294)
);

BUFx12f_ASAP7_75t_L g2295 ( 
.A(n_2131),
.Y(n_2295)
);

BUFx3_ASAP7_75t_L g2296 ( 
.A(n_2141),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2139),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2111),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2140),
.Y(n_2299)
);

BUFx12f_ASAP7_75t_L g2300 ( 
.A(n_2135),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2142),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2182),
.B(n_2246),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_2150),
.Y(n_2303)
);

INVxp67_ASAP7_75t_L g2304 ( 
.A(n_2196),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2088),
.B(n_2100),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2153),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2156),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2149),
.B(n_2010),
.Y(n_2308)
);

BUFx8_ASAP7_75t_L g2309 ( 
.A(n_2211),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2157),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2159),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_2161),
.Y(n_2312)
);

OA21x2_ASAP7_75t_L g2313 ( 
.A1(n_2083),
.A2(n_1326),
.B(n_1273),
.Y(n_2313)
);

HB1xp67_ASAP7_75t_L g2314 ( 
.A(n_2086),
.Y(n_2314)
);

INVx5_ASAP7_75t_L g2315 ( 
.A(n_2118),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2163),
.Y(n_2316)
);

OA21x2_ASAP7_75t_L g2317 ( 
.A1(n_2084),
.A2(n_1332),
.B(n_1331),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_2105),
.B(n_2180),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_2215),
.Y(n_2319)
);

OAI21x1_ASAP7_75t_L g2320 ( 
.A1(n_2240),
.A2(n_1395),
.B(n_1392),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2164),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2175),
.B(n_1669),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2185),
.B(n_1685),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2189),
.B(n_1773),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_2199),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2169),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2170),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_2171),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_2172),
.Y(n_2329)
);

OAI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2112),
.A2(n_1272),
.B1(n_1274),
.B2(n_1271),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2081),
.A2(n_1284),
.B1(n_1296),
.B2(n_1283),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2087),
.B(n_1476),
.Y(n_2332)
);

INVx6_ASAP7_75t_L g2333 ( 
.A(n_2137),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2212),
.B(n_1820),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_2173),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2244),
.B(n_1874),
.Y(n_2336)
);

BUFx2_ASAP7_75t_L g2337 ( 
.A(n_2146),
.Y(n_2337)
);

CKINVDCx6p67_ASAP7_75t_R g2338 ( 
.A(n_2160),
.Y(n_2338)
);

BUFx8_ASAP7_75t_SL g2339 ( 
.A(n_2151),
.Y(n_2339)
);

OAI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_2162),
.A2(n_2124),
.B1(n_2183),
.B2(n_2119),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2176),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2181),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_2184),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2187),
.Y(n_2344)
);

AND2x2_ASAP7_75t_R g2345 ( 
.A(n_2158),
.B(n_1695),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2188),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2231),
.B(n_1574),
.Y(n_2347)
);

AND2x6_ASAP7_75t_L g2348 ( 
.A(n_2190),
.B(n_1257),
.Y(n_2348)
);

OAI22x1_ASAP7_75t_SL g2349 ( 
.A1(n_2167),
.A2(n_1592),
.B1(n_1636),
.B2(n_1583),
.Y(n_2349)
);

OAI21x1_ASAP7_75t_L g2350 ( 
.A1(n_2085),
.A2(n_2027),
.B(n_1373),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2197),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_2198),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2191),
.B(n_1597),
.Y(n_2353)
);

OAI21x1_ASAP7_75t_L g2354 ( 
.A1(n_2089),
.A2(n_1378),
.B(n_1368),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2177),
.B(n_1626),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_2200),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2202),
.Y(n_2357)
);

INVx4_ASAP7_75t_L g2358 ( 
.A(n_2241),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2203),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2205),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2201),
.B(n_1654),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2208),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_2216),
.B(n_1704),
.Y(n_2363)
);

BUFx3_ASAP7_75t_L g2364 ( 
.A(n_2217),
.Y(n_2364)
);

INVx2_ASAP7_75t_SL g2365 ( 
.A(n_2218),
.Y(n_2365)
);

INVxp67_ASAP7_75t_L g2366 ( 
.A(n_2168),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2209),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2210),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2123),
.B(n_1720),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_SL g2370 ( 
.A1(n_2154),
.A2(n_1682),
.B1(n_1723),
.B2(n_1681),
.Y(n_2370)
);

BUFx8_ASAP7_75t_SL g2371 ( 
.A(n_2155),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_2220),
.Y(n_2372)
);

OAI21x1_ASAP7_75t_L g2373 ( 
.A1(n_2090),
.A2(n_1443),
.B(n_1387),
.Y(n_2373)
);

BUFx12f_ASAP7_75t_L g2374 ( 
.A(n_2195),
.Y(n_2374)
);

OAI22x1_ASAP7_75t_SL g2375 ( 
.A1(n_2214),
.A2(n_1741),
.B1(n_1744),
.B2(n_1733),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2093),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2095),
.Y(n_2377)
);

BUFx12f_ASAP7_75t_L g2378 ( 
.A(n_2206),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2096),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2098),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_2221),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2204),
.B(n_1444),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2099),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2102),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2223),
.Y(n_2385)
);

BUFx6f_ASAP7_75t_L g2386 ( 
.A(n_2224),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2235),
.B(n_1805),
.Y(n_2387)
);

BUFx8_ASAP7_75t_L g2388 ( 
.A(n_2225),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2148),
.A2(n_1302),
.B1(n_1303),
.B2(n_1298),
.Y(n_2389)
);

OAI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2134),
.A2(n_1311),
.B1(n_1312),
.B2(n_1305),
.Y(n_2390)
);

INVx5_ASAP7_75t_L g2391 ( 
.A(n_2178),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2103),
.Y(n_2392)
);

INVx6_ASAP7_75t_L g2393 ( 
.A(n_2204),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2109),
.B(n_1927),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_2222),
.Y(n_2395)
);

BUFx12f_ASAP7_75t_L g2396 ( 
.A(n_2186),
.Y(n_2396)
);

BUFx12f_ASAP7_75t_L g2397 ( 
.A(n_2192),
.Y(n_2397)
);

INVx2_ASAP7_75t_SL g2398 ( 
.A(n_2226),
.Y(n_2398)
);

AOI22x1_ASAP7_75t_SL g2399 ( 
.A1(n_2227),
.A2(n_1899),
.B1(n_1906),
.B2(n_1747),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_2229),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2110),
.B(n_1958),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2106),
.Y(n_2402)
);

BUFx6f_ASAP7_75t_L g2403 ( 
.A(n_2230),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2232),
.A2(n_2037),
.B1(n_1969),
.B2(n_1320),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2233),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2204),
.B(n_2107),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2108),
.Y(n_2407)
);

OAI21x1_ASAP7_75t_L g2408 ( 
.A1(n_2234),
.A2(n_1461),
.B(n_1458),
.Y(n_2408)
);

BUFx8_ASAP7_75t_SL g2409 ( 
.A(n_2236),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_SL g2410 ( 
.A1(n_2237),
.A2(n_1925),
.B1(n_2072),
.B2(n_1913),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2238),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2239),
.Y(n_2412)
);

AOI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2242),
.A2(n_1321),
.B1(n_1323),
.B2(n_1316),
.Y(n_2413)
);

CKINVDCx6p67_ASAP7_75t_R g2414 ( 
.A(n_2204),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2243),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2097),
.B(n_1468),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_2152),
.Y(n_2417)
);

BUFx3_ASAP7_75t_L g2418 ( 
.A(n_2152),
.Y(n_2418)
);

INVx4_ASAP7_75t_L g2419 ( 
.A(n_2097),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2129),
.Y(n_2420)
);

HB1xp67_ASAP7_75t_L g2421 ( 
.A(n_2082),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_2147),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2116),
.B(n_2051),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2082),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2147),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2116),
.B(n_1610),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_2147),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2147),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2147),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_2147),
.Y(n_2430)
);

BUFx3_ASAP7_75t_L g2431 ( 
.A(n_2152),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2129),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2116),
.B(n_1991),
.Y(n_2433)
);

OAI22x1_ASAP7_75t_SL g2434 ( 
.A1(n_2104),
.A2(n_2076),
.B1(n_1325),
.B2(n_1333),
.Y(n_2434)
);

INVx5_ASAP7_75t_L g2435 ( 
.A(n_2213),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2147),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2147),
.Y(n_2437)
);

INVx3_ASAP7_75t_L g2438 ( 
.A(n_2213),
.Y(n_2438)
);

BUFx6f_ASAP7_75t_L g2439 ( 
.A(n_2147),
.Y(n_2439)
);

BUFx8_ASAP7_75t_SL g2440 ( 
.A(n_2079),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_2097),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2082),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2116),
.B(n_1611),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2152),
.Y(n_2444)
);

BUFx12f_ASAP7_75t_L g2445 ( 
.A(n_2079),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2104),
.A2(n_1342),
.B1(n_1343),
.B2(n_1324),
.Y(n_2446)
);

INVx4_ASAP7_75t_L g2447 ( 
.A(n_2097),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_2152),
.Y(n_2448)
);

AND2x6_ASAP7_75t_L g2449 ( 
.A(n_2088),
.B(n_1260),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2129),
.Y(n_2450)
);

HB1xp67_ASAP7_75t_L g2451 ( 
.A(n_2082),
.Y(n_2451)
);

BUFx3_ASAP7_75t_L g2452 ( 
.A(n_2152),
.Y(n_2452)
);

INVx3_ASAP7_75t_L g2453 ( 
.A(n_2213),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2147),
.Y(n_2454)
);

INVx4_ASAP7_75t_L g2455 ( 
.A(n_2097),
.Y(n_2455)
);

AOI22xp5_ASAP7_75t_L g2456 ( 
.A1(n_2104),
.A2(n_1348),
.B1(n_1349),
.B2(n_1347),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2129),
.Y(n_2457)
);

OAI21x1_ASAP7_75t_L g2458 ( 
.A1(n_2228),
.A2(n_1492),
.B(n_1477),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2097),
.B(n_1498),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2116),
.B(n_1612),
.Y(n_2460)
);

BUFx8_ASAP7_75t_L g2461 ( 
.A(n_2116),
.Y(n_2461)
);

BUFx12f_ASAP7_75t_L g2462 ( 
.A(n_2079),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2147),
.Y(n_2463)
);

OAI22x1_ASAP7_75t_R g2464 ( 
.A1(n_2094),
.A2(n_1356),
.B1(n_1358),
.B2(n_1353),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2129),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_2082),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2147),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2116),
.B(n_1631),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2097),
.Y(n_2469)
);

INVx5_ASAP7_75t_L g2470 ( 
.A(n_2213),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2129),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2097),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_2116),
.B(n_1504),
.Y(n_2473)
);

OA21x2_ASAP7_75t_L g2474 ( 
.A1(n_2083),
.A2(n_1567),
.B(n_1536),
.Y(n_2474)
);

INVxp67_ASAP7_75t_L g2475 ( 
.A(n_2082),
.Y(n_2475)
);

BUFx12f_ASAP7_75t_L g2476 ( 
.A(n_2079),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_2152),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2097),
.B(n_1569),
.Y(n_2478)
);

INVx6_ASAP7_75t_L g2479 ( 
.A(n_2213),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_2082),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2241),
.B(n_1292),
.Y(n_2481)
);

OAI21x1_ASAP7_75t_L g2482 ( 
.A1(n_2228),
.A2(n_1579),
.B(n_1573),
.Y(n_2482)
);

INVx5_ASAP7_75t_L g2483 ( 
.A(n_2213),
.Y(n_2483)
);

BUFx6f_ASAP7_75t_L g2484 ( 
.A(n_2147),
.Y(n_2484)
);

AOI22x1_ASAP7_75t_SL g2485 ( 
.A1(n_2094),
.A2(n_1360),
.B1(n_1363),
.B2(n_1359),
.Y(n_2485)
);

INVx2_ASAP7_75t_SL g2486 ( 
.A(n_2117),
.Y(n_2486)
);

INVx3_ASAP7_75t_L g2487 ( 
.A(n_2213),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2082),
.Y(n_2488)
);

INVx2_ASAP7_75t_SL g2489 ( 
.A(n_2117),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2147),
.Y(n_2490)
);

BUFx12f_ASAP7_75t_L g2491 ( 
.A(n_2079),
.Y(n_2491)
);

OA21x2_ASAP7_75t_L g2492 ( 
.A1(n_2083),
.A2(n_1644),
.B(n_1619),
.Y(n_2492)
);

INVx2_ASAP7_75t_SL g2493 ( 
.A(n_2117),
.Y(n_2493)
);

OA21x2_ASAP7_75t_L g2494 ( 
.A1(n_2083),
.A2(n_1660),
.B(n_1645),
.Y(n_2494)
);

INVx3_ASAP7_75t_L g2495 ( 
.A(n_2213),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2147),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_2147),
.Y(n_2497)
);

BUFx2_ASAP7_75t_L g2498 ( 
.A(n_2082),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2116),
.B(n_1679),
.Y(n_2499)
);

INVx3_ASAP7_75t_L g2500 ( 
.A(n_2213),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2147),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2129),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2129),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2097),
.B(n_1709),
.Y(n_2504)
);

BUFx8_ASAP7_75t_SL g2505 ( 
.A(n_2079),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2097),
.B(n_1713),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2082),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2129),
.Y(n_2508)
);

INVx5_ASAP7_75t_L g2509 ( 
.A(n_2213),
.Y(n_2509)
);

OAI22x1_ASAP7_75t_L g2510 ( 
.A1(n_2104),
.A2(n_1288),
.B1(n_1339),
.B2(n_1308),
.Y(n_2510)
);

INVx5_ASAP7_75t_L g2511 ( 
.A(n_2213),
.Y(n_2511)
);

INVx4_ASAP7_75t_L g2512 ( 
.A(n_2097),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2147),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2147),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2116),
.B(n_1732),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_2147),
.Y(n_2516)
);

BUFx3_ASAP7_75t_L g2517 ( 
.A(n_2152),
.Y(n_2517)
);

INVx3_ASAP7_75t_L g2518 ( 
.A(n_2213),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2104),
.A2(n_1365),
.B1(n_1374),
.B2(n_1364),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2147),
.Y(n_2520)
);

INVx5_ASAP7_75t_L g2521 ( 
.A(n_2213),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2129),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2129),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2152),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_2147),
.Y(n_2525)
);

BUFx8_ASAP7_75t_L g2526 ( 
.A(n_2116),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2147),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2147),
.Y(n_2528)
);

INVx2_ASAP7_75t_SL g2529 ( 
.A(n_2117),
.Y(n_2529)
);

INVx5_ASAP7_75t_L g2530 ( 
.A(n_2213),
.Y(n_2530)
);

AOI22xp5_ASAP7_75t_L g2531 ( 
.A1(n_2104),
.A2(n_1380),
.B1(n_1386),
.B2(n_1375),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2147),
.Y(n_2532)
);

OAI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2104),
.A2(n_1396),
.B1(n_1397),
.B2(n_1388),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2147),
.Y(n_2534)
);

BUFx3_ASAP7_75t_L g2535 ( 
.A(n_2152),
.Y(n_2535)
);

HB1xp67_ASAP7_75t_L g2536 ( 
.A(n_2082),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2147),
.Y(n_2537)
);

CKINVDCx20_ASAP7_75t_R g2538 ( 
.A(n_2094),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_2116),
.B(n_1731),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2147),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2147),
.Y(n_2541)
);

INVx5_ASAP7_75t_L g2542 ( 
.A(n_2213),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2129),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2147),
.Y(n_2544)
);

OA21x2_ASAP7_75t_L g2545 ( 
.A1(n_2083),
.A2(n_1750),
.B(n_1743),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2129),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2129),
.Y(n_2547)
);

BUFx6f_ASAP7_75t_L g2548 ( 
.A(n_2147),
.Y(n_2548)
);

BUFx2_ASAP7_75t_L g2549 ( 
.A(n_2082),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2147),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2129),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2129),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2129),
.Y(n_2553)
);

BUFx6f_ASAP7_75t_L g2554 ( 
.A(n_2147),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2130),
.B(n_1755),
.Y(n_2555)
);

BUFx8_ASAP7_75t_L g2556 ( 
.A(n_2116),
.Y(n_2556)
);

CKINVDCx16_ASAP7_75t_R g2557 ( 
.A(n_2086),
.Y(n_2557)
);

BUFx6f_ASAP7_75t_L g2558 ( 
.A(n_2147),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2097),
.B(n_1763),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2097),
.B(n_1784),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2147),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2147),
.Y(n_2562)
);

BUFx6f_ASAP7_75t_L g2563 ( 
.A(n_2147),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2116),
.B(n_1990),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2129),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2129),
.Y(n_2566)
);

AND2x4_ASAP7_75t_L g2567 ( 
.A(n_2116),
.B(n_1795),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2147),
.Y(n_2568)
);

OAI21x1_ASAP7_75t_L g2569 ( 
.A1(n_2228),
.A2(n_1813),
.B(n_1802),
.Y(n_2569)
);

AOI22x1_ASAP7_75t_SL g2570 ( 
.A1(n_2094),
.A2(n_1402),
.B1(n_1403),
.B2(n_1398),
.Y(n_2570)
);

BUFx3_ASAP7_75t_L g2571 ( 
.A(n_2152),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2147),
.Y(n_2572)
);

CKINVDCx20_ASAP7_75t_R g2573 ( 
.A(n_2094),
.Y(n_2573)
);

BUFx12f_ASAP7_75t_L g2574 ( 
.A(n_2079),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2369),
.B(n_1346),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2339),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2411),
.Y(n_2577)
);

NOR2x1_ASAP7_75t_L g2578 ( 
.A(n_2248),
.B(n_1825),
.Y(n_2578)
);

BUFx6f_ASAP7_75t_L g2579 ( 
.A(n_2254),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2275),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2280),
.Y(n_2581)
);

BUFx6f_ASAP7_75t_L g2582 ( 
.A(n_2256),
.Y(n_2582)
);

AND2x4_ASAP7_75t_L g2583 ( 
.A(n_2290),
.B(n_1995),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2412),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2296),
.B(n_1997),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2414),
.B(n_1307),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2386),
.Y(n_2587)
);

INVx3_ASAP7_75t_L g2588 ( 
.A(n_2479),
.Y(n_2588)
);

HB1xp67_ASAP7_75t_L g2589 ( 
.A(n_2391),
.Y(n_2589)
);

BUFx6f_ASAP7_75t_L g2590 ( 
.A(n_2422),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2425),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2400),
.Y(n_2592)
);

HB1xp67_ASAP7_75t_L g2593 ( 
.A(n_2251),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2263),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2271),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2322),
.B(n_2073),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2403),
.Y(n_2597)
);

BUFx3_ASAP7_75t_L g2598 ( 
.A(n_2259),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2405),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2379),
.Y(n_2600)
);

BUFx2_ASAP7_75t_L g2601 ( 
.A(n_2396),
.Y(n_2601)
);

INVxp67_ASAP7_75t_L g2602 ( 
.A(n_2249),
.Y(n_2602)
);

BUFx6f_ASAP7_75t_L g2603 ( 
.A(n_2427),
.Y(n_2603)
);

OR2x6_ASAP7_75t_L g2604 ( 
.A(n_2333),
.B(n_1276),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2247),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2323),
.B(n_1410),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2264),
.B(n_1346),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2392),
.Y(n_2608)
);

AND2x4_ASAP7_75t_L g2609 ( 
.A(n_2261),
.B(n_1337),
.Y(n_2609)
);

BUFx2_ASAP7_75t_L g2610 ( 
.A(n_2397),
.Y(n_2610)
);

OA21x2_ASAP7_75t_L g2611 ( 
.A1(n_2270),
.A2(n_1832),
.B(n_1829),
.Y(n_2611)
);

BUFx3_ASAP7_75t_L g2612 ( 
.A(n_2417),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2423),
.B(n_1391),
.Y(n_2613)
);

BUFx6f_ASAP7_75t_L g2614 ( 
.A(n_2430),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2376),
.Y(n_2615)
);

BUFx8_ASAP7_75t_L g2616 ( 
.A(n_2337),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2377),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2380),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2324),
.B(n_1411),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2383),
.Y(n_2620)
);

NAND2xp33_ASAP7_75t_SL g2621 ( 
.A(n_2486),
.B(n_1412),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2258),
.Y(n_2622)
);

BUFx3_ASAP7_75t_L g2623 ( 
.A(n_2418),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2384),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2371),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2402),
.Y(n_2626)
);

OA21x2_ASAP7_75t_L g2627 ( 
.A1(n_2320),
.A2(n_1853),
.B(n_1840),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2407),
.Y(n_2628)
);

CKINVDCx6p67_ASAP7_75t_R g2629 ( 
.A(n_2315),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2366),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2319),
.Y(n_2631)
);

BUFx6f_ASAP7_75t_L g2632 ( 
.A(n_2436),
.Y(n_2632)
);

INVx4_ASAP7_75t_L g2633 ( 
.A(n_2295),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2364),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2260),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2420),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_2437),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2334),
.B(n_1416),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2415),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2489),
.B(n_1391),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2432),
.Y(n_2641)
);

CKINVDCx9p33_ASAP7_75t_R g2642 ( 
.A(n_2399),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2431),
.B(n_1344),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2493),
.B(n_1435),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2450),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2457),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2529),
.B(n_1435),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2465),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2398),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2381),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2385),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2272),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2471),
.Y(n_2653)
);

BUFx3_ASAP7_75t_L g2654 ( 
.A(n_2444),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2287),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2306),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2336),
.B(n_1314),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2353),
.B(n_1524),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2416),
.B(n_1315),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2502),
.Y(n_2660)
);

AND2x2_ASAP7_75t_SL g2661 ( 
.A(n_2557),
.B(n_1267),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2439),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2307),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2311),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2321),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2503),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2448),
.Y(n_2667)
);

AND2x4_ASAP7_75t_L g2668 ( 
.A(n_2452),
.B(n_2477),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2508),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2361),
.B(n_1524),
.Y(n_2670)
);

AND2x6_ASAP7_75t_L g2671 ( 
.A(n_2426),
.B(n_1448),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2463),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2327),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2355),
.B(n_2363),
.Y(n_2674)
);

BUFx6f_ASAP7_75t_L g2675 ( 
.A(n_2467),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2459),
.B(n_2478),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2342),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2346),
.Y(n_2678)
);

AND2x6_ASAP7_75t_L g2679 ( 
.A(n_2443),
.B(n_1466),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2357),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2360),
.Y(n_2681)
);

OAI22xp5_ASAP7_75t_SL g2682 ( 
.A1(n_2410),
.A2(n_1520),
.B1(n_1521),
.B2(n_1489),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2368),
.Y(n_2683)
);

AND2x4_ASAP7_75t_L g2684 ( 
.A(n_2517),
.B(n_1351),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2522),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2504),
.B(n_1423),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2523),
.Y(n_2687)
);

BUFx6f_ASAP7_75t_L g2688 ( 
.A(n_2484),
.Y(n_2688)
);

BUFx2_ASAP7_75t_L g2689 ( 
.A(n_2374),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2274),
.B(n_1577),
.Y(n_2690)
);

BUFx6f_ASAP7_75t_L g2691 ( 
.A(n_2496),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2524),
.B(n_1354),
.Y(n_2692)
);

BUFx2_ASAP7_75t_L g2693 ( 
.A(n_2314),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2543),
.Y(n_2694)
);

BUFx2_ASAP7_75t_L g2695 ( 
.A(n_2424),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2546),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2547),
.Y(n_2697)
);

INVxp33_ASAP7_75t_L g2698 ( 
.A(n_2298),
.Y(n_2698)
);

CKINVDCx5p33_ASAP7_75t_R g2699 ( 
.A(n_2267),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2347),
.B(n_1577),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2332),
.B(n_1606),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2551),
.Y(n_2702)
);

INVx3_ASAP7_75t_L g2703 ( 
.A(n_2497),
.Y(n_2703)
);

BUFx6f_ASAP7_75t_L g2704 ( 
.A(n_2501),
.Y(n_2704)
);

AND2x6_ASAP7_75t_L g2705 ( 
.A(n_2460),
.B(n_1621),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2552),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2553),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2506),
.B(n_1338),
.Y(n_2708)
);

BUFx2_ASAP7_75t_L g2709 ( 
.A(n_2480),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2565),
.Y(n_2710)
);

AOI22x1_ASAP7_75t_SL g2711 ( 
.A1(n_2538),
.A2(n_1428),
.B1(n_1431),
.B2(n_1427),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2566),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2516),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2559),
.B(n_1340),
.Y(n_2714)
);

OAI22xp5_ASAP7_75t_SL g2715 ( 
.A1(n_2404),
.A2(n_1650),
.B1(n_1661),
.B2(n_1623),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2428),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2282),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2291),
.Y(n_2718)
);

OR2x6_ASAP7_75t_L g2719 ( 
.A(n_2395),
.B(n_1472),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_2288),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2325),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2560),
.B(n_1345),
.Y(n_2722)
);

INVx4_ASAP7_75t_L g2723 ( 
.A(n_2300),
.Y(n_2723)
);

NOR2xp33_ASAP7_75t_L g2724 ( 
.A(n_2276),
.B(n_1433),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2268),
.B(n_1606),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2294),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_L g2727 ( 
.A(n_2520),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2429),
.Y(n_2728)
);

BUFx2_ASAP7_75t_L g2729 ( 
.A(n_2498),
.Y(n_2729)
);

HB1xp67_ASAP7_75t_L g2730 ( 
.A(n_2304),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2305),
.B(n_1355),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_2535),
.B(n_1362),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2525),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2297),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2454),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2527),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2490),
.Y(n_2737)
);

OAI21x1_ASAP7_75t_L g2738 ( 
.A1(n_2354),
.A2(n_2373),
.B(n_2350),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2555),
.B(n_1361),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2299),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2513),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2532),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2544),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2514),
.Y(n_2744)
);

BUFx6f_ASAP7_75t_L g2745 ( 
.A(n_2548),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2301),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2528),
.Y(n_2747)
);

BUFx6f_ASAP7_75t_L g2748 ( 
.A(n_2554),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2310),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2316),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2534),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_L g2752 ( 
.A(n_2286),
.B(n_1437),
.Y(n_2752)
);

BUFx8_ASAP7_75t_L g2753 ( 
.A(n_2549),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2341),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2351),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_2441),
.Y(n_2756)
);

OA21x2_ASAP7_75t_L g2757 ( 
.A1(n_2408),
.A2(n_1889),
.B(n_1878),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2537),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2359),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2468),
.B(n_2515),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2540),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2308),
.B(n_1366),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2362),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2558),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2541),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2387),
.B(n_1369),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_SL g2767 ( 
.A(n_2285),
.B(n_1717),
.Y(n_2767)
);

INVx6_ASAP7_75t_L g2768 ( 
.A(n_2309),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2550),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2318),
.B(n_1371),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2302),
.B(n_1372),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2564),
.B(n_1618),
.Y(n_2772)
);

BUFx3_ASAP7_75t_L g2773 ( 
.A(n_2571),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2568),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2367),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2572),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2561),
.Y(n_2777)
);

AOI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2348),
.A2(n_1761),
.B1(n_1788),
.B2(n_1725),
.Y(n_2778)
);

CKINVDCx8_ASAP7_75t_R g2779 ( 
.A(n_2449),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2262),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2283),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2365),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2284),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2289),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2562),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2433),
.B(n_1379),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_L g2787 ( 
.A(n_2563),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2393),
.B(n_2406),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2293),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2421),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2442),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2303),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2372),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2394),
.B(n_1383),
.Y(n_2794)
);

HB1xp67_ASAP7_75t_L g2795 ( 
.A(n_2451),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2312),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2344),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2326),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2458),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2401),
.B(n_1401),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2328),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2329),
.Y(n_2802)
);

AND2x2_ASAP7_75t_SL g2803 ( 
.A(n_2358),
.B(n_1319),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2482),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2277),
.B(n_1618),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2569),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2466),
.Y(n_2807)
);

BUFx6f_ASAP7_75t_L g2808 ( 
.A(n_2335),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2257),
.Y(n_2809)
);

INVx2_ASAP7_75t_SL g2810 ( 
.A(n_2488),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2343),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2352),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2356),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_2507),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2382),
.B(n_2473),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2269),
.Y(n_2816)
);

AND2x4_ASAP7_75t_SL g2817 ( 
.A(n_2338),
.B(n_1771),
.Y(n_2817)
);

AND2x4_ASAP7_75t_L g2818 ( 
.A(n_2499),
.B(n_1377),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2536),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2252),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2438),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2453),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2487),
.Y(n_2823)
);

BUFx3_ASAP7_75t_L g2824 ( 
.A(n_2250),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_L g2825 ( 
.A(n_2419),
.B(n_1438),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2495),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2446),
.B(n_1771),
.Y(n_2827)
);

INVx1_ASAP7_75t_SL g2828 ( 
.A(n_2573),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2292),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2500),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2518),
.Y(n_2831)
);

HB1xp67_ASAP7_75t_L g2832 ( 
.A(n_2475),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2313),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2317),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2474),
.Y(n_2835)
);

INVx3_ASAP7_75t_L g2836 ( 
.A(n_2265),
.Y(n_2836)
);

BUFx6f_ASAP7_75t_L g2837 ( 
.A(n_2265),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2447),
.B(n_1441),
.Y(n_2838)
);

NAND2xp33_ASAP7_75t_R g2839 ( 
.A(n_2469),
.B(n_1442),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2492),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2494),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2255),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2545),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2255),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2539),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2456),
.B(n_1842),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2567),
.Y(n_2847)
);

INVx3_ASAP7_75t_L g2848 ( 
.A(n_2435),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2531),
.B(n_1842),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2273),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2470),
.Y(n_2851)
);

NAND2xp33_ASAP7_75t_L g2852 ( 
.A(n_2449),
.B(n_1268),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2455),
.B(n_1404),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2483),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2509),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2472),
.B(n_1408),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2511),
.Y(n_2857)
);

BUFx6f_ASAP7_75t_L g2858 ( 
.A(n_2521),
.Y(n_2858)
);

INVx3_ASAP7_75t_L g2859 ( 
.A(n_2530),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2512),
.B(n_1446),
.Y(n_2860)
);

INVx3_ASAP7_75t_L g2861 ( 
.A(n_2542),
.Y(n_2861)
);

NAND2xp33_ASAP7_75t_R g2862 ( 
.A(n_2485),
.B(n_1447),
.Y(n_2862)
);

CKINVDCx16_ASAP7_75t_R g2863 ( 
.A(n_2464),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2413),
.Y(n_2864)
);

OA21x2_ASAP7_75t_L g2865 ( 
.A1(n_2389),
.A2(n_1911),
.B(n_1907),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2390),
.Y(n_2866)
);

INVx2_ASAP7_75t_SL g2867 ( 
.A(n_2481),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2519),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2533),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2331),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2348),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2330),
.B(n_1413),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2510),
.Y(n_2873)
);

INVx3_ASAP7_75t_L g2874 ( 
.A(n_2409),
.Y(n_2874)
);

BUFx8_ASAP7_75t_L g2875 ( 
.A(n_2279),
.Y(n_2875)
);

BUFx2_ASAP7_75t_L g2876 ( 
.A(n_2461),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2340),
.B(n_1414),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2370),
.B(n_1935),
.Y(n_2878)
);

CKINVDCx5p33_ASAP7_75t_R g2879 ( 
.A(n_2281),
.Y(n_2879)
);

BUFx8_ASAP7_75t_L g2880 ( 
.A(n_2574),
.Y(n_2880)
);

AND2x4_ASAP7_75t_L g2881 ( 
.A(n_2345),
.B(n_1382),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2378),
.B(n_1935),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2388),
.Y(n_2883)
);

NOR2x1_ASAP7_75t_L g2884 ( 
.A(n_2434),
.B(n_1915),
.Y(n_2884)
);

INVx3_ASAP7_75t_L g2885 ( 
.A(n_2526),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2556),
.B(n_1425),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2570),
.Y(n_2887)
);

INVxp67_ASAP7_75t_L g2888 ( 
.A(n_2253),
.Y(n_2888)
);

BUFx6f_ASAP7_75t_L g2889 ( 
.A(n_2579),
.Y(n_2889)
);

OAI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2674),
.A2(n_1812),
.B1(n_1988),
.B2(n_1794),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2760),
.B(n_1430),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2579),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2605),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2577),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2584),
.Y(n_2895)
);

BUFx2_ASAP7_75t_L g2896 ( 
.A(n_2593),
.Y(n_2896)
);

BUFx6f_ASAP7_75t_L g2897 ( 
.A(n_2582),
.Y(n_2897)
);

INVx5_ASAP7_75t_L g2898 ( 
.A(n_2858),
.Y(n_2898)
);

BUFx10_ASAP7_75t_L g2899 ( 
.A(n_2576),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2652),
.Y(n_2900)
);

INVx3_ASAP7_75t_L g2901 ( 
.A(n_2582),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2622),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2575),
.B(n_2060),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2676),
.B(n_1942),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2635),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2636),
.Y(n_2906)
);

INVx4_ASAP7_75t_L g2907 ( 
.A(n_2858),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2686),
.B(n_1948),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2641),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2645),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2646),
.Y(n_2911)
);

INVx1_ASAP7_75t_SL g2912 ( 
.A(n_2630),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2607),
.B(n_2060),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2590),
.Y(n_2914)
);

BUFx6f_ASAP7_75t_L g2915 ( 
.A(n_2590),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2655),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2648),
.Y(n_2917)
);

INVxp67_ASAP7_75t_L g2918 ( 
.A(n_2613),
.Y(n_2918)
);

BUFx2_ASAP7_75t_L g2919 ( 
.A(n_2695),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2653),
.Y(n_2920)
);

OR2x6_ASAP7_75t_L g2921 ( 
.A(n_2768),
.B(n_2445),
.Y(n_2921)
);

AND3x2_ASAP7_75t_L g2922 ( 
.A(n_2689),
.B(n_1335),
.C(n_1334),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2656),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2660),
.Y(n_2924)
);

AOI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2866),
.A2(n_1449),
.B1(n_1451),
.B2(n_1432),
.Y(n_2925)
);

INVx3_ASAP7_75t_L g2926 ( 
.A(n_2603),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2602),
.B(n_2462),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2663),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2606),
.B(n_1970),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2699),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2664),
.Y(n_2931)
);

INVx3_ASAP7_75t_L g2932 ( 
.A(n_2603),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2666),
.Y(n_2933)
);

INVx1_ASAP7_75t_SL g2934 ( 
.A(n_2709),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2619),
.B(n_2638),
.Y(n_2935)
);

BUFx3_ASAP7_75t_L g2936 ( 
.A(n_2598),
.Y(n_2936)
);

INVx8_ASAP7_75t_L g2937 ( 
.A(n_2604),
.Y(n_2937)
);

BUFx3_ASAP7_75t_L g2938 ( 
.A(n_2612),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2669),
.Y(n_2939)
);

NOR2xp33_ASAP7_75t_L g2940 ( 
.A(n_2739),
.B(n_2266),
.Y(n_2940)
);

INVx2_ASAP7_75t_SL g2941 ( 
.A(n_2729),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2665),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2673),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2677),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2596),
.B(n_1976),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2678),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2685),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2680),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2767),
.B(n_1467),
.Y(n_2949)
);

AOI22xp5_ASAP7_75t_L g2950 ( 
.A1(n_2868),
.A2(n_1470),
.B1(n_1473),
.B2(n_1469),
.Y(n_2950)
);

INVxp33_ASAP7_75t_L g2951 ( 
.A(n_2790),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2681),
.Y(n_2952)
);

OR2x6_ASAP7_75t_L g2953 ( 
.A(n_2876),
.B(n_2476),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2725),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2683),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2702),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2724),
.B(n_1478),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2752),
.B(n_1983),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2706),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2717),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2687),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2718),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2698),
.B(n_2349),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2614),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2772),
.B(n_2491),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2694),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2815),
.B(n_2002),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2726),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2734),
.Y(n_2969)
);

INVx5_ASAP7_75t_L g2970 ( 
.A(n_2842),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2740),
.Y(n_2971)
);

AND2x6_ASAP7_75t_L g2972 ( 
.A(n_2833),
.B(n_2016),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2690),
.B(n_1453),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2746),
.Y(n_2974)
);

BUFx10_ASAP7_75t_L g2975 ( 
.A(n_2625),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2788),
.B(n_2032),
.Y(n_2976)
);

BUFx3_ASAP7_75t_L g2977 ( 
.A(n_2623),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2696),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2614),
.Y(n_2979)
);

AOI22xp33_ASAP7_75t_L g2980 ( 
.A1(n_2834),
.A2(n_2835),
.B1(n_2841),
.B2(n_2840),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2749),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2697),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_SL g2983 ( 
.A(n_2700),
.B(n_1479),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2750),
.Y(n_2984)
);

CKINVDCx5p33_ASAP7_75t_R g2985 ( 
.A(n_2720),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2707),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2754),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2710),
.Y(n_2988)
);

CKINVDCx5p33_ASAP7_75t_R g2989 ( 
.A(n_2721),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2659),
.B(n_2040),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2632),
.Y(n_2991)
);

AND2x2_ASAP7_75t_SL g2992 ( 
.A(n_2863),
.B(n_2375),
.Y(n_2992)
);

INVx1_ASAP7_75t_SL g2993 ( 
.A(n_2693),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2755),
.Y(n_2994)
);

INVx2_ASAP7_75t_SL g2995 ( 
.A(n_2583),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_R g2996 ( 
.A(n_2879),
.B(n_1487),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2819),
.B(n_2278),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2759),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2763),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2658),
.B(n_1455),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2712),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2803),
.B(n_1491),
.Y(n_3002)
);

AOI22xp33_ASAP7_75t_L g3003 ( 
.A1(n_2843),
.A2(n_2064),
.B1(n_2056),
.B2(n_1327),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2600),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2708),
.B(n_1496),
.Y(n_3005)
);

INVx4_ASAP7_75t_L g3006 ( 
.A(n_2789),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2670),
.B(n_1456),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2701),
.B(n_2640),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2775),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2608),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2639),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2816),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2644),
.B(n_1462),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2615),
.Y(n_3014)
);

NAND2xp33_ASAP7_75t_L g3015 ( 
.A(n_2714),
.B(n_1518),
.Y(n_3015)
);

CKINVDCx5p33_ASAP7_75t_R g3016 ( 
.A(n_2756),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2722),
.B(n_1529),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2617),
.Y(n_3018)
);

BUFx6f_ASAP7_75t_L g3019 ( 
.A(n_2632),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_SL g3020 ( 
.A(n_2864),
.B(n_1538),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2780),
.Y(n_3021)
);

INVx2_ASAP7_75t_SL g3022 ( 
.A(n_2585),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2618),
.Y(n_3023)
);

OR2x6_ASAP7_75t_L g3024 ( 
.A(n_2883),
.B(n_2633),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2580),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2581),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2620),
.Y(n_3027)
);

INVx2_ASAP7_75t_SL g3028 ( 
.A(n_2791),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2624),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2626),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_2839),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2628),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_SL g3033 ( 
.A(n_2825),
.B(n_1542),
.Y(n_3033)
);

INVx1_ASAP7_75t_SL g3034 ( 
.A(n_2795),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2716),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2728),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2735),
.Y(n_3037)
);

INVx2_ASAP7_75t_SL g3038 ( 
.A(n_2807),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2737),
.Y(n_3039)
);

INVxp67_ASAP7_75t_L g3040 ( 
.A(n_2647),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2650),
.Y(n_3041)
);

INVx2_ASAP7_75t_SL g3042 ( 
.A(n_2814),
.Y(n_3042)
);

AND2x4_ASAP7_75t_L g3043 ( 
.A(n_2668),
.B(n_1389),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_2629),
.Y(n_3044)
);

CKINVDCx5p33_ASAP7_75t_R g3045 ( 
.A(n_2828),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2829),
.B(n_2440),
.Y(n_3046)
);

BUFx2_ASAP7_75t_L g3047 ( 
.A(n_2671),
.Y(n_3047)
);

BUFx10_ASAP7_75t_L g3048 ( 
.A(n_2817),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2805),
.B(n_1474),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2869),
.A2(n_1327),
.B1(n_1385),
.B2(n_1357),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2741),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2744),
.Y(n_3052)
);

BUFx4f_ASAP7_75t_L g3053 ( 
.A(n_2871),
.Y(n_3053)
);

INVx4_ASAP7_75t_L g3054 ( 
.A(n_2789),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2651),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2747),
.Y(n_3056)
);

INVx2_ASAP7_75t_SL g3057 ( 
.A(n_2810),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2832),
.B(n_1475),
.Y(n_3058)
);

INVx3_ASAP7_75t_L g3059 ( 
.A(n_2672),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2657),
.B(n_2505),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2751),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2762),
.B(n_1551),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2758),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2761),
.Y(n_3064)
);

BUFx6f_ASAP7_75t_SL g3065 ( 
.A(n_2723),
.Y(n_3065)
);

CKINVDCx16_ASAP7_75t_R g3066 ( 
.A(n_2719),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_SL g3067 ( 
.A(n_2838),
.B(n_1557),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2765),
.Y(n_3068)
);

BUFx6f_ASAP7_75t_L g3069 ( 
.A(n_2672),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2769),
.Y(n_3070)
);

CKINVDCx5p33_ASAP7_75t_R g3071 ( 
.A(n_2875),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2774),
.Y(n_3072)
);

AOI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2799),
.A2(n_1399),
.B(n_1393),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2776),
.Y(n_3074)
);

INVxp67_ASAP7_75t_SL g3075 ( 
.A(n_2793),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2860),
.B(n_1565),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2809),
.Y(n_3077)
);

INVx8_ASAP7_75t_L g3078 ( 
.A(n_2671),
.Y(n_3078)
);

INVx2_ASAP7_75t_SL g3079 ( 
.A(n_2609),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2770),
.B(n_1571),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_2880),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2796),
.Y(n_3082)
);

CKINVDCx5p33_ASAP7_75t_R g3083 ( 
.A(n_2616),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2872),
.B(n_1587),
.Y(n_3084)
);

INVx2_ASAP7_75t_SL g3085 ( 
.A(n_2643),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2797),
.Y(n_3086)
);

INVx2_ASAP7_75t_SL g3087 ( 
.A(n_2684),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2661),
.B(n_1482),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2870),
.B(n_1493),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2820),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2586),
.B(n_1591),
.Y(n_3091)
);

INVx4_ASAP7_75t_L g3092 ( 
.A(n_2808),
.Y(n_3092)
);

NAND3xp33_ASAP7_75t_L g3093 ( 
.A(n_2852),
.B(n_1495),
.C(n_1494),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2821),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2822),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2823),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2826),
.Y(n_3097)
);

BUFx3_ASAP7_75t_L g3098 ( 
.A(n_2654),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2830),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2831),
.Y(n_3100)
);

INVx5_ASAP7_75t_L g3101 ( 
.A(n_2842),
.Y(n_3101)
);

NAND2xp33_ASAP7_75t_L g3102 ( 
.A(n_2871),
.B(n_2867),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2631),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2634),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2587),
.Y(n_3105)
);

INVx1_ASAP7_75t_SL g3106 ( 
.A(n_2730),
.Y(n_3106)
);

OR2x6_ASAP7_75t_L g3107 ( 
.A(n_2601),
.B(n_1400),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2592),
.Y(n_3108)
);

BUFx6f_ASAP7_75t_L g3109 ( 
.A(n_2675),
.Y(n_3109)
);

OR2x6_ASAP7_75t_L g3110 ( 
.A(n_2610),
.B(n_1406),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2597),
.Y(n_3111)
);

INVx3_ASAP7_75t_L g3112 ( 
.A(n_2675),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2594),
.Y(n_3113)
);

NOR2xp33_ASAP7_75t_L g3114 ( 
.A(n_2877),
.B(n_1497),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2827),
.B(n_1499),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2595),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2781),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2783),
.Y(n_3118)
);

OAI22xp5_ASAP7_75t_L g3119 ( 
.A1(n_2731),
.A2(n_1600),
.B1(n_1602),
.B2(n_1593),
.Y(n_3119)
);

AOI22xp5_ASAP7_75t_L g3120 ( 
.A1(n_2679),
.A2(n_2705),
.B1(n_2873),
.B2(n_2800),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2784),
.Y(n_3121)
);

NAND2xp33_ASAP7_75t_L g3122 ( 
.A(n_2679),
.B(n_1608),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2599),
.Y(n_3123)
);

CKINVDCx20_ASAP7_75t_R g3124 ( 
.A(n_2753),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_2667),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2692),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2688),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2792),
.Y(n_3128)
);

INVx3_ASAP7_75t_L g3129 ( 
.A(n_2688),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2894),
.Y(n_3130)
);

INVx4_ASAP7_75t_L g3131 ( 
.A(n_2898),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_2896),
.B(n_2846),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2893),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2902),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2895),
.Y(n_3135)
);

AND2x6_ASAP7_75t_L g3136 ( 
.A(n_3008),
.B(n_2887),
.Y(n_3136)
);

OR2x6_ASAP7_75t_L g3137 ( 
.A(n_2937),
.B(n_2773),
.Y(n_3137)
);

CKINVDCx5p33_ASAP7_75t_R g3138 ( 
.A(n_2930),
.Y(n_3138)
);

BUFx3_ASAP7_75t_L g3139 ( 
.A(n_2889),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2900),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_L g3141 ( 
.A(n_2935),
.B(n_2856),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_2918),
.B(n_2779),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2904),
.B(n_2908),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_2889),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2916),
.Y(n_3145)
);

NAND2x1p5_ASAP7_75t_L g3146 ( 
.A(n_2936),
.B(n_2808),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2903),
.B(n_2849),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2905),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2906),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2913),
.B(n_2845),
.Y(n_3150)
);

AND2x4_ASAP7_75t_L g3151 ( 
.A(n_2938),
.B(n_2588),
.Y(n_3151)
);

NAND2x1p5_ASAP7_75t_L g3152 ( 
.A(n_2977),
.B(n_2812),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2923),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2928),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_3098),
.B(n_2847),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2909),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2910),
.Y(n_3157)
);

AO22x2_ASAP7_75t_L g3158 ( 
.A1(n_3115),
.A2(n_2878),
.B1(n_2888),
.B2(n_2711),
.Y(n_3158)
);

INVx3_ASAP7_75t_L g3159 ( 
.A(n_2897),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_2912),
.B(n_2771),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2931),
.Y(n_3161)
);

BUFx3_ASAP7_75t_L g3162 ( 
.A(n_2897),
.Y(n_3162)
);

NAND2x1p5_ASAP7_75t_L g3163 ( 
.A(n_3006),
.B(n_2812),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2942),
.Y(n_3164)
);

BUFx3_ASAP7_75t_L g3165 ( 
.A(n_2915),
.Y(n_3165)
);

BUFx2_ASAP7_75t_L g3166 ( 
.A(n_2919),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2973),
.B(n_2818),
.Y(n_3167)
);

AND2x2_ASAP7_75t_SL g3168 ( 
.A(n_2992),
.B(n_2874),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2943),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2911),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2929),
.B(n_2853),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2944),
.Y(n_3172)
);

BUFx6f_ASAP7_75t_L g3173 ( 
.A(n_2915),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2917),
.Y(n_3174)
);

INVx4_ASAP7_75t_L g3175 ( 
.A(n_2898),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_2964),
.Y(n_3176)
);

INVx1_ASAP7_75t_SL g3177 ( 
.A(n_2934),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_3031),
.B(n_2649),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2958),
.B(n_2794),
.Y(n_3179)
);

AND3x4_ASAP7_75t_L g3180 ( 
.A(n_3043),
.B(n_2884),
.C(n_2881),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2920),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2967),
.B(n_2865),
.Y(n_3182)
);

OA22x2_ASAP7_75t_L g3183 ( 
.A1(n_3120),
.A2(n_2682),
.B1(n_2778),
.B2(n_2715),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2946),
.Y(n_3184)
);

HB1xp67_ASAP7_75t_L g3185 ( 
.A(n_2941),
.Y(n_3185)
);

BUFx6f_ASAP7_75t_L g3186 ( 
.A(n_2964),
.Y(n_3186)
);

INVx4_ASAP7_75t_L g3187 ( 
.A(n_2970),
.Y(n_3187)
);

INVx6_ASAP7_75t_L g3188 ( 
.A(n_2970),
.Y(n_3188)
);

INVx3_ASAP7_75t_L g3189 ( 
.A(n_3019),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2980),
.B(n_2786),
.Y(n_3190)
);

AO22x2_ASAP7_75t_L g3191 ( 
.A1(n_3088),
.A2(n_2766),
.B1(n_2882),
.B2(n_1417),
.Y(n_3191)
);

AOI22xp5_ASAP7_75t_SL g3192 ( 
.A1(n_2985),
.A2(n_3016),
.B1(n_2989),
.B2(n_2940),
.Y(n_3192)
);

INVx3_ASAP7_75t_L g3193 ( 
.A(n_3019),
.Y(n_3193)
);

AND2x4_ASAP7_75t_L g3194 ( 
.A(n_2907),
.B(n_2732),
.Y(n_3194)
);

BUFx6f_ASAP7_75t_L g3195 ( 
.A(n_3069),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2924),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_3005),
.B(n_2705),
.Y(n_3197)
);

AOI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_3114),
.A2(n_2621),
.B1(n_2782),
.B2(n_2804),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2948),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2952),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2955),
.Y(n_3201)
);

OR2x6_ASAP7_75t_L g3202 ( 
.A(n_2937),
.B(n_2885),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3004),
.Y(n_3203)
);

BUFx2_ASAP7_75t_L g3204 ( 
.A(n_2993),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3010),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3056),
.Y(n_3206)
);

INVx4_ASAP7_75t_L g3207 ( 
.A(n_3101),
.Y(n_3207)
);

BUFx2_ASAP7_75t_L g3208 ( 
.A(n_3045),
.Y(n_3208)
);

AND2x4_ASAP7_75t_L g3209 ( 
.A(n_3054),
.B(n_2798),
.Y(n_3209)
);

CKINVDCx5p33_ASAP7_75t_R g3210 ( 
.A(n_2996),
.Y(n_3210)
);

OR2x2_ASAP7_75t_L g3211 ( 
.A(n_3034),
.B(n_2886),
.Y(n_3211)
);

BUFx2_ASAP7_75t_L g3212 ( 
.A(n_3028),
.Y(n_3212)
);

INVx2_ASAP7_75t_SL g3213 ( 
.A(n_3038),
.Y(n_3213)
);

NAND3xp33_ASAP7_75t_L g3214 ( 
.A(n_3089),
.B(n_2578),
.C(n_2862),
.Y(n_3214)
);

INVx4_ASAP7_75t_L g3215 ( 
.A(n_3101),
.Y(n_3215)
);

INVx2_ASAP7_75t_SL g3216 ( 
.A(n_3042),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3017),
.B(n_2976),
.Y(n_3217)
);

CKINVDCx20_ASAP7_75t_R g3218 ( 
.A(n_2899),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3013),
.B(n_3057),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2933),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_L g3221 ( 
.A1(n_2972),
.A2(n_2806),
.B1(n_1327),
.B2(n_2627),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2939),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_2947),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2956),
.Y(n_3224)
);

INVx8_ASAP7_75t_L g3225 ( 
.A(n_3078),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_L g3226 ( 
.A(n_3069),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2959),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_3106),
.B(n_2801),
.Y(n_3228)
);

INVx6_ASAP7_75t_L g3229 ( 
.A(n_3109),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3061),
.Y(n_3230)
);

INVx3_ASAP7_75t_L g3231 ( 
.A(n_3109),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3063),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3070),
.Y(n_3233)
);

BUFx6f_ASAP7_75t_L g3234 ( 
.A(n_3127),
.Y(n_3234)
);

INVx3_ASAP7_75t_L g3235 ( 
.A(n_3127),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_3058),
.B(n_2589),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2960),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3062),
.B(n_1615),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2962),
.Y(n_3239)
);

BUFx6f_ASAP7_75t_L g3240 ( 
.A(n_3092),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_2951),
.B(n_2802),
.Y(n_3241)
);

AND2x4_ASAP7_75t_L g3242 ( 
.A(n_2995),
.B(n_2811),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3076),
.B(n_1616),
.Y(n_3243)
);

AND2x4_ASAP7_75t_L g3244 ( 
.A(n_3022),
.B(n_2813),
.Y(n_3244)
);

CKINVDCx5p33_ASAP7_75t_R g3245 ( 
.A(n_3125),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3074),
.Y(n_3246)
);

AND2x4_ASAP7_75t_L g3247 ( 
.A(n_3079),
.B(n_2591),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_2968),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2969),
.Y(n_3249)
);

BUFx2_ASAP7_75t_L g3250 ( 
.A(n_3047),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_2972),
.A2(n_2611),
.B1(n_2757),
.B2(n_1384),
.Y(n_3251)
);

BUFx3_ASAP7_75t_L g3252 ( 
.A(n_3053),
.Y(n_3252)
);

AND2x2_ASAP7_75t_SL g3253 ( 
.A(n_3046),
.B(n_2691),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2990),
.B(n_1620),
.Y(n_3254)
);

BUFx3_ASAP7_75t_L g3255 ( 
.A(n_2892),
.Y(n_3255)
);

BUFx10_ASAP7_75t_L g3256 ( 
.A(n_2997),
.Y(n_3256)
);

BUFx6f_ASAP7_75t_L g3257 ( 
.A(n_2901),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2961),
.Y(n_3258)
);

BUFx6f_ASAP7_75t_L g3259 ( 
.A(n_2914),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2971),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_3040),
.B(n_2850),
.Y(n_3261)
);

BUFx6f_ASAP7_75t_L g3262 ( 
.A(n_2926),
.Y(n_3262)
);

INVx4_ASAP7_75t_L g3263 ( 
.A(n_3044),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2966),
.Y(n_3264)
);

HB1xp67_ASAP7_75t_L g3265 ( 
.A(n_2954),
.Y(n_3265)
);

INVx3_ASAP7_75t_L g3266 ( 
.A(n_2932),
.Y(n_3266)
);

OR2x2_ASAP7_75t_L g3267 ( 
.A(n_3000),
.B(n_3007),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_2974),
.Y(n_3268)
);

NAND2x1p5_ASAP7_75t_L g3269 ( 
.A(n_2965),
.B(n_2637),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_2981),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_3085),
.B(n_2662),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2978),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_2945),
.B(n_1627),
.Y(n_3273)
);

BUFx3_ASAP7_75t_L g3274 ( 
.A(n_2979),
.Y(n_3274)
);

INVx4_ASAP7_75t_L g3275 ( 
.A(n_2991),
.Y(n_3275)
);

INVx1_ASAP7_75t_SL g3276 ( 
.A(n_3049),
.Y(n_3276)
);

OR2x6_ASAP7_75t_L g3277 ( 
.A(n_2921),
.B(n_2691),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2984),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3091),
.B(n_1628),
.Y(n_3279)
);

AND2x4_ASAP7_75t_L g3280 ( 
.A(n_3087),
.B(n_2703),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_2927),
.B(n_2704),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2982),
.Y(n_3282)
);

AND2x4_ASAP7_75t_L g3283 ( 
.A(n_3126),
.B(n_2764),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2986),
.Y(n_3284)
);

AND2x4_ASAP7_75t_L g3285 ( 
.A(n_3059),
.B(n_2777),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3075),
.B(n_1634),
.Y(n_3286)
);

AND2x6_ASAP7_75t_L g3287 ( 
.A(n_3060),
.B(n_2851),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2987),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2988),
.Y(n_3289)
);

AND2x4_ASAP7_75t_L g3290 ( 
.A(n_3151),
.B(n_3112),
.Y(n_3290)
);

NOR2xp33_ASAP7_75t_L g3291 ( 
.A(n_3141),
.B(n_2963),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3133),
.Y(n_3292)
);

BUFx3_ASAP7_75t_L g3293 ( 
.A(n_3229),
.Y(n_3293)
);

BUFx6f_ASAP7_75t_SL g3294 ( 
.A(n_3252),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3143),
.B(n_2957),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3179),
.B(n_2890),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3134),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3130),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_SL g3299 ( 
.A(n_3267),
.B(n_2925),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_L g3300 ( 
.A(n_3177),
.B(n_3020),
.Y(n_3300)
);

INVx2_ASAP7_75t_SL g3301 ( 
.A(n_3204),
.Y(n_3301)
);

AO221x1_ASAP7_75t_L g3302 ( 
.A1(n_3191),
.A2(n_3119),
.B1(n_3129),
.B2(n_3105),
.C(n_3111),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_3276),
.B(n_2950),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_3147),
.B(n_3103),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_3217),
.B(n_2994),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_SL g3306 ( 
.A(n_3219),
.B(n_3104),
.Y(n_3306)
);

NOR2xp67_ASAP7_75t_L g3307 ( 
.A(n_3263),
.B(n_3093),
.Y(n_3307)
);

AND2x6_ASAP7_75t_L g3308 ( 
.A(n_3167),
.B(n_3041),
.Y(n_3308)
);

NOR3xp33_ASAP7_75t_L g3309 ( 
.A(n_3214),
.B(n_3122),
.C(n_2949),
.Y(n_3309)
);

NAND2xp33_ASAP7_75t_L g3310 ( 
.A(n_3287),
.B(n_2972),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3171),
.B(n_2998),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3135),
.Y(n_3312)
);

OR2x2_ASAP7_75t_L g3313 ( 
.A(n_3166),
.B(n_2891),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_SL g3314 ( 
.A(n_3138),
.B(n_3083),
.Y(n_3314)
);

INVx3_ASAP7_75t_L g3315 ( 
.A(n_3188),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3140),
.B(n_2999),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_3197),
.B(n_2983),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3148),
.Y(n_3318)
);

BUFx8_ASAP7_75t_L g3319 ( 
.A(n_3208),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3145),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3183),
.A2(n_3086),
.B1(n_3055),
.B2(n_3011),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3153),
.B(n_3009),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3154),
.B(n_3001),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3161),
.B(n_3029),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_3132),
.B(n_3002),
.Y(n_3325)
);

INVx2_ASAP7_75t_SL g3326 ( 
.A(n_3212),
.Y(n_3326)
);

INVx2_ASAP7_75t_SL g3327 ( 
.A(n_3213),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3164),
.B(n_3030),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3169),
.B(n_3014),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3149),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3172),
.Y(n_3331)
);

INVxp67_ASAP7_75t_SL g3332 ( 
.A(n_3185),
.Y(n_3332)
);

AOI22xp33_ASAP7_75t_L g3333 ( 
.A1(n_3184),
.A2(n_3023),
.B1(n_3027),
.B2(n_3018),
.Y(n_3333)
);

AND2x6_ASAP7_75t_SL g3334 ( 
.A(n_3202),
.B(n_2953),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3199),
.B(n_3032),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3200),
.B(n_3012),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3201),
.B(n_3033),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_3211),
.B(n_3084),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3203),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3205),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3206),
.Y(n_3341)
);

INVxp67_ASAP7_75t_L g3342 ( 
.A(n_3236),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3245),
.B(n_3082),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_3216),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3230),
.Y(n_3345)
);

INVx3_ASAP7_75t_L g3346 ( 
.A(n_3131),
.Y(n_3346)
);

NAND3xp33_ASAP7_75t_SL g3347 ( 
.A(n_3210),
.B(n_3124),
.C(n_3081),
.Y(n_3347)
);

INVx1_ASAP7_75t_SL g3348 ( 
.A(n_3250),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3232),
.B(n_3067),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3233),
.B(n_3050),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_SL g3351 ( 
.A(n_3150),
.B(n_3198),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_3160),
.B(n_3078),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3156),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3246),
.B(n_3080),
.Y(n_3354)
);

OAI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_3190),
.A2(n_3003),
.B(n_3073),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3258),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3281),
.B(n_3107),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3264),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3157),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3170),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3174),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3272),
.B(n_3282),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_3253),
.B(n_3284),
.Y(n_3363)
);

INVx3_ASAP7_75t_L g3364 ( 
.A(n_3175),
.Y(n_3364)
);

AND2x6_ASAP7_75t_SL g3365 ( 
.A(n_3277),
.B(n_2953),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3289),
.B(n_3035),
.Y(n_3366)
);

AOI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3180),
.A2(n_3015),
.B1(n_3021),
.B2(n_3036),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3254),
.B(n_3037),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3142),
.B(n_3039),
.Y(n_3369)
);

HB1xp67_ASAP7_75t_L g3370 ( 
.A(n_3234),
.Y(n_3370)
);

AOI22xp33_ASAP7_75t_L g3371 ( 
.A1(n_3181),
.A2(n_3052),
.B1(n_3064),
.B2(n_3051),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_3288),
.A2(n_3072),
.B1(n_3068),
.B2(n_3026),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_SL g3373 ( 
.A(n_3286),
.B(n_3077),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3273),
.B(n_3025),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_3178),
.B(n_3102),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3238),
.B(n_3094),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3261),
.B(n_3107),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3265),
.B(n_3095),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3196),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3279),
.B(n_3099),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3220),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3243),
.B(n_3090),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3192),
.B(n_3096),
.Y(n_3383)
);

OR2x2_ASAP7_75t_L g3384 ( 
.A(n_3228),
.B(n_3066),
.Y(n_3384)
);

BUFx6f_ASAP7_75t_L g3385 ( 
.A(n_3234),
.Y(n_3385)
);

BUFx3_ASAP7_75t_L g3386 ( 
.A(n_3144),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3222),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3155),
.B(n_3241),
.Y(n_3388)
);

OR2x2_ASAP7_75t_L g3389 ( 
.A(n_3223),
.B(n_3113),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_3224),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3227),
.B(n_3097),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3237),
.B(n_3100),
.Y(n_3392)
);

A2O1A1Ixp33_ASAP7_75t_L g3393 ( 
.A1(n_3182),
.A2(n_3108),
.B(n_3123),
.C(n_3116),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3239),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_SL g3395 ( 
.A(n_3248),
.B(n_3117),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3249),
.Y(n_3396)
);

INVx3_ASAP7_75t_L g3397 ( 
.A(n_3240),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3260),
.B(n_3118),
.Y(n_3398)
);

AOI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_3287),
.A2(n_3128),
.B1(n_3121),
.B2(n_1643),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3268),
.B(n_3270),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_3275),
.B(n_2975),
.Y(n_3401)
);

A2O1A1Ixp33_ASAP7_75t_L g3402 ( 
.A1(n_3278),
.A2(n_2738),
.B(n_1419),
.C(n_1420),
.Y(n_3402)
);

INVxp67_ASAP7_75t_L g3403 ( 
.A(n_3173),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_3136),
.A2(n_1384),
.B1(n_1405),
.B2(n_1268),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3266),
.B(n_1642),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_SL g3406 ( 
.A(n_3194),
.B(n_3048),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3136),
.B(n_1648),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3242),
.Y(n_3408)
);

AOI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_3244),
.A2(n_1655),
.B1(n_1656),
.B2(n_1653),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3159),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3176),
.Y(n_3411)
);

AOI22xp33_ASAP7_75t_L g3412 ( 
.A1(n_3168),
.A2(n_1405),
.B1(n_1421),
.B2(n_1384),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3189),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3259),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3256),
.B(n_3110),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3158),
.A2(n_1668),
.B1(n_1670),
.B2(n_1662),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3193),
.B(n_1689),
.Y(n_3417)
);

NOR2xp33_ASAP7_75t_SL g3418 ( 
.A(n_3218),
.B(n_3071),
.Y(n_3418)
);

A2O1A1Ixp33_ASAP7_75t_L g3419 ( 
.A1(n_3221),
.A2(n_1415),
.B(n_1429),
.C(n_1426),
.Y(n_3419)
);

OAI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3251),
.A2(n_1698),
.B(n_1690),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3231),
.B(n_1699),
.Y(n_3421)
);

AOI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_3291),
.A2(n_3338),
.B1(n_3325),
.B2(n_3300),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3296),
.B(n_3209),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3388),
.A2(n_3110),
.B1(n_3283),
.B2(n_3271),
.Y(n_3424)
);

INVx3_ASAP7_75t_L g3425 ( 
.A(n_3293),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3295),
.B(n_3235),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_3301),
.B(n_3186),
.Y(n_3427)
);

INVx1_ASAP7_75t_SL g3428 ( 
.A(n_3348),
.Y(n_3428)
);

INVx3_ASAP7_75t_L g3429 ( 
.A(n_3315),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3298),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3312),
.Y(n_3431)
);

BUFx3_ASAP7_75t_L g3432 ( 
.A(n_3385),
.Y(n_3432)
);

BUFx2_ASAP7_75t_L g3433 ( 
.A(n_3326),
.Y(n_3433)
);

HB1xp67_ASAP7_75t_L g3434 ( 
.A(n_3385),
.Y(n_3434)
);

INVx3_ASAP7_75t_L g3435 ( 
.A(n_3397),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3320),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3311),
.B(n_3259),
.Y(n_3437)
);

AOI22xp5_ASAP7_75t_L g3438 ( 
.A1(n_3317),
.A2(n_3303),
.B1(n_3299),
.B2(n_3357),
.Y(n_3438)
);

BUFx4f_ASAP7_75t_L g3439 ( 
.A(n_3308),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3331),
.Y(n_3440)
);

CKINVDCx5p33_ASAP7_75t_R g3441 ( 
.A(n_3294),
.Y(n_3441)
);

INVx4_ASAP7_75t_L g3442 ( 
.A(n_3386),
.Y(n_3442)
);

BUFx2_ASAP7_75t_L g3443 ( 
.A(n_3332),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3305),
.B(n_3376),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3339),
.Y(n_3445)
);

BUFx2_ASAP7_75t_L g3446 ( 
.A(n_3370),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_3342),
.B(n_3269),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3380),
.B(n_3257),
.Y(n_3448)
);

BUFx2_ASAP7_75t_L g3449 ( 
.A(n_3377),
.Y(n_3449)
);

NOR2xp33_ASAP7_75t_L g3450 ( 
.A(n_3363),
.B(n_3187),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3340),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3341),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_3378),
.B(n_3195),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3368),
.B(n_3362),
.Y(n_3454)
);

OR2x2_ASAP7_75t_L g3455 ( 
.A(n_3313),
.B(n_3146),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3374),
.B(n_3262),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3345),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3290),
.Y(n_3458)
);

AOI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3375),
.A2(n_3247),
.B1(n_3280),
.B2(n_3065),
.Y(n_3459)
);

OR2x6_ASAP7_75t_L g3460 ( 
.A(n_3327),
.B(n_3225),
.Y(n_3460)
);

AOI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3309),
.A2(n_3024),
.B1(n_3285),
.B2(n_3137),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3382),
.B(n_3139),
.Y(n_3462)
);

AOI22xp5_ASAP7_75t_L g3463 ( 
.A1(n_3369),
.A2(n_3024),
.B1(n_2921),
.B2(n_3152),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3356),
.B(n_3162),
.Y(n_3464)
);

HB1xp67_ASAP7_75t_L g3465 ( 
.A(n_3344),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_3337),
.B(n_3226),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3358),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3323),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3324),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3328),
.Y(n_3470)
);

OAI22xp5_ASAP7_75t_L g3471 ( 
.A1(n_3351),
.A2(n_3274),
.B1(n_3255),
.B2(n_3165),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_SL g3472 ( 
.A(n_3349),
.B(n_3207),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3316),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3366),
.B(n_3163),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3302),
.A2(n_1439),
.B1(n_1440),
.B2(n_1436),
.Y(n_3475)
);

CKINVDCx5p33_ASAP7_75t_R g3476 ( 
.A(n_3319),
.Y(n_3476)
);

INVx5_ASAP7_75t_L g3477 ( 
.A(n_3365),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3321),
.B(n_3215),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3322),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3292),
.Y(n_3480)
);

AND2x4_ASAP7_75t_L g3481 ( 
.A(n_3414),
.B(n_2704),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3297),
.Y(n_3482)
);

BUFx3_ASAP7_75t_L g3483 ( 
.A(n_3346),
.Y(n_3483)
);

INVx5_ASAP7_75t_L g3484 ( 
.A(n_3334),
.Y(n_3484)
);

AOI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3314),
.A2(n_1701),
.B1(n_1702),
.B2(n_1700),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3336),
.Y(n_3486)
);

OR2x6_ASAP7_75t_L g3487 ( 
.A(n_3403),
.B(n_2713),
.Y(n_3487)
);

BUFx2_ASAP7_75t_L g3488 ( 
.A(n_3384),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3318),
.Y(n_3489)
);

INVx5_ASAP7_75t_L g3490 ( 
.A(n_3364),
.Y(n_3490)
);

BUFx8_ASAP7_75t_L g3491 ( 
.A(n_3410),
.Y(n_3491)
);

AND2x4_ASAP7_75t_L g3492 ( 
.A(n_3408),
.B(n_2713),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3329),
.Y(n_3493)
);

INVx5_ASAP7_75t_L g3494 ( 
.A(n_3308),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3354),
.B(n_1711),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3335),
.B(n_1712),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3330),
.Y(n_3497)
);

AND3x1_ASAP7_75t_L g3498 ( 
.A(n_3416),
.B(n_2642),
.C(n_2855),
.Y(n_3498)
);

HB1xp67_ASAP7_75t_SL g3499 ( 
.A(n_3415),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3353),
.Y(n_3500)
);

INVx2_ASAP7_75t_SL g3501 ( 
.A(n_3406),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3400),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3308),
.B(n_1714),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3379),
.Y(n_3504)
);

BUFx3_ASAP7_75t_L g3505 ( 
.A(n_3411),
.Y(n_3505)
);

AOI22xp33_ASAP7_75t_L g3506 ( 
.A1(n_3412),
.A2(n_1465),
.B1(n_1471),
.B2(n_1464),
.Y(n_3506)
);

BUFx6f_ASAP7_75t_L g3507 ( 
.A(n_3413),
.Y(n_3507)
);

AOI22xp5_ASAP7_75t_SL g3508 ( 
.A1(n_3352),
.A2(n_1501),
.B1(n_1502),
.B2(n_1500),
.Y(n_3508)
);

INVx2_ASAP7_75t_SL g3509 ( 
.A(n_3343),
.Y(n_3509)
);

INVx2_ASAP7_75t_SL g3510 ( 
.A(n_3383),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3359),
.Y(n_3511)
);

HB1xp67_ASAP7_75t_L g3512 ( 
.A(n_3306),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_SL g3513 ( 
.A(n_3367),
.B(n_2727),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3360),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3304),
.B(n_2922),
.Y(n_3515)
);

INVx5_ASAP7_75t_L g3516 ( 
.A(n_3361),
.Y(n_3516)
);

BUFx6f_ASAP7_75t_L g3517 ( 
.A(n_3401),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3381),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3387),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3390),
.Y(n_3520)
);

INVxp67_ASAP7_75t_L g3521 ( 
.A(n_3418),
.Y(n_3521)
);

INVx3_ASAP7_75t_L g3522 ( 
.A(n_3389),
.Y(n_3522)
);

AOI22xp5_ASAP7_75t_L g3523 ( 
.A1(n_3347),
.A2(n_1730),
.B1(n_1739),
.B2(n_1718),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3394),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3420),
.A2(n_1484),
.B1(n_1486),
.B2(n_1481),
.Y(n_3525)
);

AND3x1_ASAP7_75t_SL g3526 ( 
.A(n_3396),
.B(n_1490),
.C(n_1488),
.Y(n_3526)
);

BUFx3_ASAP7_75t_L g3527 ( 
.A(n_3417),
.Y(n_3527)
);

CKINVDCx5p33_ASAP7_75t_R g3528 ( 
.A(n_3407),
.Y(n_3528)
);

OAI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_3422),
.A2(n_3409),
.B1(n_3333),
.B2(n_3371),
.Y(n_3529)
);

BUFx2_ASAP7_75t_L g3530 ( 
.A(n_3433),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3444),
.B(n_3350),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3445),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_SL g3533 ( 
.A(n_3438),
.B(n_3399),
.Y(n_3533)
);

AOI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3454),
.A2(n_3355),
.B(n_3310),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_SL g3535 ( 
.A(n_3510),
.B(n_3509),
.Y(n_3535)
);

AND2x2_ASAP7_75t_L g3536 ( 
.A(n_3522),
.B(n_3372),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3467),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3468),
.B(n_3391),
.Y(n_3538)
);

AND2x4_ASAP7_75t_L g3539 ( 
.A(n_3425),
.B(n_3442),
.Y(n_3539)
);

OAI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_3478),
.A2(n_3421),
.B1(n_3405),
.B2(n_3404),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3423),
.A2(n_3402),
.B(n_3373),
.Y(n_3541)
);

OAI22xp5_ASAP7_75t_L g3542 ( 
.A1(n_3469),
.A2(n_3307),
.B1(n_3392),
.B2(n_3393),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3470),
.B(n_3398),
.Y(n_3543)
);

AO32x2_ASAP7_75t_L g3544 ( 
.A1(n_3471),
.A2(n_3419),
.A3(n_3395),
.B1(n_3),
.B2(n_1),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3430),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3480),
.Y(n_3546)
);

NOR3xp33_ASAP7_75t_SL g3547 ( 
.A(n_3528),
.B(n_1507),
.C(n_1505),
.Y(n_3547)
);

HB1xp67_ASAP7_75t_L g3548 ( 
.A(n_3428),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_R g3549 ( 
.A(n_3441),
.B(n_2727),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3525),
.A2(n_1421),
.B(n_1405),
.Y(n_3550)
);

OAI21x1_ASAP7_75t_L g3551 ( 
.A1(n_3475),
.A2(n_1506),
.B(n_1503),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_R g3552 ( 
.A(n_3476),
.B(n_3429),
.Y(n_3552)
);

AND2x4_ASAP7_75t_L g3553 ( 
.A(n_3435),
.B(n_2733),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3486),
.B(n_1508),
.Y(n_3554)
);

HB1xp67_ASAP7_75t_L g3555 ( 
.A(n_3443),
.Y(n_3555)
);

O2A1O1Ixp5_ASAP7_75t_SL g3556 ( 
.A1(n_3513),
.A2(n_1516),
.B(n_1527),
.C(n_1512),
.Y(n_3556)
);

INVx4_ASAP7_75t_L g3557 ( 
.A(n_3490),
.Y(n_3557)
);

INVx1_ASAP7_75t_SL g3558 ( 
.A(n_3488),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3493),
.B(n_1509),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3473),
.B(n_1511),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3482),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_SL g3562 ( 
.A(n_3527),
.B(n_2733),
.Y(n_3562)
);

A2O1A1Ixp33_ASAP7_75t_SL g3563 ( 
.A1(n_3515),
.A2(n_2857),
.B(n_2854),
.C(n_1422),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3479),
.B(n_1513),
.Y(n_3564)
);

INVx3_ASAP7_75t_L g3565 ( 
.A(n_3483),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3502),
.B(n_1519),
.Y(n_3566)
);

OR2x6_ASAP7_75t_L g3567 ( 
.A(n_3460),
.B(n_2736),
.Y(n_3567)
);

NOR2xp33_ASAP7_75t_L g3568 ( 
.A(n_3449),
.B(n_2736),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3439),
.A2(n_1561),
.B(n_1421),
.Y(n_3569)
);

INVx4_ASAP7_75t_L g3570 ( 
.A(n_3490),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_SL g3571 ( 
.A(n_3450),
.B(n_2742),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3446),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3516),
.A2(n_1523),
.B1(n_1525),
.B2(n_1522),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3506),
.A2(n_1533),
.B1(n_1534),
.B2(n_1532),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3462),
.B(n_1526),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3426),
.B(n_1530),
.Y(n_3576)
);

OAI21xp33_ASAP7_75t_L g3577 ( 
.A1(n_3495),
.A2(n_3463),
.B(n_3496),
.Y(n_3577)
);

BUFx3_ASAP7_75t_L g3578 ( 
.A(n_3432),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3472),
.A2(n_2054),
.B(n_1561),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3431),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3494),
.A2(n_2054),
.B(n_1561),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3448),
.B(n_1535),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_3494),
.A2(n_2054),
.B(n_1753),
.Y(n_3583)
);

O2A1O1Ixp5_ASAP7_75t_L g3584 ( 
.A1(n_3466),
.A2(n_1545),
.B(n_1547),
.C(n_1544),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3489),
.Y(n_3585)
);

OAI21xp33_ASAP7_75t_L g3586 ( 
.A1(n_3456),
.A2(n_1540),
.B(n_1537),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3474),
.A2(n_1769),
.B(n_1742),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_3503),
.A2(n_1779),
.B(n_1770),
.Y(n_3588)
);

INVx3_ASAP7_75t_L g3589 ( 
.A(n_3517),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3437),
.B(n_1541),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3512),
.B(n_1543),
.Y(n_3591)
);

OAI22xp5_ASAP7_75t_L g3592 ( 
.A1(n_3516),
.A2(n_1548),
.B1(n_1549),
.B2(n_1546),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_SL g3593 ( 
.A(n_3517),
.B(n_2742),
.Y(n_3593)
);

HB1xp67_ASAP7_75t_L g3594 ( 
.A(n_3465),
.Y(n_3594)
);

NAND3xp33_ASAP7_75t_L g3595 ( 
.A(n_3508),
.B(n_1555),
.C(n_1554),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3521),
.B(n_2743),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3436),
.A2(n_3451),
.B(n_3440),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_3447),
.B(n_1553),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3452),
.A2(n_1792),
.B(n_1790),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3455),
.B(n_1558),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_SL g3601 ( 
.A(n_3459),
.B(n_2743),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3497),
.B(n_1559),
.Y(n_3602)
);

OAI22x1_ASAP7_75t_L g3603 ( 
.A1(n_3461),
.A2(n_1562),
.B1(n_1576),
.B2(n_1563),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3500),
.B(n_1560),
.Y(n_3604)
);

O2A1O1Ixp33_ASAP7_75t_L g3605 ( 
.A1(n_3453),
.A2(n_1584),
.B(n_1596),
.C(n_1581),
.Y(n_3605)
);

A2O1A1Ixp33_ASAP7_75t_L g3606 ( 
.A1(n_3501),
.A2(n_1613),
.B(n_1640),
.C(n_1599),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_3457),
.A2(n_1797),
.B(n_1796),
.Y(n_3607)
);

CKINVDCx16_ASAP7_75t_R g3608 ( 
.A(n_3499),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3504),
.A2(n_1810),
.B(n_1803),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3511),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3518),
.A2(n_1818),
.B(n_1817),
.Y(n_3611)
);

INVxp67_ASAP7_75t_L g3612 ( 
.A(n_3434),
.Y(n_3612)
);

NAND3xp33_ASAP7_75t_SL g3613 ( 
.A(n_3424),
.B(n_1570),
.C(n_1568),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3514),
.B(n_3520),
.Y(n_3614)
);

AND2x6_ASAP7_75t_L g3615 ( 
.A(n_3519),
.B(n_1641),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3524),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3464),
.A2(n_1837),
.B(n_1821),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3498),
.B(n_1646),
.Y(n_3618)
);

AOI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_3427),
.A2(n_1846),
.B(n_1838),
.Y(n_3619)
);

BUFx2_ASAP7_75t_L g3620 ( 
.A(n_3487),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_3523),
.A2(n_1850),
.B(n_1848),
.Y(n_3621)
);

AND2x4_ASAP7_75t_L g3622 ( 
.A(n_3460),
.B(n_2745),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3507),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3485),
.A2(n_1857),
.B(n_1856),
.Y(n_3624)
);

O2A1O1Ixp5_ASAP7_75t_L g3625 ( 
.A1(n_3492),
.A2(n_1659),
.B(n_1665),
.C(n_1647),
.Y(n_3625)
);

NAND2x1p5_ASAP7_75t_L g3626 ( 
.A(n_3505),
.B(n_2745),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3507),
.A2(n_1865),
.B(n_1863),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3481),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3487),
.Y(n_3629)
);

A2O1A1Ixp33_ASAP7_75t_L g3630 ( 
.A1(n_3526),
.A2(n_1674),
.B(n_1675),
.C(n_1672),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_3484),
.A2(n_1886),
.B(n_1872),
.Y(n_3631)
);

O2A1O1Ixp33_ASAP7_75t_L g3632 ( 
.A1(n_3484),
.A2(n_1705),
.B(n_1716),
.C(n_1687),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3458),
.B(n_1572),
.Y(n_3633)
);

O2A1O1Ixp33_ASAP7_75t_L g3634 ( 
.A1(n_3477),
.A2(n_1721),
.B(n_1722),
.C(n_1719),
.Y(n_3634)
);

BUFx6f_ASAP7_75t_L g3635 ( 
.A(n_3458),
.Y(n_3635)
);

OAI22xp5_ASAP7_75t_SL g3636 ( 
.A1(n_3477),
.A2(n_1582),
.B1(n_1585),
.B2(n_1575),
.Y(n_3636)
);

BUFx6f_ASAP7_75t_L g3637 ( 
.A(n_3491),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3444),
.B(n_1586),
.Y(n_3638)
);

INVx4_ASAP7_75t_L g3639 ( 
.A(n_3490),
.Y(n_3639)
);

BUFx2_ASAP7_75t_L g3640 ( 
.A(n_3572),
.Y(n_3640)
);

INVx4_ASAP7_75t_L g3641 ( 
.A(n_3539),
.Y(n_3641)
);

INVx3_ASAP7_75t_L g3642 ( 
.A(n_3589),
.Y(n_3642)
);

OAI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_3595),
.A2(n_2785),
.B1(n_2787),
.B2(n_2748),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3577),
.A2(n_1589),
.B1(n_1590),
.B2(n_1588),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3531),
.B(n_1595),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3545),
.Y(n_3646)
);

CKINVDCx5p33_ASAP7_75t_R g3647 ( 
.A(n_3552),
.Y(n_3647)
);

OR2x2_ASAP7_75t_L g3648 ( 
.A(n_3558),
.B(n_3555),
.Y(n_3648)
);

OAI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3608),
.A2(n_1603),
.B1(n_1607),
.B2(n_1598),
.Y(n_3649)
);

INVx3_ASAP7_75t_L g3650 ( 
.A(n_3565),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3580),
.Y(n_3651)
);

BUFx6f_ASAP7_75t_L g3652 ( 
.A(n_3578),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3635),
.Y(n_3653)
);

INVx3_ASAP7_75t_L g3654 ( 
.A(n_3557),
.Y(n_3654)
);

BUFx2_ASAP7_75t_L g3655 ( 
.A(n_3530),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3532),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3570),
.Y(n_3657)
);

AOI222xp33_ASAP7_75t_L g3658 ( 
.A1(n_3603),
.A2(n_1736),
.B1(n_1727),
.B2(n_1738),
.C1(n_1728),
.C2(n_1724),
.Y(n_3658)
);

INVx2_ASAP7_75t_SL g3659 ( 
.A(n_3635),
.Y(n_3659)
);

BUFx6f_ASAP7_75t_L g3660 ( 
.A(n_3639),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_SL g3661 ( 
.A1(n_3618),
.A2(n_1751),
.B1(n_1754),
.B2(n_1746),
.Y(n_3661)
);

INVx1_ASAP7_75t_SL g3662 ( 
.A(n_3548),
.Y(n_3662)
);

INVx5_ASAP7_75t_L g3663 ( 
.A(n_3567),
.Y(n_3663)
);

BUFx8_ASAP7_75t_L g3664 ( 
.A(n_3637),
.Y(n_3664)
);

INVx1_ASAP7_75t_SL g3665 ( 
.A(n_3594),
.Y(n_3665)
);

CKINVDCx20_ASAP7_75t_R g3666 ( 
.A(n_3549),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3616),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3536),
.B(n_1759),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3537),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3546),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3597),
.Y(n_3671)
);

AOI22xp33_ASAP7_75t_SL g3672 ( 
.A1(n_3529),
.A2(n_1765),
.B1(n_1785),
.B2(n_1764),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3538),
.B(n_1609),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3598),
.B(n_1804),
.Y(n_3674)
);

INVx3_ASAP7_75t_L g3675 ( 
.A(n_3623),
.Y(n_3675)
);

BUFx6f_ASAP7_75t_L g3676 ( 
.A(n_3620),
.Y(n_3676)
);

A2O1A1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_3533),
.A2(n_1811),
.B(n_1819),
.C(n_1809),
.Y(n_3677)
);

OR2x6_ASAP7_75t_L g3678 ( 
.A(n_3637),
.B(n_2748),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3561),
.Y(n_3679)
);

OR2x6_ASAP7_75t_L g3680 ( 
.A(n_3567),
.B(n_2785),
.Y(n_3680)
);

BUFx6f_ASAP7_75t_L g3681 ( 
.A(n_3553),
.Y(n_3681)
);

INVx3_ASAP7_75t_L g3682 ( 
.A(n_3626),
.Y(n_3682)
);

NAND2x1p5_ASAP7_75t_L g3683 ( 
.A(n_3535),
.B(n_2787),
.Y(n_3683)
);

CKINVDCx5p33_ASAP7_75t_R g3684 ( 
.A(n_3547),
.Y(n_3684)
);

BUFx12f_ASAP7_75t_L g3685 ( 
.A(n_3622),
.Y(n_3685)
);

AOI22xp5_ASAP7_75t_L g3686 ( 
.A1(n_3613),
.A2(n_1622),
.B1(n_1624),
.B2(n_1614),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3585),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3543),
.B(n_1625),
.Y(n_3688)
);

BUFx6f_ASAP7_75t_L g3689 ( 
.A(n_3593),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3534),
.A2(n_1888),
.B(n_1887),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3610),
.Y(n_3691)
);

BUFx6f_ASAP7_75t_L g3692 ( 
.A(n_3568),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3614),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3638),
.B(n_1630),
.Y(n_3694)
);

NOR2x1_ASAP7_75t_R g3695 ( 
.A(n_3601),
.B(n_2824),
.Y(n_3695)
);

O2A1O1Ixp33_ASAP7_75t_L g3696 ( 
.A1(n_3563),
.A2(n_3630),
.B(n_3634),
.C(n_3632),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3628),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3544),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3551),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3544),
.Y(n_3700)
);

AOI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_3615),
.A2(n_1633),
.B1(n_1635),
.B2(n_1632),
.Y(n_3701)
);

O2A1O1Ixp33_ASAP7_75t_SL g3702 ( 
.A1(n_3571),
.A2(n_1826),
.B(n_1830),
.C(n_1822),
.Y(n_3702)
);

NOR2xp67_ASAP7_75t_SL g3703 ( 
.A(n_3569),
.B(n_2848),
.Y(n_3703)
);

HB1xp67_ASAP7_75t_L g3704 ( 
.A(n_3612),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3576),
.B(n_1651),
.Y(n_3705)
);

INVx5_ASAP7_75t_L g3706 ( 
.A(n_3615),
.Y(n_3706)
);

AOI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3615),
.A2(n_1657),
.B1(n_1658),
.B2(n_1652),
.Y(n_3707)
);

BUFx6f_ASAP7_75t_L g3708 ( 
.A(n_3629),
.Y(n_3708)
);

BUFx8_ASAP7_75t_SL g3709 ( 
.A(n_3600),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_3541),
.A2(n_1898),
.B(n_1891),
.Y(n_3710)
);

BUFx3_ASAP7_75t_L g3711 ( 
.A(n_3596),
.Y(n_3711)
);

BUFx3_ASAP7_75t_L g3712 ( 
.A(n_3633),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3605),
.Y(n_3713)
);

NOR2xp33_ASAP7_75t_L g3714 ( 
.A(n_3582),
.B(n_2859),
.Y(n_3714)
);

BUFx6f_ASAP7_75t_L g3715 ( 
.A(n_3562),
.Y(n_3715)
);

INVx4_ASAP7_75t_L g3716 ( 
.A(n_3627),
.Y(n_3716)
);

INVx3_ASAP7_75t_L g3717 ( 
.A(n_3591),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3602),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3604),
.Y(n_3719)
);

O2A1O1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_3606),
.A2(n_1833),
.B(n_1839),
.C(n_1831),
.Y(n_3720)
);

OR2x2_ASAP7_75t_L g3721 ( 
.A(n_3590),
.B(n_1845),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3575),
.B(n_1852),
.Y(n_3722)
);

OAI22xp33_ASAP7_75t_L g3723 ( 
.A1(n_3554),
.A2(n_1664),
.B1(n_1666),
.B2(n_1663),
.Y(n_3723)
);

BUFx2_ASAP7_75t_L g3724 ( 
.A(n_3566),
.Y(n_3724)
);

AOI22xp33_ASAP7_75t_SL g3725 ( 
.A1(n_3540),
.A2(n_1859),
.B1(n_1870),
.B2(n_1855),
.Y(n_3725)
);

OR2x6_ASAP7_75t_SL g3726 ( 
.A(n_3542),
.B(n_1667),
.Y(n_3726)
);

BUFx6f_ASAP7_75t_L g3727 ( 
.A(n_3559),
.Y(n_3727)
);

BUFx2_ASAP7_75t_L g3728 ( 
.A(n_3560),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3564),
.B(n_3586),
.Y(n_3729)
);

BUFx2_ASAP7_75t_L g3730 ( 
.A(n_3573),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3584),
.B(n_1884),
.Y(n_3731)
);

AND2x4_ASAP7_75t_L g3732 ( 
.A(n_3587),
.B(n_2844),
.Y(n_3732)
);

INVx3_ASAP7_75t_L g3733 ( 
.A(n_3583),
.Y(n_3733)
);

A2O1A1Ixp33_ASAP7_75t_L g3734 ( 
.A1(n_3696),
.A2(n_3625),
.B(n_3550),
.C(n_3621),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3672),
.A2(n_3624),
.B1(n_1897),
.B2(n_1900),
.Y(n_3735)
);

AO32x2_ASAP7_75t_L g3736 ( 
.A1(n_3643),
.A2(n_3636),
.A3(n_3592),
.B1(n_3556),
.B2(n_3),
.Y(n_3736)
);

AOI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_3671),
.A2(n_3579),
.B(n_3588),
.Y(n_3737)
);

OAI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_3725),
.A2(n_3617),
.B(n_3611),
.Y(n_3738)
);

AOI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_3710),
.A2(n_3581),
.B(n_3609),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3667),
.Y(n_3740)
);

BUFx3_ASAP7_75t_L g3741 ( 
.A(n_3652),
.Y(n_3741)
);

OR2x6_ASAP7_75t_L g3742 ( 
.A(n_3641),
.B(n_3599),
.Y(n_3742)
);

AO31x2_ASAP7_75t_L g3743 ( 
.A1(n_3699),
.A2(n_3607),
.A3(n_1905),
.B(n_1909),
.Y(n_3743)
);

NOR2xp33_ASAP7_75t_L g3744 ( 
.A(n_3727),
.B(n_3631),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3662),
.B(n_3619),
.Y(n_3745)
);

AOI22xp5_ASAP7_75t_L g3746 ( 
.A1(n_3730),
.A2(n_3574),
.B1(n_1673),
.B2(n_1677),
.Y(n_3746)
);

CKINVDCx20_ASAP7_75t_R g3747 ( 
.A(n_3664),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3729),
.A2(n_3690),
.B(n_3716),
.Y(n_3748)
);

AO31x2_ASAP7_75t_L g3749 ( 
.A1(n_3698),
.A2(n_1914),
.A3(n_1924),
.B(n_1896),
.Y(n_3749)
);

O2A1O1Ixp33_ASAP7_75t_L g3750 ( 
.A1(n_3677),
.A2(n_1933),
.B(n_1939),
.C(n_1932),
.Y(n_3750)
);

AOI22xp5_ASAP7_75t_L g3751 ( 
.A1(n_3684),
.A2(n_1678),
.B1(n_1683),
.B2(n_1671),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3733),
.A2(n_1916),
.B(n_1901),
.Y(n_3752)
);

OAI21xp5_ASAP7_75t_L g3753 ( 
.A1(n_3686),
.A2(n_1941),
.B(n_1940),
.Y(n_3753)
);

CKINVDCx20_ASAP7_75t_R g3754 ( 
.A(n_3709),
.Y(n_3754)
);

INVx3_ASAP7_75t_L g3755 ( 
.A(n_3652),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3713),
.A2(n_1960),
.B1(n_1966),
.B2(n_1944),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3693),
.B(n_1684),
.Y(n_3757)
);

INVx3_ASAP7_75t_L g3758 ( 
.A(n_3692),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3718),
.A2(n_3719),
.B(n_3645),
.Y(n_3759)
);

BUFx2_ASAP7_75t_L g3760 ( 
.A(n_3640),
.Y(n_3760)
);

AOI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3732),
.A2(n_3694),
.B(n_3724),
.Y(n_3761)
);

BUFx6f_ASAP7_75t_L g3762 ( 
.A(n_3681),
.Y(n_3762)
);

O2A1O1Ixp33_ASAP7_75t_L g3763 ( 
.A1(n_3723),
.A2(n_1975),
.B(n_1989),
.C(n_1973),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3665),
.B(n_1686),
.Y(n_3764)
);

OAI21x1_ASAP7_75t_L g3765 ( 
.A1(n_3669),
.A2(n_2005),
.B(n_1992),
.Y(n_3765)
);

A2O1A1Ixp33_ASAP7_75t_L g3766 ( 
.A1(n_3720),
.A2(n_2020),
.B(n_2022),
.C(n_2018),
.Y(n_3766)
);

BUFx2_ASAP7_75t_R g3767 ( 
.A(n_3647),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_3728),
.A2(n_1922),
.B(n_1919),
.Y(n_3768)
);

O2A1O1Ixp33_ASAP7_75t_L g3769 ( 
.A1(n_3649),
.A2(n_2025),
.B(n_2030),
.C(n_2024),
.Y(n_3769)
);

INVx1_ASAP7_75t_SL g3770 ( 
.A(n_3711),
.Y(n_3770)
);

OAI21xp5_ASAP7_75t_SL g3771 ( 
.A1(n_3661),
.A2(n_2036),
.B(n_2034),
.Y(n_3771)
);

OAI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3644),
.A2(n_2049),
.B(n_1452),
.Y(n_3772)
);

A2O1A1Ixp33_ASAP7_75t_L g3773 ( 
.A1(n_3714),
.A2(n_1510),
.B(n_1514),
.C(n_1434),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3648),
.B(n_1688),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3646),
.Y(n_3775)
);

CKINVDCx20_ASAP7_75t_R g3776 ( 
.A(n_3666),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3651),
.Y(n_3777)
);

AO31x2_ASAP7_75t_L g3778 ( 
.A1(n_3700),
.A2(n_1637),
.A3(n_1638),
.B(n_1617),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3668),
.B(n_1691),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3687),
.Y(n_3780)
);

AO31x2_ASAP7_75t_L g3781 ( 
.A1(n_3691),
.A2(n_1707),
.A3(n_1766),
.B(n_1649),
.Y(n_3781)
);

OAI21x1_ASAP7_75t_L g3782 ( 
.A1(n_3656),
.A2(n_1782),
.B(n_1772),
.Y(n_3782)
);

AOI21xp5_ASAP7_75t_L g3783 ( 
.A1(n_3705),
.A2(n_1936),
.B(n_1929),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3670),
.B(n_1693),
.Y(n_3784)
);

HB1xp67_ASAP7_75t_L g3785 ( 
.A(n_3655),
.Y(n_3785)
);

AOI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_3673),
.A2(n_1938),
.B(n_1937),
.Y(n_3786)
);

O2A1O1Ixp33_ASAP7_75t_SL g3787 ( 
.A1(n_3688),
.A2(n_1882),
.B(n_1931),
.C(n_1836),
.Y(n_3787)
);

O2A1O1Ixp33_ASAP7_75t_SL g3788 ( 
.A1(n_3726),
.A2(n_2007),
.B(n_4),
.C(n_1),
.Y(n_3788)
);

OAI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_3701),
.A2(n_1945),
.B(n_1943),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_3727),
.B(n_1694),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3717),
.A2(n_1952),
.B(n_1946),
.Y(n_3791)
);

O2A1O1Ixp33_ASAP7_75t_SL g3792 ( 
.A1(n_3721),
.A2(n_6),
.B(n_2),
.C(n_5),
.Y(n_3792)
);

OAI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3706),
.A2(n_1706),
.B1(n_1708),
.B2(n_1703),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3679),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3697),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_3731),
.A2(n_1956),
.B(n_1953),
.Y(n_3796)
);

OAI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3683),
.A2(n_2836),
.B(n_2861),
.Y(n_3797)
);

OAI21xp33_ASAP7_75t_L g3798 ( 
.A1(n_3707),
.A2(n_1734),
.B(n_1729),
.Y(n_3798)
);

INVx2_ASAP7_75t_SL g3799 ( 
.A(n_3653),
.Y(n_3799)
);

O2A1O1Ixp33_ASAP7_75t_SL g3800 ( 
.A1(n_3704),
.A2(n_13),
.B(n_22),
.C(n_5),
.Y(n_3800)
);

AND2x4_ASAP7_75t_L g3801 ( 
.A(n_3676),
.B(n_982),
.Y(n_3801)
);

AO32x2_ASAP7_75t_L g3802 ( 
.A1(n_3659),
.A2(n_3658),
.A3(n_3708),
.B1(n_3715),
.B2(n_3689),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3695),
.A2(n_1963),
.B(n_1957),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_3706),
.A2(n_1972),
.B(n_1967),
.Y(n_3804)
);

NAND2xp33_ASAP7_75t_L g3805 ( 
.A(n_3660),
.B(n_1735),
.Y(n_3805)
);

O2A1O1Ixp33_ASAP7_75t_L g3806 ( 
.A1(n_3702),
.A2(n_1740),
.B(n_1748),
.C(n_1737),
.Y(n_3806)
);

O2A1O1Ixp33_ASAP7_75t_SL g3807 ( 
.A1(n_3654),
.A2(n_14),
.B(n_24),
.C(n_6),
.Y(n_3807)
);

AO31x2_ASAP7_75t_L g3808 ( 
.A1(n_3703),
.A2(n_9),
.A3(n_7),
.B(n_8),
.Y(n_3808)
);

NOR3xp33_ASAP7_75t_L g3809 ( 
.A(n_3722),
.B(n_1758),
.C(n_1757),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3775),
.Y(n_3810)
);

OAI222xp33_ASAP7_75t_L g3811 ( 
.A1(n_3761),
.A2(n_3663),
.B1(n_3674),
.B2(n_3712),
.C1(n_3675),
.C2(n_3680),
.Y(n_3811)
);

AO21x2_ASAP7_75t_L g3812 ( 
.A1(n_3748),
.A2(n_3663),
.B(n_3715),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3759),
.B(n_3676),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3760),
.B(n_3708),
.Y(n_3814)
);

OR2x2_ASAP7_75t_L g3815 ( 
.A(n_3785),
.B(n_3692),
.Y(n_3815)
);

AOI22xp33_ASAP7_75t_L g3816 ( 
.A1(n_3738),
.A2(n_3685),
.B1(n_3689),
.B2(n_3650),
.Y(n_3816)
);

AOI22xp33_ASAP7_75t_SL g3817 ( 
.A1(n_3772),
.A2(n_3682),
.B1(n_3657),
.B2(n_3642),
.Y(n_3817)
);

OAI22xp33_ASAP7_75t_L g3818 ( 
.A1(n_3770),
.A2(n_3660),
.B1(n_3681),
.B2(n_3678),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3777),
.Y(n_3819)
);

OAI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3742),
.A2(n_2055),
.B1(n_2057),
.B2(n_2050),
.Y(n_3820)
);

AND2x4_ASAP7_75t_SL g3821 ( 
.A(n_3758),
.B(n_2837),
.Y(n_3821)
);

AOI22xp33_ASAP7_75t_L g3822 ( 
.A1(n_3809),
.A2(n_1768),
.B1(n_1774),
.B2(n_1760),
.Y(n_3822)
);

CKINVDCx5p33_ASAP7_75t_R g3823 ( 
.A(n_3776),
.Y(n_3823)
);

NOR2x2_ASAP7_75t_L g3824 ( 
.A(n_3767),
.B(n_8),
.Y(n_3824)
);

CKINVDCx5p33_ASAP7_75t_R g3825 ( 
.A(n_3747),
.Y(n_3825)
);

AOI22xp33_ASAP7_75t_L g3826 ( 
.A1(n_3798),
.A2(n_1776),
.B1(n_1777),
.B2(n_1775),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3744),
.A2(n_1781),
.B1(n_1783),
.B2(n_1780),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3735),
.A2(n_1787),
.B1(n_1789),
.B2(n_1786),
.Y(n_3828)
);

OAI221xp5_ASAP7_75t_L g3829 ( 
.A1(n_3753),
.A2(n_1800),
.B1(n_1801),
.B2(n_1798),
.C(n_1793),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3780),
.B(n_3795),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3740),
.Y(n_3831)
);

INVx4_ASAP7_75t_L g3832 ( 
.A(n_3762),
.Y(n_3832)
);

INVx4_ASAP7_75t_L g3833 ( 
.A(n_3762),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3794),
.Y(n_3834)
);

AOI22xp33_ASAP7_75t_L g3835 ( 
.A1(n_3796),
.A2(n_1807),
.B1(n_1814),
.B2(n_1806),
.Y(n_3835)
);

INVx2_ASAP7_75t_SL g3836 ( 
.A(n_3741),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3745),
.B(n_1816),
.Y(n_3837)
);

OAI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3756),
.A2(n_3734),
.B1(n_3746),
.B2(n_3773),
.Y(n_3838)
);

NOR2xp33_ASAP7_75t_SL g3839 ( 
.A(n_3754),
.B(n_2068),
.Y(n_3839)
);

AOI22xp33_ASAP7_75t_L g3840 ( 
.A1(n_3790),
.A2(n_1824),
.B1(n_1827),
.B2(n_1823),
.Y(n_3840)
);

O2A1O1Ixp33_ASAP7_75t_L g3841 ( 
.A1(n_3788),
.A2(n_1835),
.B(n_1841),
.C(n_1834),
.Y(n_3841)
);

AOI22xp33_ASAP7_75t_L g3842 ( 
.A1(n_3786),
.A2(n_1844),
.B1(n_1847),
.B2(n_1843),
.Y(n_3842)
);

OR2x2_ASAP7_75t_L g3843 ( 
.A(n_3778),
.B(n_9),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3799),
.B(n_983),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3778),
.Y(n_3845)
);

AOI22xp33_ASAP7_75t_L g3846 ( 
.A1(n_3768),
.A2(n_1851),
.B1(n_1854),
.B2(n_1849),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3774),
.B(n_1858),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3781),
.Y(n_3848)
);

NAND2x1_ASAP7_75t_L g3849 ( 
.A(n_3755),
.B(n_2837),
.Y(n_3849)
);

OAI21x1_ASAP7_75t_L g3850 ( 
.A1(n_3737),
.A2(n_987),
.B(n_985),
.Y(n_3850)
);

AOI22xp33_ASAP7_75t_L g3851 ( 
.A1(n_3783),
.A2(n_1862),
.B1(n_1864),
.B2(n_1861),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3739),
.A2(n_1868),
.B(n_1866),
.Y(n_3852)
);

AOI22xp33_ASAP7_75t_SL g3853 ( 
.A1(n_3789),
.A2(n_1873),
.B1(n_1875),
.B2(n_1871),
.Y(n_3853)
);

AOI22xp33_ASAP7_75t_L g3854 ( 
.A1(n_3779),
.A2(n_1879),
.B1(n_1880),
.B2(n_1877),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3802),
.B(n_3749),
.Y(n_3855)
);

NOR2xp33_ASAP7_75t_L g3856 ( 
.A(n_3757),
.B(n_1881),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3749),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3791),
.A2(n_1885),
.B1(n_1892),
.B2(n_1883),
.Y(n_3858)
);

OAI22xp33_ASAP7_75t_L g3859 ( 
.A1(n_3802),
.A2(n_2075),
.B1(n_1894),
.B2(n_1895),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3781),
.Y(n_3860)
);

OAI22xp33_ASAP7_75t_L g3861 ( 
.A1(n_3771),
.A2(n_2041),
.B1(n_2042),
.B2(n_2039),
.Y(n_3861)
);

A2O1A1Ixp33_ASAP7_75t_L g3862 ( 
.A1(n_3806),
.A2(n_2044),
.B(n_2046),
.C(n_2043),
.Y(n_3862)
);

AOI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3752),
.A2(n_1902),
.B1(n_1903),
.B2(n_1893),
.Y(n_3863)
);

OAI22xp5_ASAP7_75t_L g3864 ( 
.A1(n_3766),
.A2(n_1910),
.B1(n_1912),
.B2(n_1904),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_3764),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3765),
.Y(n_3866)
);

A2O1A1Ixp33_ASAP7_75t_L g3867 ( 
.A1(n_3763),
.A2(n_2065),
.B(n_1918),
.C(n_1968),
.Y(n_3867)
);

OAI211xp5_ASAP7_75t_SL g3868 ( 
.A1(n_3769),
.A2(n_1920),
.B(n_1921),
.C(n_1917),
.Y(n_3868)
);

CKINVDCx5p33_ASAP7_75t_R g3869 ( 
.A(n_3801),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3808),
.Y(n_3870)
);

HB1xp67_ASAP7_75t_L g3871 ( 
.A(n_3782),
.Y(n_3871)
);

BUFx6f_ASAP7_75t_L g3872 ( 
.A(n_3797),
.Y(n_3872)
);

OAI22xp5_ASAP7_75t_L g3873 ( 
.A1(n_3751),
.A2(n_1926),
.B1(n_1928),
.B2(n_1923),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3743),
.Y(n_3874)
);

A2O1A1Ixp33_ASAP7_75t_L g3875 ( 
.A1(n_3750),
.A2(n_2047),
.B(n_2048),
.C(n_2035),
.Y(n_3875)
);

OAI22xp33_ASAP7_75t_L g3876 ( 
.A1(n_3784),
.A2(n_2061),
.B1(n_2059),
.B2(n_1947),
.Y(n_3876)
);

AOI22xp5_ASAP7_75t_L g3877 ( 
.A1(n_3787),
.A2(n_1949),
.B1(n_1951),
.B2(n_1930),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3808),
.B(n_10),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3743),
.Y(n_3879)
);

BUFx2_ASAP7_75t_L g3880 ( 
.A(n_3736),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3792),
.B(n_3800),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3736),
.Y(n_3882)
);

OAI21xp33_ASAP7_75t_L g3883 ( 
.A1(n_3793),
.A2(n_1955),
.B(n_1954),
.Y(n_3883)
);

AND2x4_ASAP7_75t_L g3884 ( 
.A(n_3804),
.B(n_11),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3803),
.B(n_12),
.Y(n_3885)
);

BUFx2_ASAP7_75t_L g3886 ( 
.A(n_3805),
.Y(n_3886)
);

INVx3_ASAP7_75t_L g3887 ( 
.A(n_3807),
.Y(n_3887)
);

AOI22xp33_ASAP7_75t_L g3888 ( 
.A1(n_3738),
.A2(n_1961),
.B1(n_1962),
.B2(n_1959),
.Y(n_3888)
);

INVxp67_ASAP7_75t_SL g3889 ( 
.A(n_3813),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3810),
.Y(n_3890)
);

AOI22xp33_ASAP7_75t_L g3891 ( 
.A1(n_3880),
.A2(n_2029),
.B1(n_2023),
.B2(n_1977),
.Y(n_3891)
);

INVx1_ASAP7_75t_SL g3892 ( 
.A(n_3815),
.Y(n_3892)
);

AOI22xp33_ASAP7_75t_SL g3893 ( 
.A1(n_3838),
.A2(n_1979),
.B1(n_1980),
.B2(n_1965),
.Y(n_3893)
);

OA21x2_ASAP7_75t_L g3894 ( 
.A1(n_3855),
.A2(n_1986),
.B(n_1982),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3819),
.Y(n_3895)
);

HB1xp67_ASAP7_75t_L g3896 ( 
.A(n_3830),
.Y(n_3896)
);

HB1xp67_ASAP7_75t_L g3897 ( 
.A(n_3831),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3834),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_3837),
.B(n_1987),
.Y(n_3899)
);

INVx3_ASAP7_75t_L g3900 ( 
.A(n_3832),
.Y(n_3900)
);

BUFx2_ASAP7_75t_L g3901 ( 
.A(n_3814),
.Y(n_3901)
);

INVxp67_ASAP7_75t_L g3902 ( 
.A(n_3836),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3833),
.B(n_12),
.Y(n_3903)
);

INVx1_ASAP7_75t_SL g3904 ( 
.A(n_3823),
.Y(n_3904)
);

OAI21x1_ASAP7_75t_L g3905 ( 
.A1(n_3848),
.A2(n_13),
.B(n_15),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3870),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3816),
.B(n_3812),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3857),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3845),
.Y(n_3909)
);

AO31x2_ASAP7_75t_L g3910 ( 
.A1(n_3882),
.A2(n_17),
.A3(n_15),
.B(n_16),
.Y(n_3910)
);

OAI21x1_ASAP7_75t_L g3911 ( 
.A1(n_3860),
.A2(n_16),
.B(n_17),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3879),
.Y(n_3912)
);

INVx3_ASAP7_75t_L g3913 ( 
.A(n_3821),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3874),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3865),
.B(n_1993),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3866),
.Y(n_3916)
);

BUFx2_ASAP7_75t_L g3917 ( 
.A(n_3869),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3871),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3872),
.Y(n_3919)
);

HB1xp67_ASAP7_75t_L g3920 ( 
.A(n_3843),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3872),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3878),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3859),
.B(n_1994),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3872),
.Y(n_3924)
);

INVx3_ASAP7_75t_L g3925 ( 
.A(n_3849),
.Y(n_3925)
);

INVxp67_ASAP7_75t_SL g3926 ( 
.A(n_3887),
.Y(n_3926)
);

INVxp67_ASAP7_75t_L g3927 ( 
.A(n_3847),
.Y(n_3927)
);

OAI21x1_ASAP7_75t_L g3928 ( 
.A1(n_3850),
.A2(n_19),
.B(n_20),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3881),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3818),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3885),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3884),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3884),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3844),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3886),
.B(n_19),
.Y(n_3935)
);

OAI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3852),
.A2(n_1999),
.B(n_1996),
.Y(n_3936)
);

INVx2_ASAP7_75t_SL g3937 ( 
.A(n_3825),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3817),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3824),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3841),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3820),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3856),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3877),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3888),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3876),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3827),
.Y(n_3946)
);

OAI21x1_ASAP7_75t_L g3947 ( 
.A1(n_3811),
.A2(n_20),
.B(n_21),
.Y(n_3947)
);

BUFx6f_ASAP7_75t_L g3948 ( 
.A(n_3839),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3862),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3854),
.B(n_21),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3829),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3873),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3864),
.Y(n_3953)
);

INVx1_ASAP7_75t_SL g3954 ( 
.A(n_3853),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3828),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3875),
.Y(n_3956)
);

HB1xp67_ASAP7_75t_L g3957 ( 
.A(n_3920),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3912),
.Y(n_3958)
);

BUFx2_ASAP7_75t_L g3959 ( 
.A(n_3926),
.Y(n_3959)
);

A2O1A1Ixp33_ASAP7_75t_L g3960 ( 
.A1(n_3940),
.A2(n_3883),
.B(n_3867),
.C(n_3840),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3901),
.B(n_3835),
.Y(n_3961)
);

OA21x2_ASAP7_75t_L g3962 ( 
.A1(n_3906),
.A2(n_3908),
.B(n_3914),
.Y(n_3962)
);

AOI22xp33_ASAP7_75t_SL g3963 ( 
.A1(n_3894),
.A2(n_2004),
.B1(n_2009),
.B2(n_2003),
.Y(n_3963)
);

HB1xp67_ASAP7_75t_L g3964 ( 
.A(n_3918),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3892),
.B(n_3842),
.Y(n_3965)
);

AND2x4_ASAP7_75t_L g3966 ( 
.A(n_3933),
.B(n_3851),
.Y(n_3966)
);

AOI22xp33_ASAP7_75t_L g3967 ( 
.A1(n_3951),
.A2(n_3868),
.B1(n_3863),
.B2(n_3846),
.Y(n_3967)
);

AOI22xp33_ASAP7_75t_L g3968 ( 
.A1(n_3893),
.A2(n_3861),
.B1(n_3858),
.B2(n_3826),
.Y(n_3968)
);

AOI221xp5_ASAP7_75t_L g3969 ( 
.A1(n_3891),
.A2(n_3822),
.B1(n_2015),
.B2(n_2017),
.C(n_2013),
.Y(n_3969)
);

OAI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3929),
.A2(n_2019),
.B1(n_2011),
.B2(n_1981),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3922),
.B(n_23),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3932),
.Y(n_3972)
);

OAI22xp5_ASAP7_75t_L g3973 ( 
.A1(n_3938),
.A2(n_1984),
.B1(n_2001),
.B2(n_1978),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3890),
.Y(n_3974)
);

OAI211xp5_ASAP7_75t_SL g3975 ( 
.A1(n_3941),
.A2(n_3954),
.B(n_3923),
.C(n_3943),
.Y(n_3975)
);

AOI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_3936),
.A2(n_2008),
.B(n_2006),
.Y(n_3976)
);

OA21x2_ASAP7_75t_L g3977 ( 
.A1(n_3909),
.A2(n_2021),
.B(n_2012),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3889),
.B(n_23),
.Y(n_3978)
);

OAI22xp33_ASAP7_75t_L g3979 ( 
.A1(n_3930),
.A2(n_2031),
.B1(n_2033),
.B2(n_2026),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3944),
.A2(n_2045),
.B1(n_2053),
.B2(n_2038),
.Y(n_3980)
);

BUFx3_ASAP7_75t_L g3981 ( 
.A(n_3917),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_3931),
.B(n_24),
.Y(n_3982)
);

CKINVDCx5p33_ASAP7_75t_R g3983 ( 
.A(n_3904),
.Y(n_3983)
);

AOI33xp33_ASAP7_75t_L g3984 ( 
.A1(n_3946),
.A2(n_28),
.A3(n_30),
.B1(n_26),
.B2(n_27),
.B3(n_29),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3895),
.Y(n_3985)
);

BUFx3_ASAP7_75t_L g3986 ( 
.A(n_3937),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_SL g3987 ( 
.A1(n_3939),
.A2(n_2066),
.B1(n_2063),
.B2(n_32),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3898),
.Y(n_3988)
);

OAI22xp5_ASAP7_75t_L g3989 ( 
.A1(n_3949),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_3989)
);

AOI22xp33_ASAP7_75t_L g3990 ( 
.A1(n_3907),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_3990)
);

HB1xp67_ASAP7_75t_L g3991 ( 
.A(n_3896),
.Y(n_3991)
);

OAI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3945),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_3992)
);

AOI22xp33_ASAP7_75t_L g3993 ( 
.A1(n_3956),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_3993)
);

AOI22xp33_ASAP7_75t_L g3994 ( 
.A1(n_3952),
.A2(n_41),
.B1(n_37),
.B2(n_40),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_L g3995 ( 
.A1(n_3953),
.A2(n_3955),
.B1(n_3942),
.B2(n_3950),
.Y(n_3995)
);

OAI22xp5_ASAP7_75t_L g3996 ( 
.A1(n_3902),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3897),
.B(n_43),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3916),
.Y(n_3998)
);

OAI22xp5_ASAP7_75t_L g3999 ( 
.A1(n_3927),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3999)
);

AOI22xp33_ASAP7_75t_L g4000 ( 
.A1(n_3899),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_4000)
);

AOI22xp33_ASAP7_75t_SL g4001 ( 
.A1(n_3947),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_4001)
);

OAI22xp5_ASAP7_75t_L g4002 ( 
.A1(n_3934),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_4002)
);

AOI22xp33_ASAP7_75t_L g4003 ( 
.A1(n_3948),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_4003)
);

INVx2_ASAP7_75t_SL g4004 ( 
.A(n_3900),
.Y(n_4004)
);

OAI221xp5_ASAP7_75t_L g4005 ( 
.A1(n_3915),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.C(n_57),
.Y(n_4005)
);

NAND2xp33_ASAP7_75t_L g4006 ( 
.A(n_3948),
.B(n_54),
.Y(n_4006)
);

OAI21xp5_ASAP7_75t_L g4007 ( 
.A1(n_3928),
.A2(n_56),
.B(n_57),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3919),
.B(n_58),
.Y(n_4008)
);

INVx4_ASAP7_75t_L g4009 ( 
.A(n_3913),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3925),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_4010)
);

OAI221xp5_ASAP7_75t_L g4011 ( 
.A1(n_3921),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.C(n_63),
.Y(n_4011)
);

AOI22xp33_ASAP7_75t_L g4012 ( 
.A1(n_3935),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_4012)
);

AOI221x1_ASAP7_75t_SL g4013 ( 
.A1(n_3910),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_4013)
);

CKINVDCx5p33_ASAP7_75t_R g4014 ( 
.A(n_3903),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3924),
.Y(n_4015)
);

AOI22xp33_ASAP7_75t_L g4016 ( 
.A1(n_3911),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_4016)
);

A2O1A1Ixp33_ASAP7_75t_L g4017 ( 
.A1(n_3905),
.A2(n_78),
.B(n_86),
.C(n_69),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3910),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3933),
.Y(n_4019)
);

OAI22xp33_ASAP7_75t_L g4020 ( 
.A1(n_3938),
.A2(n_74),
.B1(n_71),
.B2(n_73),
.Y(n_4020)
);

OAI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_3891),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_4021)
);

OAI211xp5_ASAP7_75t_L g4022 ( 
.A1(n_3893),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3889),
.B(n_76),
.Y(n_4023)
);

AO21x2_ASAP7_75t_L g4024 ( 
.A1(n_3912),
.A2(n_77),
.B(n_79),
.Y(n_4024)
);

OAI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3938),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_4025)
);

OAI211xp5_ASAP7_75t_SL g4026 ( 
.A1(n_3893),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_4026)
);

OAI21x1_ASAP7_75t_L g4027 ( 
.A1(n_3906),
.A2(n_83),
.B(n_84),
.Y(n_4027)
);

OR2x2_ASAP7_75t_L g4028 ( 
.A(n_3896),
.B(n_85),
.Y(n_4028)
);

BUFx6f_ASAP7_75t_L g4029 ( 
.A(n_3948),
.Y(n_4029)
);

OAI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_3893),
.A2(n_85),
.B(n_86),
.Y(n_4030)
);

A2O1A1Ixp33_ASAP7_75t_L g4031 ( 
.A1(n_3940),
.A2(n_96),
.B(n_108),
.C(n_87),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3951),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_4032)
);

OAI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3891),
.A2(n_91),
.B1(n_88),
.B2(n_90),
.Y(n_4033)
);

BUFx10_ASAP7_75t_L g4034 ( 
.A(n_3948),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3912),
.Y(n_4035)
);

AOI222xp33_ASAP7_75t_L g4036 ( 
.A1(n_3940),
.A2(n_93),
.B1(n_95),
.B2(n_91),
.C1(n_92),
.C2(n_94),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3901),
.B(n_92),
.Y(n_4037)
);

OAI22xp5_ASAP7_75t_SL g4038 ( 
.A1(n_3939),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_4038)
);

BUFx12f_ASAP7_75t_L g4039 ( 
.A(n_3948),
.Y(n_4039)
);

AOI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3951),
.A2(n_102),
.B1(n_98),
.B2(n_101),
.Y(n_4040)
);

BUFx2_ASAP7_75t_L g4041 ( 
.A(n_3926),
.Y(n_4041)
);

BUFx3_ASAP7_75t_L g4042 ( 
.A(n_3917),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3912),
.Y(n_4043)
);

AOI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_3940),
.A2(n_98),
.B(n_103),
.Y(n_4044)
);

OAI22xp33_ASAP7_75t_L g4045 ( 
.A1(n_3938),
.A2(n_108),
.B1(n_105),
.B2(n_106),
.Y(n_4045)
);

HB1xp67_ASAP7_75t_L g4046 ( 
.A(n_3920),
.Y(n_4046)
);

OAI221xp5_ASAP7_75t_L g4047 ( 
.A1(n_3893),
.A2(n_110),
.B1(n_106),
.B2(n_109),
.C(n_111),
.Y(n_4047)
);

AOI221xp5_ASAP7_75t_L g4048 ( 
.A1(n_3940),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.C(n_112),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3912),
.Y(n_4049)
);

HB1xp67_ASAP7_75t_L g4050 ( 
.A(n_3920),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3889),
.B(n_112),
.Y(n_4051)
);

OAI211xp5_ASAP7_75t_L g4052 ( 
.A1(n_3893),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_4052)
);

OAI22xp5_ASAP7_75t_L g4053 ( 
.A1(n_3891),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_4053)
);

INVx2_ASAP7_75t_L g4054 ( 
.A(n_3933),
.Y(n_4054)
);

OAI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3893),
.A2(n_116),
.B(n_117),
.Y(n_4055)
);

AOI22xp33_ASAP7_75t_L g4056 ( 
.A1(n_3951),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3912),
.Y(n_4057)
);

AND2x4_ASAP7_75t_L g4058 ( 
.A(n_3933),
.B(n_119),
.Y(n_4058)
);

AOI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3951),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_L g4060 ( 
.A1(n_3951),
.A2(n_127),
.B1(n_124),
.B2(n_126),
.Y(n_4060)
);

OAI22xp5_ASAP7_75t_L g4061 ( 
.A1(n_3891),
.A2(n_128),
.B1(n_124),
.B2(n_126),
.Y(n_4061)
);

OAI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3891),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_4062)
);

OAI22xp5_ASAP7_75t_L g4063 ( 
.A1(n_3891),
.A2(n_132),
.B1(n_129),
.B2(n_130),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_L g4064 ( 
.A1(n_3951),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_4064)
);

AO31x2_ASAP7_75t_L g4065 ( 
.A1(n_3906),
.A2(n_137),
.A3(n_133),
.B(n_136),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3933),
.Y(n_4066)
);

AOI21xp33_ASAP7_75t_L g4067 ( 
.A1(n_3940),
.A2(n_137),
.B(n_138),
.Y(n_4067)
);

OR2x6_ASAP7_75t_L g4068 ( 
.A(n_3917),
.B(n_138),
.Y(n_4068)
);

OAI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_3891),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_4069)
);

CKINVDCx20_ASAP7_75t_R g4070 ( 
.A(n_3937),
.Y(n_4070)
);

HB1xp67_ASAP7_75t_L g4071 ( 
.A(n_3920),
.Y(n_4071)
);

AOI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_3951),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_4072)
);

OAI21x1_ASAP7_75t_L g4073 ( 
.A1(n_3906),
.A2(n_142),
.B(n_143),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_3957),
.B(n_143),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3962),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3958),
.Y(n_4076)
);

AND2x4_ASAP7_75t_L g4077 ( 
.A(n_4004),
.B(n_144),
.Y(n_4077)
);

OR2x2_ASAP7_75t_L g4078 ( 
.A(n_4046),
.B(n_145),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_4035),
.Y(n_4079)
);

AND2x2_ASAP7_75t_L g4080 ( 
.A(n_3959),
.B(n_145),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_4041),
.B(n_146),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_3991),
.B(n_146),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_4043),
.Y(n_4083)
);

AO31x2_ASAP7_75t_L g4084 ( 
.A1(n_3978),
.A2(n_149),
.A3(n_147),
.B(n_148),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_4019),
.B(n_147),
.Y(n_4085)
);

HB1xp67_ASAP7_75t_L g4086 ( 
.A(n_4050),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_4049),
.Y(n_4087)
);

AOI21xp5_ASAP7_75t_L g4088 ( 
.A1(n_4044),
.A2(n_149),
.B(n_150),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_4057),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3974),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3988),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4071),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3998),
.Y(n_4093)
);

BUFx2_ASAP7_75t_L g4094 ( 
.A(n_3981),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_3962),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3995),
.B(n_4023),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_4054),
.B(n_151),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3964),
.Y(n_4098)
);

OR2x2_ASAP7_75t_L g4099 ( 
.A(n_3972),
.B(n_4066),
.Y(n_4099)
);

OR2x2_ASAP7_75t_L g4100 ( 
.A(n_3985),
.B(n_152),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_4065),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4065),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_4009),
.B(n_153),
.Y(n_4103)
);

HB1xp67_ASAP7_75t_L g4104 ( 
.A(n_4015),
.Y(n_4104)
);

INVx2_ASAP7_75t_SL g4105 ( 
.A(n_4042),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3961),
.B(n_153),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_3965),
.B(n_3997),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_3966),
.B(n_154),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_4028),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_4051),
.B(n_154),
.Y(n_4110)
);

AND2x4_ASAP7_75t_L g4111 ( 
.A(n_3986),
.B(n_155),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_4008),
.Y(n_4112)
);

OR2x2_ASAP7_75t_L g4113 ( 
.A(n_3982),
.B(n_155),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_3971),
.B(n_156),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_4058),
.Y(n_4115)
);

INVxp67_ASAP7_75t_L g4116 ( 
.A(n_4068),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_4034),
.Y(n_4117)
);

NAND3xp33_ASAP7_75t_L g4118 ( 
.A(n_3963),
.B(n_156),
.C(n_157),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4024),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_4027),
.Y(n_4120)
);

AND2x4_ASAP7_75t_L g4121 ( 
.A(n_4037),
.B(n_158),
.Y(n_4121)
);

AND2x4_ASAP7_75t_L g4122 ( 
.A(n_4070),
.B(n_158),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4073),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3977),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_4014),
.B(n_159),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_4029),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_4068),
.B(n_160),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3977),
.Y(n_4128)
);

HB1xp67_ASAP7_75t_L g4129 ( 
.A(n_4007),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_4029),
.B(n_160),
.Y(n_4130)
);

AND2x4_ASAP7_75t_L g4131 ( 
.A(n_3983),
.B(n_162),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3975),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_4039),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_4013),
.B(n_162),
.Y(n_4134)
);

NOR2xp33_ASAP7_75t_L g4135 ( 
.A(n_3987),
.B(n_163),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_4002),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_4038),
.Y(n_4137)
);

BUFx2_ASAP7_75t_L g4138 ( 
.A(n_4017),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3990),
.B(n_163),
.Y(n_4139)
);

INVx3_ASAP7_75t_L g4140 ( 
.A(n_4006),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4018),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_4001),
.B(n_164),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_4072),
.Y(n_4143)
);

AND2x2_ASAP7_75t_L g4144 ( 
.A(n_4016),
.B(n_164),
.Y(n_4144)
);

BUFx3_ASAP7_75t_L g4145 ( 
.A(n_4005),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3984),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_4012),
.B(n_3967),
.Y(n_4147)
);

INVxp67_ASAP7_75t_SL g4148 ( 
.A(n_4020),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_4011),
.Y(n_4149)
);

BUFx3_ASAP7_75t_L g4150 ( 
.A(n_3996),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4067),
.B(n_165),
.Y(n_4151)
);

OR2x2_ASAP7_75t_L g4152 ( 
.A(n_3992),
.B(n_167),
.Y(n_4152)
);

INVxp67_ASAP7_75t_L g4153 ( 
.A(n_3999),
.Y(n_4153)
);

AND2x2_ASAP7_75t_L g4154 ( 
.A(n_3960),
.B(n_167),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4025),
.B(n_168),
.Y(n_4155)
);

HB1xp67_ASAP7_75t_L g4156 ( 
.A(n_4010),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_3973),
.B(n_169),
.Y(n_4157)
);

NAND3xp33_ASAP7_75t_L g4158 ( 
.A(n_4048),
.B(n_169),
.C(n_170),
.Y(n_4158)
);

INVx1_ASAP7_75t_SL g4159 ( 
.A(n_3989),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_4036),
.B(n_4031),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4032),
.B(n_170),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4045),
.B(n_171),
.Y(n_4162)
);

OR2x2_ASAP7_75t_L g4163 ( 
.A(n_4040),
.B(n_172),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3970),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4021),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4033),
.Y(n_4166)
);

OR2x2_ASAP7_75t_L g4167 ( 
.A(n_4056),
.B(n_172),
.Y(n_4167)
);

AND2x4_ASAP7_75t_L g4168 ( 
.A(n_4030),
.B(n_174),
.Y(n_4168)
);

BUFx2_ASAP7_75t_L g4169 ( 
.A(n_4055),
.Y(n_4169)
);

BUFx3_ASAP7_75t_L g4170 ( 
.A(n_4047),
.Y(n_4170)
);

AND2x2_ASAP7_75t_L g4171 ( 
.A(n_4059),
.B(n_174),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_4053),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4061),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4060),
.B(n_175),
.Y(n_4174)
);

OR2x2_ASAP7_75t_L g4175 ( 
.A(n_4064),
.B(n_175),
.Y(n_4175)
);

AO21x2_ASAP7_75t_L g4176 ( 
.A1(n_3979),
.A2(n_177),
.B(n_178),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_4026),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4062),
.Y(n_4178)
);

OR2x2_ASAP7_75t_L g4179 ( 
.A(n_3994),
.B(n_3993),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4063),
.Y(n_4180)
);

INVxp67_ASAP7_75t_SL g4181 ( 
.A(n_4003),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_4000),
.B(n_179),
.Y(n_4182)
);

BUFx3_ASAP7_75t_L g4183 ( 
.A(n_4069),
.Y(n_4183)
);

HB1xp67_ASAP7_75t_L g4184 ( 
.A(n_4022),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4052),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_3980),
.Y(n_4186)
);

INVx2_ASAP7_75t_L g4187 ( 
.A(n_3968),
.Y(n_4187)
);

AND2x4_ASAP7_75t_L g4188 ( 
.A(n_3976),
.B(n_180),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_3969),
.Y(n_4189)
);

INVx2_ASAP7_75t_SL g4190 ( 
.A(n_3981),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_3959),
.B(n_180),
.Y(n_4191)
);

INVxp67_ASAP7_75t_L g4192 ( 
.A(n_3957),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_3959),
.B(n_181),
.Y(n_4193)
);

INVx5_ASAP7_75t_L g4194 ( 
.A(n_4068),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_3959),
.B(n_182),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3959),
.B(n_182),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_3957),
.B(n_183),
.Y(n_4197)
);

BUFx6f_ASAP7_75t_L g4198 ( 
.A(n_4039),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_3962),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_3959),
.B(n_184),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_3959),
.B(n_184),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_3959),
.B(n_185),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_3958),
.Y(n_4203)
);

AOI22xp33_ASAP7_75t_L g4204 ( 
.A1(n_3975),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_3959),
.B(n_186),
.Y(n_4205)
);

HB1xp67_ASAP7_75t_L g4206 ( 
.A(n_3957),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3958),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_3959),
.B(n_187),
.Y(n_4208)
);

NAND4xp25_ASAP7_75t_L g4209 ( 
.A(n_4013),
.B(n_190),
.C(n_188),
.D(n_189),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3958),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_3959),
.B(n_190),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_3959),
.B(n_191),
.Y(n_4212)
);

AND2x2_ASAP7_75t_L g4213 ( 
.A(n_3959),
.B(n_191),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_3959),
.B(n_193),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_3959),
.B(n_193),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_3962),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3958),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_3959),
.B(n_194),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3958),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3958),
.Y(n_4220)
);

BUFx6f_ASAP7_75t_L g4221 ( 
.A(n_4039),
.Y(n_4221)
);

BUFx2_ASAP7_75t_L g4222 ( 
.A(n_3959),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_3959),
.B(n_194),
.Y(n_4223)
);

OAI31xp33_ASAP7_75t_SL g4224 ( 
.A1(n_3975),
.A2(n_198),
.A3(n_195),
.B(n_196),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3962),
.Y(n_4225)
);

INVx2_ASAP7_75t_L g4226 ( 
.A(n_3962),
.Y(n_4226)
);

INVx3_ASAP7_75t_L g4227 ( 
.A(n_3981),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_3962),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_3959),
.B(n_196),
.Y(n_4229)
);

HB1xp67_ASAP7_75t_L g4230 ( 
.A(n_3957),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3958),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_3958),
.Y(n_4232)
);

OR2x2_ASAP7_75t_L g4233 ( 
.A(n_3957),
.B(n_199),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_3962),
.Y(n_4234)
);

INVx2_ASAP7_75t_SL g4235 ( 
.A(n_4198),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4076),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4079),
.Y(n_4237)
);

AOI22xp33_ASAP7_75t_L g4238 ( 
.A1(n_4145),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4083),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4094),
.Y(n_4240)
);

OAI21xp5_ASAP7_75t_L g4241 ( 
.A1(n_4160),
.A2(n_201),
.B(n_204),
.Y(n_4241)
);

AOI222xp33_ASAP7_75t_L g4242 ( 
.A1(n_4169),
.A2(n_207),
.B1(n_209),
.B2(n_204),
.C1(n_205),
.C2(n_208),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_4117),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4227),
.Y(n_4244)
);

OAI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_4129),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4132),
.B(n_4107),
.Y(n_4246)
);

INVx2_ASAP7_75t_L g4247 ( 
.A(n_4105),
.Y(n_4247)
);

AOI22xp33_ASAP7_75t_L g4248 ( 
.A1(n_4170),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_4248)
);

HB1xp67_ASAP7_75t_L g4249 ( 
.A(n_4086),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4190),
.Y(n_4250)
);

BUFx2_ASAP7_75t_L g4251 ( 
.A(n_4222),
.Y(n_4251)
);

HB1xp67_ASAP7_75t_L g4252 ( 
.A(n_4206),
.Y(n_4252)
);

AOI33xp33_ASAP7_75t_L g4253 ( 
.A1(n_4146),
.A2(n_213),
.A3(n_215),
.B1(n_210),
.B2(n_211),
.B3(n_214),
.Y(n_4253)
);

HB1xp67_ASAP7_75t_L g4254 ( 
.A(n_4230),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_4133),
.Y(n_4255)
);

NAND3xp33_ASAP7_75t_L g4256 ( 
.A(n_4224),
.B(n_213),
.C(n_214),
.Y(n_4256)
);

INVxp67_ASAP7_75t_L g4257 ( 
.A(n_4184),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4087),
.Y(n_4258)
);

INVx3_ASAP7_75t_L g4259 ( 
.A(n_4198),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4126),
.B(n_216),
.Y(n_4260)
);

NOR2xp33_ASAP7_75t_L g4261 ( 
.A(n_4221),
.B(n_216),
.Y(n_4261)
);

AOI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_4138),
.A2(n_220),
.B1(n_217),
.B2(n_219),
.Y(n_4262)
);

INVx5_ASAP7_75t_L g4263 ( 
.A(n_4221),
.Y(n_4263)
);

OAI22xp5_ASAP7_75t_L g4264 ( 
.A1(n_4148),
.A2(n_222),
.B1(n_219),
.B2(n_221),
.Y(n_4264)
);

OAI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_4158),
.A2(n_221),
.B(n_223),
.Y(n_4265)
);

INVx2_ASAP7_75t_SL g4266 ( 
.A(n_4194),
.Y(n_4266)
);

NOR2xp33_ASAP7_75t_L g4267 ( 
.A(n_4116),
.B(n_224),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4089),
.Y(n_4268)
);

BUFx2_ASAP7_75t_L g4269 ( 
.A(n_4194),
.Y(n_4269)
);

AOI22xp5_ASAP7_75t_L g4270 ( 
.A1(n_4209),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_4270)
);

AOI31xp33_ASAP7_75t_L g4271 ( 
.A1(n_4154),
.A2(n_229),
.A3(n_225),
.B(n_228),
.Y(n_4271)
);

NOR2x1_ASAP7_75t_L g4272 ( 
.A(n_4119),
.B(n_229),
.Y(n_4272)
);

INVxp67_ASAP7_75t_SL g4273 ( 
.A(n_4140),
.Y(n_4273)
);

OR2x2_ASAP7_75t_L g4274 ( 
.A(n_4092),
.B(n_230),
.Y(n_4274)
);

AOI22xp33_ASAP7_75t_L g4275 ( 
.A1(n_4183),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_4275)
);

AOI221xp5_ASAP7_75t_L g4276 ( 
.A1(n_4147),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.C(n_236),
.Y(n_4276)
);

BUFx3_ASAP7_75t_L g4277 ( 
.A(n_4131),
.Y(n_4277)
);

AO21x2_ASAP7_75t_L g4278 ( 
.A1(n_4074),
.A2(n_233),
.B(n_236),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4090),
.Y(n_4279)
);

AO21x2_ASAP7_75t_L g4280 ( 
.A1(n_4075),
.A2(n_237),
.B(n_239),
.Y(n_4280)
);

NAND4xp25_ASAP7_75t_L g4281 ( 
.A(n_4135),
.B(n_241),
.C(n_242),
.D(n_240),
.Y(n_4281)
);

AOI21xp33_ASAP7_75t_SL g4282 ( 
.A1(n_4137),
.A2(n_237),
.B(n_240),
.Y(n_4282)
);

OAI22xp5_ASAP7_75t_L g4283 ( 
.A1(n_4156),
.A2(n_244),
.B1(n_241),
.B2(n_243),
.Y(n_4283)
);

AO21x2_ASAP7_75t_L g4284 ( 
.A1(n_4095),
.A2(n_243),
.B(n_244),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4091),
.Y(n_4285)
);

BUFx3_ASAP7_75t_L g4286 ( 
.A(n_4111),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4093),
.Y(n_4287)
);

INVxp67_ASAP7_75t_SL g4288 ( 
.A(n_4192),
.Y(n_4288)
);

NOR2xp33_ASAP7_75t_L g4289 ( 
.A(n_4187),
.B(n_245),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4203),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4112),
.B(n_246),
.Y(n_4291)
);

OAI221xp5_ASAP7_75t_L g4292 ( 
.A1(n_4096),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.C(n_249),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4207),
.Y(n_4293)
);

OAI221xp5_ASAP7_75t_L g4294 ( 
.A1(n_4141),
.A2(n_4181),
.B1(n_4134),
.B2(n_4124),
.C(n_4128),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_4099),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4210),
.Y(n_4296)
);

AOI221xp5_ASAP7_75t_L g4297 ( 
.A1(n_4153),
.A2(n_4159),
.B1(n_4185),
.B2(n_4149),
.C(n_4166),
.Y(n_4297)
);

NAND5xp2_ASAP7_75t_SL g4298 ( 
.A(n_4204),
.B(n_252),
.C(n_250),
.D(n_251),
.E(n_253),
.Y(n_4298)
);

INVxp67_ASAP7_75t_L g4299 ( 
.A(n_4120),
.Y(n_4299)
);

OAI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_4088),
.A2(n_4162),
.B(n_4155),
.Y(n_4300)
);

AOI22xp5_ASAP7_75t_L g4301 ( 
.A1(n_4168),
.A2(n_254),
.B1(n_250),
.B2(n_253),
.Y(n_4301)
);

AOI21x1_ASAP7_75t_L g4302 ( 
.A1(n_4080),
.A2(n_255),
.B(n_256),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4100),
.Y(n_4303)
);

AOI22xp33_ASAP7_75t_L g4304 ( 
.A1(n_4189),
.A2(n_259),
.B1(n_256),
.B2(n_258),
.Y(n_4304)
);

INVxp67_ASAP7_75t_L g4305 ( 
.A(n_4123),
.Y(n_4305)
);

AOI22xp5_ASAP7_75t_L g4306 ( 
.A1(n_4143),
.A2(n_262),
.B1(n_259),
.B2(n_260),
.Y(n_4306)
);

OAI31xp33_ASAP7_75t_SL g4307 ( 
.A1(n_4118),
.A2(n_265),
.A3(n_266),
.B(n_263),
.Y(n_4307)
);

OAI211xp5_ASAP7_75t_L g4308 ( 
.A1(n_4142),
.A2(n_267),
.B(n_262),
.C(n_266),
.Y(n_4308)
);

OA21x2_ASAP7_75t_L g4309 ( 
.A1(n_4199),
.A2(n_267),
.B(n_268),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4217),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4109),
.B(n_269),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4115),
.B(n_269),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4165),
.B(n_270),
.Y(n_4313)
);

AND2x4_ASAP7_75t_L g4314 ( 
.A(n_4103),
.B(n_4098),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4104),
.B(n_270),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4219),
.Y(n_4316)
);

NOR3xp33_ASAP7_75t_L g4317 ( 
.A(n_4139),
.B(n_271),
.C(n_272),
.Y(n_4317)
);

AOI22xp33_ASAP7_75t_L g4318 ( 
.A1(n_4172),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_4318)
);

INVx3_ASAP7_75t_L g4319 ( 
.A(n_4077),
.Y(n_4319)
);

AO21x2_ASAP7_75t_L g4320 ( 
.A1(n_4216),
.A2(n_273),
.B(n_275),
.Y(n_4320)
);

AOI22xp33_ASAP7_75t_L g4321 ( 
.A1(n_4173),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_4321)
);

OAI21x1_ASAP7_75t_L g4322 ( 
.A1(n_4225),
.A2(n_4228),
.B(n_4226),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4220),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4231),
.Y(n_4324)
);

OA21x2_ASAP7_75t_L g4325 ( 
.A1(n_4234),
.A2(n_276),
.B(n_277),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4136),
.B(n_278),
.Y(n_4326)
);

OAI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4178),
.A2(n_278),
.B(n_279),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4232),
.Y(n_4328)
);

OAI211xp5_ASAP7_75t_SL g4329 ( 
.A1(n_4180),
.A2(n_282),
.B(n_280),
.C(n_281),
.Y(n_4329)
);

AOI22xp33_ASAP7_75t_SL g4330 ( 
.A1(n_4150),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4330)
);

INVx1_ASAP7_75t_SL g4331 ( 
.A(n_4081),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4085),
.Y(n_4332)
);

OAI221xp5_ASAP7_75t_SL g4333 ( 
.A1(n_4177),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_4333)
);

OAI211xp5_ASAP7_75t_L g4334 ( 
.A1(n_4152),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4101),
.Y(n_4335)
);

INVx1_ASAP7_75t_SL g4336 ( 
.A(n_4191),
.Y(n_4336)
);

AOI22xp33_ASAP7_75t_L g4337 ( 
.A1(n_4179),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_4337)
);

AOI33xp33_ASAP7_75t_L g4338 ( 
.A1(n_4164),
.A2(n_4182),
.A3(n_4171),
.B1(n_4161),
.B2(n_4174),
.B3(n_4151),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4193),
.B(n_288),
.Y(n_4339)
);

AOI22xp33_ASAP7_75t_SL g4340 ( 
.A1(n_4144),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_4340)
);

INVxp67_ASAP7_75t_SL g4341 ( 
.A(n_4102),
.Y(n_4341)
);

INVx3_ASAP7_75t_L g4342 ( 
.A(n_4078),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4097),
.Y(n_4343)
);

NAND3xp33_ASAP7_75t_L g4344 ( 
.A(n_4186),
.B(n_290),
.C(n_292),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4197),
.Y(n_4345)
);

BUFx3_ASAP7_75t_L g4346 ( 
.A(n_4130),
.Y(n_4346)
);

AOI22xp33_ASAP7_75t_L g4347 ( 
.A1(n_4176),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_4347)
);

OR2x2_ASAP7_75t_L g4348 ( 
.A(n_4233),
.B(n_293),
.Y(n_4348)
);

OAI222xp33_ASAP7_75t_L g4349 ( 
.A1(n_4163),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.C1(n_295),
.C2(n_298),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4195),
.B(n_4196),
.Y(n_4350)
);

AOI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_4188),
.A2(n_4106),
.B1(n_4157),
.B2(n_4108),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4200),
.B(n_294),
.Y(n_4352)
);

NOR2xp33_ASAP7_75t_L g4353 ( 
.A(n_4113),
.B(n_295),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4084),
.Y(n_4354)
);

OR2x2_ASAP7_75t_L g4355 ( 
.A(n_4082),
.B(n_4201),
.Y(n_4355)
);

OAI211xp5_ASAP7_75t_L g4356 ( 
.A1(n_4167),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_4356)
);

NAND3xp33_ASAP7_75t_L g4357 ( 
.A(n_4175),
.B(n_301),
.C(n_302),
.Y(n_4357)
);

INVx3_ASAP7_75t_L g4358 ( 
.A(n_4121),
.Y(n_4358)
);

AO21x2_ASAP7_75t_L g4359 ( 
.A1(n_4202),
.A2(n_301),
.B(n_303),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_4205),
.B(n_303),
.Y(n_4360)
);

OAI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_4110),
.A2(n_304),
.B(n_305),
.Y(n_4361)
);

OAI322xp33_ASAP7_75t_L g4362 ( 
.A1(n_4208),
.A2(n_309),
.A3(n_308),
.B1(n_306),
.B2(n_304),
.C1(n_305),
.C2(n_307),
.Y(n_4362)
);

AOI22xp5_ASAP7_75t_L g4363 ( 
.A1(n_4127),
.A2(n_4212),
.B1(n_4213),
.B2(n_4211),
.Y(n_4363)
);

AND2x4_ASAP7_75t_SL g4364 ( 
.A(n_4122),
.B(n_306),
.Y(n_4364)
);

BUFx2_ASAP7_75t_L g4365 ( 
.A(n_4214),
.Y(n_4365)
);

OAI221xp5_ASAP7_75t_L g4366 ( 
.A1(n_4229),
.A2(n_311),
.B1(n_307),
.B2(n_310),
.C(n_312),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4084),
.Y(n_4367)
);

OAI33xp33_ASAP7_75t_L g4368 ( 
.A1(n_4215),
.A2(n_312),
.A3(n_314),
.B1(n_310),
.B2(n_311),
.B3(n_313),
.Y(n_4368)
);

OAI31xp33_ASAP7_75t_L g4369 ( 
.A1(n_4218),
.A2(n_318),
.A3(n_316),
.B(n_317),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4223),
.Y(n_4370)
);

AOI221xp5_ASAP7_75t_L g4371 ( 
.A1(n_4114),
.A2(n_319),
.B1(n_316),
.B2(n_317),
.C(n_320),
.Y(n_4371)
);

OAI221xp5_ASAP7_75t_L g4372 ( 
.A1(n_4125),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.C(n_322),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4094),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4076),
.Y(n_4374)
);

INVx4_ASAP7_75t_L g4375 ( 
.A(n_4198),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4132),
.B(n_321),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4076),
.Y(n_4377)
);

AOI22xp33_ASAP7_75t_L g4378 ( 
.A1(n_4145),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_4378)
);

NAND4xp25_ASAP7_75t_L g4379 ( 
.A(n_4209),
.B(n_325),
.C(n_326),
.D(n_324),
.Y(n_4379)
);

OAI221xp5_ASAP7_75t_L g4380 ( 
.A1(n_4169),
.A2(n_326),
.B1(n_323),
.B2(n_325),
.C(n_327),
.Y(n_4380)
);

A2O1A1Ixp33_ASAP7_75t_L g4381 ( 
.A1(n_4138),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4076),
.Y(n_4382)
);

OAI31xp33_ASAP7_75t_L g4383 ( 
.A1(n_4138),
.A2(n_332),
.A3(n_329),
.B(n_330),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_4117),
.B(n_330),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_L g4385 ( 
.A1(n_4145),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_4385)
);

BUFx3_ASAP7_75t_L g4386 ( 
.A(n_4198),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_4145),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_4387)
);

OR2x2_ASAP7_75t_L g4388 ( 
.A(n_4092),
.B(n_336),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4094),
.Y(n_4389)
);

INVxp67_ASAP7_75t_L g4390 ( 
.A(n_4094),
.Y(n_4390)
);

OAI22xp5_ASAP7_75t_L g4391 ( 
.A1(n_4169),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_4391)
);

AOI22xp33_ASAP7_75t_L g4392 ( 
.A1(n_4145),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4094),
.B(n_339),
.Y(n_4393)
);

OAI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_4160),
.A2(n_340),
.B(n_341),
.Y(n_4394)
);

AOI22xp33_ASAP7_75t_SL g4395 ( 
.A1(n_4169),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_4395)
);

OAI22xp5_ASAP7_75t_L g4396 ( 
.A1(n_4169),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_4396)
);

AOI221xp5_ASAP7_75t_L g4397 ( 
.A1(n_4138),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.C(n_346),
.Y(n_4397)
);

NOR4xp25_ASAP7_75t_L g4398 ( 
.A(n_4209),
.B(n_347),
.C(n_345),
.D(n_346),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4094),
.B(n_348),
.Y(n_4399)
);

OAI31xp33_ASAP7_75t_L g4400 ( 
.A1(n_4138),
.A2(n_353),
.A3(n_350),
.B(n_352),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4094),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_4198),
.B(n_352),
.Y(n_4402)
);

AOI331xp33_ASAP7_75t_L g4403 ( 
.A1(n_4146),
.A2(n_359),
.A3(n_358),
.B1(n_355),
.B2(n_353),
.B3(n_354),
.C1(n_356),
.Y(n_4403)
);

OAI211xp5_ASAP7_75t_SL g4404 ( 
.A1(n_4096),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4076),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4094),
.Y(n_4406)
);

AOI322xp5_ASAP7_75t_L g4407 ( 
.A1(n_4160),
.A2(n_364),
.A3(n_363),
.B1(n_361),
.B2(n_359),
.C1(n_360),
.C2(n_362),
.Y(n_4407)
);

AOI22xp33_ASAP7_75t_L g4408 ( 
.A1(n_4145),
.A2(n_363),
.B1(n_360),
.B2(n_361),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_SL g4409 ( 
.A(n_4194),
.B(n_364),
.Y(n_4409)
);

AOI22xp33_ASAP7_75t_L g4410 ( 
.A1(n_4145),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_4410)
);

NOR2x1_ASAP7_75t_R g4411 ( 
.A(n_4194),
.B(n_365),
.Y(n_4411)
);

AOI221xp5_ASAP7_75t_L g4412 ( 
.A1(n_4138),
.A2(n_369),
.B1(n_366),
.B2(n_368),
.C(n_370),
.Y(n_4412)
);

AOI22xp33_ASAP7_75t_L g4413 ( 
.A1(n_4145),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_4413)
);

AND2x4_ASAP7_75t_SL g4414 ( 
.A(n_4198),
.B(n_372),
.Y(n_4414)
);

OAI221xp5_ASAP7_75t_L g4415 ( 
.A1(n_4169),
.A2(n_377),
.B1(n_373),
.B2(n_374),
.C(n_378),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4076),
.Y(n_4416)
);

OAI211xp5_ASAP7_75t_SL g4417 ( 
.A1(n_4096),
.A2(n_380),
.B(n_373),
.C(n_379),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4094),
.Y(n_4418)
);

AOI22xp33_ASAP7_75t_L g4419 ( 
.A1(n_4145),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4076),
.Y(n_4420)
);

OR2x2_ASAP7_75t_L g4421 ( 
.A(n_4092),
.B(n_383),
.Y(n_4421)
);

OR2x6_ASAP7_75t_L g4422 ( 
.A(n_4094),
.B(n_384),
.Y(n_4422)
);

OAI22xp5_ASAP7_75t_L g4423 ( 
.A1(n_4169),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_4094),
.Y(n_4424)
);

OAI211xp5_ASAP7_75t_L g4425 ( 
.A1(n_4209),
.A2(n_390),
.B(n_388),
.C(n_389),
.Y(n_4425)
);

OAI22xp5_ASAP7_75t_L g4426 ( 
.A1(n_4169),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4094),
.B(n_391),
.Y(n_4427)
);

OAI21xp5_ASAP7_75t_SL g4428 ( 
.A1(n_4169),
.A2(n_394),
.B(n_393),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4076),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_4251),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_4266),
.B(n_392),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4249),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_4386),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4252),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4269),
.B(n_392),
.Y(n_4435)
);

AND2x2_ASAP7_75t_SL g4436 ( 
.A(n_4398),
.B(n_393),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4273),
.B(n_394),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_4259),
.Y(n_4438)
);

OR2x2_ASAP7_75t_L g4439 ( 
.A(n_4246),
.B(n_395),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4254),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4365),
.B(n_396),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4335),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4235),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4288),
.Y(n_4444)
);

INVx2_ASAP7_75t_L g4445 ( 
.A(n_4277),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4346),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_4286),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4341),
.Y(n_4448)
);

AND2x4_ASAP7_75t_SL g4449 ( 
.A(n_4375),
.B(n_396),
.Y(n_4449)
);

O2A1O1Ixp33_ASAP7_75t_L g4450 ( 
.A1(n_4271),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_4450)
);

BUFx2_ASAP7_75t_L g4451 ( 
.A(n_4390),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4328),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4236),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4240),
.B(n_4373),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4237),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4239),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_4331),
.B(n_398),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4358),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4258),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4268),
.Y(n_4460)
);

HB1xp67_ASAP7_75t_L g4461 ( 
.A(n_4336),
.Y(n_4461)
);

AND2x2_ASAP7_75t_L g4462 ( 
.A(n_4389),
.B(n_399),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4279),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4285),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4287),
.Y(n_4465)
);

BUFx3_ASAP7_75t_L g4466 ( 
.A(n_4263),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4319),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4401),
.B(n_400),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_4406),
.Y(n_4469)
);

INVx2_ASAP7_75t_L g4470 ( 
.A(n_4418),
.Y(n_4470)
);

NOR2xp33_ASAP7_75t_L g4471 ( 
.A(n_4263),
.B(n_401),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4257),
.B(n_401),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4424),
.Y(n_4473)
);

AND2x2_ASAP7_75t_L g4474 ( 
.A(n_4255),
.B(n_402),
.Y(n_4474)
);

BUFx2_ASAP7_75t_L g4475 ( 
.A(n_4422),
.Y(n_4475)
);

BUFx12f_ASAP7_75t_L g4476 ( 
.A(n_4263),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4290),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4293),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4247),
.B(n_403),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4370),
.B(n_403),
.Y(n_4480)
);

AND3x1_ASAP7_75t_L g4481 ( 
.A(n_4409),
.B(n_404),
.C(n_405),
.Y(n_4481)
);

INVxp33_ASAP7_75t_L g4482 ( 
.A(n_4411),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4296),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4310),
.Y(n_4484)
);

OR2x2_ASAP7_75t_L g4485 ( 
.A(n_4342),
.B(n_405),
.Y(n_4485)
);

BUFx2_ASAP7_75t_L g4486 ( 
.A(n_4422),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4316),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4250),
.B(n_406),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4244),
.B(n_407),
.Y(n_4489)
);

INVxp67_ASAP7_75t_SL g4490 ( 
.A(n_4272),
.Y(n_4490)
);

AND2x4_ASAP7_75t_L g4491 ( 
.A(n_4314),
.B(n_407),
.Y(n_4491)
);

INVx1_ASAP7_75t_SL g4492 ( 
.A(n_4414),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_4332),
.B(n_408),
.Y(n_4493)
);

AND2x4_ASAP7_75t_SL g4494 ( 
.A(n_4384),
.B(n_408),
.Y(n_4494)
);

HB1xp67_ASAP7_75t_L g4495 ( 
.A(n_4309),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4323),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4243),
.B(n_409),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4324),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4350),
.B(n_409),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_SL g4500 ( 
.A(n_4297),
.B(n_410),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4343),
.B(n_410),
.Y(n_4501)
);

INVxp67_ASAP7_75t_L g4502 ( 
.A(n_4355),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4303),
.B(n_411),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4345),
.B(n_412),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4295),
.B(n_413),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4374),
.Y(n_4506)
);

NAND4xp25_ASAP7_75t_L g4507 ( 
.A(n_4270),
.B(n_416),
.C(n_413),
.D(n_414),
.Y(n_4507)
);

AND2x4_ASAP7_75t_SL g4508 ( 
.A(n_4393),
.B(n_4399),
.Y(n_4508)
);

BUFx2_ASAP7_75t_L g4509 ( 
.A(n_4309),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4377),
.Y(n_4510)
);

BUFx2_ASAP7_75t_L g4511 ( 
.A(n_4325),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_4322),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4382),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4338),
.B(n_4278),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4405),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4416),
.Y(n_4516)
);

AND2x2_ASAP7_75t_L g4517 ( 
.A(n_4326),
.B(n_416),
.Y(n_4517)
);

INVx2_ASAP7_75t_SL g4518 ( 
.A(n_4427),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4300),
.B(n_417),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4420),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4429),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4359),
.B(n_417),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4274),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_4351),
.B(n_419),
.Y(n_4524)
);

NAND3xp33_ASAP7_75t_L g4525 ( 
.A(n_4307),
.B(n_419),
.C(n_420),
.Y(n_4525)
);

BUFx3_ASAP7_75t_L g4526 ( 
.A(n_4364),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4325),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4388),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4421),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4315),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4280),
.Y(n_4531)
);

INVx2_ASAP7_75t_SL g4532 ( 
.A(n_4260),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4428),
.B(n_4354),
.Y(n_4533)
);

AOI22xp33_ASAP7_75t_L g4534 ( 
.A1(n_4379),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4363),
.B(n_421),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_L g4536 ( 
.A(n_4367),
.B(n_424),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4241),
.B(n_425),
.Y(n_4537)
);

AND2x2_ASAP7_75t_L g4538 ( 
.A(n_4311),
.B(n_425),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4312),
.B(n_426),
.Y(n_4539)
);

INVx5_ASAP7_75t_L g4540 ( 
.A(n_4291),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4394),
.B(n_426),
.Y(n_4541)
);

INVx2_ASAP7_75t_L g4542 ( 
.A(n_4284),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4320),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4313),
.Y(n_4544)
);

HB1xp67_ASAP7_75t_L g4545 ( 
.A(n_4299),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4339),
.B(n_4352),
.Y(n_4546)
);

AND2x4_ASAP7_75t_L g4547 ( 
.A(n_4305),
.B(n_427),
.Y(n_4547)
);

BUFx6f_ASAP7_75t_L g4548 ( 
.A(n_4348),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4267),
.B(n_428),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4353),
.B(n_428),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4376),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4289),
.B(n_429),
.Y(n_4552)
);

HB1xp67_ASAP7_75t_L g4553 ( 
.A(n_4302),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4282),
.B(n_430),
.Y(n_4554)
);

AND2x4_ASAP7_75t_L g4555 ( 
.A(n_4357),
.B(n_430),
.Y(n_4555)
);

HB1xp67_ASAP7_75t_L g4556 ( 
.A(n_4294),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4360),
.Y(n_4557)
);

BUFx6f_ASAP7_75t_L g4558 ( 
.A(n_4261),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4402),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_SL g4560 ( 
.A(n_4256),
.B(n_432),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4361),
.B(n_432),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4264),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4344),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4283),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4262),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4317),
.B(n_433),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4245),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4475),
.B(n_4486),
.Y(n_4568)
);

INVxp67_ASAP7_75t_L g4569 ( 
.A(n_4430),
.Y(n_4569)
);

AOI221xp5_ASAP7_75t_L g4570 ( 
.A1(n_4556),
.A2(n_4425),
.B1(n_4292),
.B2(n_4349),
.C(n_4396),
.Y(n_4570)
);

OAI21xp33_ASAP7_75t_L g4571 ( 
.A1(n_4436),
.A2(n_4253),
.B(n_4407),
.Y(n_4571)
);

AOI33xp33_ASAP7_75t_L g4572 ( 
.A1(n_4444),
.A2(n_4395),
.A3(n_4330),
.B1(n_4340),
.B2(n_4248),
.B3(n_4337),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4461),
.Y(n_4573)
);

BUFx2_ASAP7_75t_L g4574 ( 
.A(n_4476),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4433),
.B(n_4327),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4466),
.Y(n_4576)
);

AOI22xp33_ASAP7_75t_L g4577 ( 
.A1(n_4514),
.A2(n_4525),
.B1(n_4565),
.B2(n_4533),
.Y(n_4577)
);

AOI221xp5_ASAP7_75t_L g4578 ( 
.A1(n_4490),
.A2(n_4426),
.B1(n_4423),
.B2(n_4391),
.C(n_4412),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4495),
.Y(n_4579)
);

OR2x2_ASAP7_75t_L g4580 ( 
.A(n_4451),
.B(n_4281),
.Y(n_4580)
);

AND2x4_ASAP7_75t_L g4581 ( 
.A(n_4526),
.B(n_4265),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4540),
.Y(n_4582)
);

INVx3_ASAP7_75t_L g4583 ( 
.A(n_4431),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4509),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4511),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4505),
.Y(n_4586)
);

AOI22xp33_ASAP7_75t_L g4587 ( 
.A1(n_4500),
.A2(n_4404),
.B1(n_4417),
.B2(n_4276),
.Y(n_4587)
);

OAI22xp5_ASAP7_75t_L g4588 ( 
.A1(n_4534),
.A2(n_4347),
.B1(n_4301),
.B2(n_4381),
.Y(n_4588)
);

OAI222xp33_ASAP7_75t_L g4589 ( 
.A1(n_4553),
.A2(n_4380),
.B1(n_4415),
.B2(n_4306),
.C1(n_4366),
.C2(n_4372),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_4546),
.B(n_4518),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4540),
.B(n_4369),
.Y(n_4591)
);

HB1xp67_ASAP7_75t_L g4592 ( 
.A(n_4548),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4508),
.B(n_4383),
.Y(n_4593)
);

HB1xp67_ASAP7_75t_L g4594 ( 
.A(n_4548),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4432),
.Y(n_4595)
);

NAND3xp33_ASAP7_75t_L g4596 ( 
.A(n_4450),
.B(n_4242),
.C(n_4397),
.Y(n_4596)
);

AND2x2_ASAP7_75t_L g4597 ( 
.A(n_4443),
.B(n_4400),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4532),
.B(n_4334),
.Y(n_4598)
);

AOI22xp5_ASAP7_75t_L g4599 ( 
.A1(n_4563),
.A2(n_4368),
.B1(n_4356),
.B2(n_4308),
.Y(n_4599)
);

AND2x4_ASAP7_75t_L g4600 ( 
.A(n_4438),
.B(n_4275),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4434),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4445),
.B(n_4318),
.Y(n_4602)
);

OR2x2_ASAP7_75t_L g4603 ( 
.A(n_4530),
.B(n_4321),
.Y(n_4603)
);

AND2x4_ASAP7_75t_L g4604 ( 
.A(n_4447),
.B(n_4238),
.Y(n_4604)
);

BUFx2_ASAP7_75t_L g4605 ( 
.A(n_4558),
.Y(n_4605)
);

OR2x2_ASAP7_75t_L g4606 ( 
.A(n_4440),
.B(n_4567),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4454),
.B(n_4413),
.Y(n_4607)
);

HB1xp67_ASAP7_75t_L g4608 ( 
.A(n_4527),
.Y(n_4608)
);

OR2x2_ASAP7_75t_L g4609 ( 
.A(n_4469),
.B(n_4378),
.Y(n_4609)
);

AOI22xp33_ASAP7_75t_L g4610 ( 
.A1(n_4446),
.A2(n_4298),
.B1(n_4329),
.B2(n_4371),
.Y(n_4610)
);

AND4x1_ASAP7_75t_L g4611 ( 
.A(n_4471),
.B(n_4385),
.C(n_4387),
.D(n_4392),
.Y(n_4611)
);

OAI211xp5_ASAP7_75t_L g4612 ( 
.A1(n_4560),
.A2(n_4408),
.B(n_4419),
.C(n_4410),
.Y(n_4612)
);

OAI33xp33_ASAP7_75t_L g4613 ( 
.A1(n_4448),
.A2(n_4403),
.A3(n_4362),
.B1(n_4333),
.B2(n_4304),
.B3(n_436),
.Y(n_4613)
);

OAI31xp33_ASAP7_75t_L g4614 ( 
.A1(n_4507),
.A2(n_436),
.A3(n_434),
.B(n_435),
.Y(n_4614)
);

NOR3xp33_ASAP7_75t_L g4615 ( 
.A(n_4519),
.B(n_437),
.C(n_438),
.Y(n_4615)
);

BUFx2_ASAP7_75t_L g4616 ( 
.A(n_4558),
.Y(n_4616)
);

AOI22xp5_ASAP7_75t_L g4617 ( 
.A1(n_4562),
.A2(n_440),
.B1(n_438),
.B2(n_439),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4503),
.Y(n_4618)
);

AND2x4_ASAP7_75t_L g4619 ( 
.A(n_4458),
.B(n_439),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4492),
.B(n_440),
.Y(n_4620)
);

OAI21x1_ASAP7_75t_L g4621 ( 
.A1(n_4512),
.A2(n_441),
.B(n_442),
.Y(n_4621)
);

INVx2_ASAP7_75t_L g4622 ( 
.A(n_4467),
.Y(n_4622)
);

BUFx3_ASAP7_75t_L g4623 ( 
.A(n_4449),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4435),
.Y(n_4624)
);

AOI22xp5_ASAP7_75t_L g4625 ( 
.A1(n_4481),
.A2(n_4564),
.B1(n_4502),
.B2(n_4555),
.Y(n_4625)
);

AOI22xp33_ASAP7_75t_SL g4626 ( 
.A1(n_4531),
.A2(n_444),
.B1(n_445),
.B2(n_443),
.Y(n_4626)
);

AOI221xp5_ASAP7_75t_L g4627 ( 
.A1(n_4545),
.A2(n_4542),
.B1(n_4543),
.B2(n_4473),
.C(n_4470),
.Y(n_4627)
);

OAI31xp33_ASAP7_75t_L g4628 ( 
.A1(n_4537),
.A2(n_446),
.A3(n_442),
.B(n_443),
.Y(n_4628)
);

INVx3_ASAP7_75t_L g4629 ( 
.A(n_4491),
.Y(n_4629)
);

AND2x4_ASAP7_75t_L g4630 ( 
.A(n_4462),
.B(n_447),
.Y(n_4630)
);

OAI221xp5_ASAP7_75t_L g4631 ( 
.A1(n_4541),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.C(n_450),
.Y(n_4631)
);

AND3x2_ASAP7_75t_L g4632 ( 
.A(n_4441),
.B(n_448),
.C(n_449),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4523),
.B(n_453),
.Y(n_4633)
);

OAI21xp33_ASAP7_75t_L g4634 ( 
.A1(n_4482),
.A2(n_453),
.B(n_454),
.Y(n_4634)
);

OAI33xp33_ASAP7_75t_L g4635 ( 
.A1(n_4453),
.A2(n_457),
.A3(n_459),
.B1(n_455),
.B2(n_456),
.B3(n_458),
.Y(n_4635)
);

INVx2_ASAP7_75t_L g4636 ( 
.A(n_4468),
.Y(n_4636)
);

OA21x2_ASAP7_75t_L g4637 ( 
.A1(n_4536),
.A2(n_457),
.B(n_460),
.Y(n_4637)
);

AOI221xp5_ASAP7_75t_L g4638 ( 
.A1(n_4566),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.C(n_464),
.Y(n_4638)
);

NOR2xp33_ASAP7_75t_SL g4639 ( 
.A(n_4559),
.B(n_4437),
.Y(n_4639)
);

INVx4_ASAP7_75t_L g4640 ( 
.A(n_4494),
.Y(n_4640)
);

AOI22xp33_ASAP7_75t_L g4641 ( 
.A1(n_4557),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4497),
.Y(n_4642)
);

OAI33xp33_ASAP7_75t_L g4643 ( 
.A1(n_4455),
.A2(n_467),
.A3(n_469),
.B1(n_465),
.B2(n_466),
.B3(n_468),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4528),
.B(n_465),
.Y(n_4644)
);

AOI211xp5_ASAP7_75t_L g4645 ( 
.A1(n_4522),
.A2(n_469),
.B(n_466),
.C(n_467),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4504),
.Y(n_4646)
);

AND2x4_ASAP7_75t_L g4647 ( 
.A(n_4479),
.B(n_470),
.Y(n_4647)
);

AOI22xp5_ASAP7_75t_L g4648 ( 
.A1(n_4551),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.Y(n_4648)
);

HB1xp67_ASAP7_75t_L g4649 ( 
.A(n_4529),
.Y(n_4649)
);

INVx5_ASAP7_75t_L g4650 ( 
.A(n_4488),
.Y(n_4650)
);

OAI21xp5_ASAP7_75t_L g4651 ( 
.A1(n_4554),
.A2(n_4472),
.B(n_4561),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4544),
.B(n_4499),
.Y(n_4652)
);

CKINVDCx16_ASAP7_75t_R g4653 ( 
.A(n_4524),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4442),
.Y(n_4654)
);

INVxp67_ASAP7_75t_SL g4655 ( 
.A(n_4457),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4501),
.Y(n_4656)
);

INVxp67_ASAP7_75t_SL g4657 ( 
.A(n_4485),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4489),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4493),
.Y(n_4659)
);

AND2x4_ASAP7_75t_L g4660 ( 
.A(n_4547),
.B(n_472),
.Y(n_4660)
);

INVx1_ASAP7_75t_SL g4661 ( 
.A(n_4517),
.Y(n_4661)
);

OAI31xp33_ASAP7_75t_L g4662 ( 
.A1(n_4571),
.A2(n_4535),
.A3(n_4439),
.B(n_4552),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4608),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4582),
.B(n_4452),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4623),
.Y(n_4665)
);

AOI22xp33_ASAP7_75t_L g4666 ( 
.A1(n_4596),
.A2(n_4459),
.B1(n_4460),
.B2(n_4456),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4568),
.B(n_4474),
.Y(n_4667)
);

INVx2_ASAP7_75t_L g4668 ( 
.A(n_4574),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4649),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4573),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4579),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4653),
.B(n_4480),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4583),
.B(n_4550),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4650),
.B(n_4625),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4584),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4585),
.Y(n_4676)
);

AND2x2_ASAP7_75t_L g4677 ( 
.A(n_4640),
.B(n_4538),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4576),
.B(n_4539),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_L g4679 ( 
.A(n_4650),
.B(n_4463),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4605),
.B(n_4549),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4620),
.Y(n_4681)
);

OAI321xp33_ASAP7_75t_L g4682 ( 
.A1(n_4577),
.A2(n_4516),
.A3(n_4513),
.B1(n_4520),
.B2(n_4515),
.C(n_4510),
.Y(n_4682)
);

AND2x4_ASAP7_75t_L g4683 ( 
.A(n_4650),
.B(n_4464),
.Y(n_4683)
);

AOI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4570),
.A2(n_4589),
.B(n_4591),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4644),
.Y(n_4685)
);

AND2x4_ASAP7_75t_L g4686 ( 
.A(n_4616),
.B(n_4465),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4592),
.Y(n_4687)
);

AND3x2_ASAP7_75t_L g4688 ( 
.A(n_4645),
.B(n_4478),
.C(n_4477),
.Y(n_4688)
);

OAI33xp33_ASAP7_75t_L g4689 ( 
.A1(n_4569),
.A2(n_4496),
.A3(n_4484),
.B1(n_4498),
.B2(n_4487),
.B3(n_4483),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4594),
.B(n_4506),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4624),
.B(n_4521),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4657),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4646),
.Y(n_4693)
);

INVx2_ASAP7_75t_SL g4694 ( 
.A(n_4660),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4606),
.Y(n_4695)
);

OR2x2_ASAP7_75t_L g4696 ( 
.A(n_4580),
.B(n_473),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4581),
.B(n_473),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4656),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4632),
.B(n_474),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4586),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4618),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4659),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4590),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4629),
.B(n_474),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4595),
.Y(n_4705)
);

OR2x2_ASAP7_75t_L g4706 ( 
.A(n_4661),
.B(n_475),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4639),
.B(n_475),
.Y(n_4707)
);

BUFx2_ASAP7_75t_L g4708 ( 
.A(n_4637),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4601),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4619),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4633),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4597),
.B(n_476),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4593),
.B(n_476),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4575),
.B(n_478),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4652),
.Y(n_4715)
);

NOR2x1_ASAP7_75t_L g4716 ( 
.A(n_4598),
.B(n_479),
.Y(n_4716)
);

OR2x2_ASAP7_75t_L g4717 ( 
.A(n_4636),
.B(n_480),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4587),
.B(n_481),
.Y(n_4718)
);

AOI22xp33_ASAP7_75t_L g4719 ( 
.A1(n_4578),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4602),
.B(n_482),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4642),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4658),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4647),
.Y(n_4723)
);

BUFx3_ASAP7_75t_L g4724 ( 
.A(n_4665),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4668),
.B(n_4599),
.Y(n_4725)
);

AOI221xp5_ASAP7_75t_L g4726 ( 
.A1(n_4684),
.A2(n_4682),
.B1(n_4627),
.B2(n_4708),
.C(n_4674),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4681),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4663),
.Y(n_4728)
);

AND2x2_ASAP7_75t_SL g4729 ( 
.A(n_4680),
.B(n_4615),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4677),
.B(n_4604),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4713),
.B(n_4600),
.Y(n_4731)
);

NAND4xp25_ASAP7_75t_L g4732 ( 
.A(n_4662),
.B(n_4667),
.C(n_4666),
.D(n_4672),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4694),
.B(n_4607),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4673),
.B(n_4622),
.Y(n_4734)
);

INVx1_ASAP7_75t_SL g4735 ( 
.A(n_4706),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4669),
.Y(n_4736)
);

OR2x2_ASAP7_75t_L g4737 ( 
.A(n_4712),
.B(n_4687),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4688),
.B(n_4678),
.Y(n_4738)
);

AND2x2_ASAP7_75t_L g4739 ( 
.A(n_4710),
.B(n_4655),
.Y(n_4739)
);

AOI22xp33_ASAP7_75t_SL g4740 ( 
.A1(n_4695),
.A2(n_4588),
.B1(n_4612),
.B2(n_4631),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4692),
.Y(n_4741)
);

O2A1O1Ixp33_ASAP7_75t_L g4742 ( 
.A1(n_4707),
.A2(n_4628),
.B(n_4651),
.C(n_4634),
.Y(n_4742)
);

NOR3xp33_ASAP7_75t_L g4743 ( 
.A(n_4703),
.B(n_4638),
.C(n_4609),
.Y(n_4743)
);

INVx1_ASAP7_75t_SL g4744 ( 
.A(n_4716),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4683),
.Y(n_4745)
);

INVxp67_ASAP7_75t_SL g4746 ( 
.A(n_4699),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4704),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4720),
.B(n_4603),
.Y(n_4748)
);

NAND2x1_ASAP7_75t_SL g4749 ( 
.A(n_4714),
.B(n_4617),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4715),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4697),
.B(n_4630),
.Y(n_4751)
);

HB1xp67_ASAP7_75t_L g4752 ( 
.A(n_4686),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4723),
.Y(n_4753)
);

OR2x2_ASAP7_75t_L g4754 ( 
.A(n_4696),
.B(n_4654),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4685),
.B(n_4621),
.Y(n_4755)
);

OR2x2_ASAP7_75t_L g4756 ( 
.A(n_4664),
.B(n_4610),
.Y(n_4756)
);

OR2x2_ASAP7_75t_L g4757 ( 
.A(n_4690),
.B(n_4614),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4686),
.B(n_4572),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4717),
.Y(n_4759)
);

HB1xp67_ASAP7_75t_L g4760 ( 
.A(n_4679),
.Y(n_4760)
);

INVxp67_ASAP7_75t_L g4761 ( 
.A(n_4718),
.Y(n_4761)
);

INVx2_ASAP7_75t_L g4762 ( 
.A(n_4675),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4676),
.Y(n_4763)
);

AND2x2_ASAP7_75t_L g4764 ( 
.A(n_4722),
.B(n_4611),
.Y(n_4764)
);

OAI21xp5_ASAP7_75t_L g4765 ( 
.A1(n_4719),
.A2(n_4626),
.B(n_4648),
.Y(n_4765)
);

NOR2xp67_ASAP7_75t_L g4766 ( 
.A(n_4671),
.B(n_4641),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4691),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4670),
.B(n_4721),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4693),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4698),
.B(n_4635),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4711),
.B(n_4643),
.Y(n_4771)
);

INVxp67_ASAP7_75t_L g4772 ( 
.A(n_4752),
.Y(n_4772)
);

NOR2xp33_ASAP7_75t_L g4773 ( 
.A(n_4744),
.B(n_4689),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4730),
.B(n_4700),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4733),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4724),
.B(n_4701),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4745),
.Y(n_4777)
);

INVx4_ASAP7_75t_L g4778 ( 
.A(n_4753),
.Y(n_4778)
);

OR2x2_ASAP7_75t_L g4779 ( 
.A(n_4732),
.B(n_4702),
.Y(n_4779)
);

AND2x2_ASAP7_75t_L g4780 ( 
.A(n_4731),
.B(n_4748),
.Y(n_4780)
);

AND2x2_ASAP7_75t_L g4781 ( 
.A(n_4734),
.B(n_4705),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4739),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4760),
.Y(n_4783)
);

AND2x4_ASAP7_75t_L g4784 ( 
.A(n_4751),
.B(n_4709),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4747),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4754),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4729),
.B(n_4613),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4767),
.Y(n_4788)
);

NOR2x1p5_ASAP7_75t_SL g4789 ( 
.A(n_4757),
.B(n_483),
.Y(n_4789)
);

INVxp67_ASAP7_75t_L g4790 ( 
.A(n_4738),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4746),
.B(n_4726),
.Y(n_4791)
);

NAND2x1p5_ASAP7_75t_L g4792 ( 
.A(n_4735),
.B(n_485),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4755),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4737),
.Y(n_4794)
);

INVxp67_ASAP7_75t_SL g4795 ( 
.A(n_4749),
.Y(n_4795)
);

AND2x2_ASAP7_75t_L g4796 ( 
.A(n_4764),
.B(n_484),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4771),
.B(n_485),
.Y(n_4797)
);

AO21x2_ASAP7_75t_L g4798 ( 
.A1(n_4725),
.A2(n_488),
.B(n_487),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4741),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4759),
.B(n_486),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4727),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4762),
.Y(n_4802)
);

AND2x4_ASAP7_75t_L g4803 ( 
.A(n_4750),
.B(n_488),
.Y(n_4803)
);

BUFx3_ASAP7_75t_L g4804 ( 
.A(n_4728),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4768),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4766),
.B(n_489),
.Y(n_4806)
);

NOR2xp33_ASAP7_75t_L g4807 ( 
.A(n_4758),
.B(n_489),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4736),
.Y(n_4808)
);

INVx3_ASAP7_75t_L g4809 ( 
.A(n_4763),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4761),
.B(n_490),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4765),
.B(n_490),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4769),
.Y(n_4812)
);

AOI22xp5_ASAP7_75t_L g4813 ( 
.A1(n_4743),
.A2(n_4740),
.B1(n_4770),
.B2(n_4756),
.Y(n_4813)
);

INVx2_ASAP7_75t_L g4814 ( 
.A(n_4742),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4730),
.B(n_492),
.Y(n_4815)
);

OAI31xp33_ASAP7_75t_SL g4816 ( 
.A1(n_4726),
.A2(n_494),
.A3(n_492),
.B(n_493),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4730),
.B(n_493),
.Y(n_4817)
);

INVx1_ASAP7_75t_SL g4818 ( 
.A(n_4744),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4752),
.B(n_495),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_L g4820 ( 
.A(n_4752),
.B(n_496),
.Y(n_4820)
);

INVx3_ASAP7_75t_L g4821 ( 
.A(n_4778),
.Y(n_4821)
);

OR2x2_ASAP7_75t_L g4822 ( 
.A(n_4792),
.B(n_496),
.Y(n_4822)
);

OAI211xp5_ASAP7_75t_L g4823 ( 
.A1(n_4813),
.A2(n_501),
.B(n_497),
.C(n_499),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4780),
.Y(n_4824)
);

NOR2xp33_ASAP7_75t_SL g4825 ( 
.A(n_4818),
.B(n_497),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4795),
.B(n_499),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4774),
.Y(n_4827)
);

AND2x2_ASAP7_75t_L g4828 ( 
.A(n_4815),
.B(n_501),
.Y(n_4828)
);

AND2x2_ASAP7_75t_L g4829 ( 
.A(n_4817),
.B(n_502),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4772),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4820),
.Y(n_4831)
);

NAND3xp33_ASAP7_75t_SL g4832 ( 
.A(n_4773),
.B(n_4791),
.C(n_4787),
.Y(n_4832)
);

INVx1_ASAP7_75t_SL g4833 ( 
.A(n_4806),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4777),
.B(n_502),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4793),
.B(n_503),
.Y(n_4835)
);

INVx2_ASAP7_75t_L g4836 ( 
.A(n_4784),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4816),
.B(n_503),
.Y(n_4837)
);

OAI21xp33_ASAP7_75t_L g4838 ( 
.A1(n_4790),
.A2(n_504),
.B(n_505),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4819),
.Y(n_4839)
);

OR2x2_ASAP7_75t_L g4840 ( 
.A(n_4797),
.B(n_505),
.Y(n_4840)
);

INVx2_ASAP7_75t_L g4841 ( 
.A(n_4781),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4796),
.B(n_507),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4789),
.B(n_507),
.Y(n_4843)
);

INVx2_ASAP7_75t_SL g4844 ( 
.A(n_4803),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4776),
.Y(n_4845)
);

AOI322xp5_ASAP7_75t_L g4846 ( 
.A1(n_4814),
.A2(n_514),
.A3(n_513),
.B1(n_511),
.B2(n_508),
.C1(n_509),
.C2(n_512),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4782),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4811),
.B(n_512),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4800),
.Y(n_4849)
);

OAI21xp5_ASAP7_75t_L g4850 ( 
.A1(n_4807),
.A2(n_514),
.B(n_515),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4804),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4783),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4785),
.B(n_516),
.Y(n_4853)
);

INVxp67_ASAP7_75t_SL g4854 ( 
.A(n_4786),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4810),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4794),
.B(n_516),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4788),
.Y(n_4857)
);

INVxp67_ASAP7_75t_L g4858 ( 
.A(n_4798),
.Y(n_4858)
);

NOR2xp33_ASAP7_75t_L g4859 ( 
.A(n_4779),
.B(n_517),
.Y(n_4859)
);

AND2x2_ASAP7_75t_L g4860 ( 
.A(n_4775),
.B(n_517),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4802),
.B(n_518),
.Y(n_4861)
);

NOR2xp33_ASAP7_75t_L g4862 ( 
.A(n_4809),
.B(n_519),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_4808),
.B(n_519),
.Y(n_4863)
);

AND2x4_ASAP7_75t_L g4864 ( 
.A(n_4801),
.B(n_520),
.Y(n_4864)
);

NAND2xp33_ASAP7_75t_L g4865 ( 
.A(n_4805),
.B(n_520),
.Y(n_4865)
);

HB1xp67_ASAP7_75t_L g4866 ( 
.A(n_4799),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4812),
.Y(n_4867)
);

OR2x2_ASAP7_75t_L g4868 ( 
.A(n_4792),
.B(n_521),
.Y(n_4868)
);

OR2x2_ASAP7_75t_L g4869 ( 
.A(n_4792),
.B(n_521),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_L g4870 ( 
.A(n_4780),
.B(n_522),
.Y(n_4870)
);

OR2x6_ASAP7_75t_L g4871 ( 
.A(n_4772),
.B(n_523),
.Y(n_4871)
);

INVx2_ASAP7_75t_SL g4872 ( 
.A(n_4774),
.Y(n_4872)
);

AND2x4_ASAP7_75t_L g4873 ( 
.A(n_4780),
.B(n_523),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4792),
.Y(n_4874)
);

INVx1_ASAP7_75t_SL g4875 ( 
.A(n_4780),
.Y(n_4875)
);

INVx2_ASAP7_75t_L g4876 ( 
.A(n_4780),
.Y(n_4876)
);

INVxp67_ASAP7_75t_SL g4877 ( 
.A(n_4792),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4877),
.Y(n_4878)
);

AOI211x1_ASAP7_75t_L g4879 ( 
.A1(n_4823),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_4879)
);

AOI22xp5_ASAP7_75t_L g4880 ( 
.A1(n_4832),
.A2(n_527),
.B1(n_524),
.B2(n_526),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4875),
.B(n_527),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4824),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4876),
.Y(n_4883)
);

AND2x2_ASAP7_75t_L g4884 ( 
.A(n_4872),
.B(n_528),
.Y(n_4884)
);

AND2x2_ASAP7_75t_L g4885 ( 
.A(n_4836),
.B(n_529),
.Y(n_4885)
);

OAI22xp33_ASAP7_75t_L g4886 ( 
.A1(n_4825),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_4886)
);

INVxp67_ASAP7_75t_L g4887 ( 
.A(n_4822),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4868),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4833),
.B(n_530),
.Y(n_4889)
);

OAI22xp33_ASAP7_75t_L g4890 ( 
.A1(n_4874),
.A2(n_534),
.B1(n_531),
.B2(n_533),
.Y(n_4890)
);

AOI222xp33_ASAP7_75t_L g4891 ( 
.A1(n_4858),
.A2(n_537),
.B1(n_539),
.B2(n_533),
.C1(n_535),
.C2(n_538),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4869),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4842),
.Y(n_4893)
);

INVx2_ASAP7_75t_L g4894 ( 
.A(n_4871),
.Y(n_4894)
);

INVxp67_ASAP7_75t_SL g4895 ( 
.A(n_4821),
.Y(n_4895)
);

OR2x2_ASAP7_75t_L g4896 ( 
.A(n_4827),
.B(n_537),
.Y(n_4896)
);

INVxp67_ASAP7_75t_L g4897 ( 
.A(n_4843),
.Y(n_4897)
);

INVxp67_ASAP7_75t_SL g4898 ( 
.A(n_4854),
.Y(n_4898)
);

AND2x2_ASAP7_75t_L g4899 ( 
.A(n_4841),
.B(n_538),
.Y(n_4899)
);

NAND3xp33_ASAP7_75t_L g4900 ( 
.A(n_4865),
.B(n_539),
.C(n_540),
.Y(n_4900)
);

AOI22xp5_ASAP7_75t_L g4901 ( 
.A1(n_4830),
.A2(n_544),
.B1(n_541),
.B2(n_542),
.Y(n_4901)
);

AOI211xp5_ASAP7_75t_L g4902 ( 
.A1(n_4859),
.A2(n_545),
.B(n_541),
.C(n_542),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4870),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4828),
.Y(n_4904)
);

OAI21xp5_ASAP7_75t_L g4905 ( 
.A1(n_4826),
.A2(n_545),
.B(n_548),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4844),
.B(n_548),
.Y(n_4906)
);

NAND3xp33_ASAP7_75t_L g4907 ( 
.A(n_4866),
.B(n_550),
.C(n_551),
.Y(n_4907)
);

OAI22xp33_ASAP7_75t_L g4908 ( 
.A1(n_4837),
.A2(n_554),
.B1(n_550),
.B2(n_552),
.Y(n_4908)
);

OAI21xp5_ASAP7_75t_SL g4909 ( 
.A1(n_4847),
.A2(n_554),
.B(n_555),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4829),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4848),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4873),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4871),
.Y(n_4913)
);

NAND2x1p5_ASAP7_75t_L g4914 ( 
.A(n_4851),
.B(n_556),
.Y(n_4914)
);

NAND2xp5_ASAP7_75t_L g4915 ( 
.A(n_4846),
.B(n_556),
.Y(n_4915)
);

OAI21xp33_ASAP7_75t_L g4916 ( 
.A1(n_4849),
.A2(n_568),
.B(n_557),
.Y(n_4916)
);

OAI322xp33_ASAP7_75t_L g4917 ( 
.A1(n_4852),
.A2(n_563),
.A3(n_562),
.B1(n_559),
.B2(n_557),
.C1(n_558),
.C2(n_561),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4856),
.Y(n_4918)
);

OAI21xp33_ASAP7_75t_L g4919 ( 
.A1(n_4845),
.A2(n_570),
.B(n_558),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4840),
.B(n_559),
.Y(n_4920)
);

OR2x2_ASAP7_75t_L g4921 ( 
.A(n_4835),
.B(n_561),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4853),
.Y(n_4922)
);

OAI222xp33_ASAP7_75t_L g4923 ( 
.A1(n_4857),
.A2(n_564),
.B1(n_569),
.B2(n_562),
.C1(n_563),
.C2(n_567),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4861),
.B(n_564),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4862),
.B(n_567),
.Y(n_4925)
);

AND2x2_ASAP7_75t_L g4926 ( 
.A(n_4855),
.B(n_571),
.Y(n_4926)
);

INVx2_ASAP7_75t_L g4927 ( 
.A(n_4864),
.Y(n_4927)
);

AOI22xp5_ASAP7_75t_L g4928 ( 
.A1(n_4838),
.A2(n_574),
.B1(n_571),
.B2(n_572),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4860),
.B(n_572),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4834),
.Y(n_4930)
);

OR2x2_ASAP7_75t_L g4931 ( 
.A(n_4863),
.B(n_574),
.Y(n_4931)
);

OAI22xp33_ASAP7_75t_L g4932 ( 
.A1(n_4831),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4839),
.B(n_576),
.Y(n_4933)
);

AOI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4867),
.A2(n_580),
.B1(n_577),
.B2(n_579),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4850),
.Y(n_4935)
);

AND2x2_ASAP7_75t_SL g4936 ( 
.A(n_4874),
.B(n_580),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4875),
.B(n_581),
.Y(n_4937)
);

AOI32xp33_ASAP7_75t_L g4938 ( 
.A1(n_4875),
.A2(n_583),
.A3(n_581),
.B1(n_582),
.B2(n_584),
.Y(n_4938)
);

INVx2_ASAP7_75t_L g4939 ( 
.A(n_4824),
.Y(n_4939)
);

AOI211xp5_ASAP7_75t_L g4940 ( 
.A1(n_4832),
.A2(n_584),
.B(n_582),
.C(n_583),
.Y(n_4940)
);

OAI222xp33_ASAP7_75t_L g4941 ( 
.A1(n_4875),
.A2(n_588),
.B1(n_591),
.B2(n_586),
.C1(n_587),
.C2(n_590),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4877),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4877),
.Y(n_4943)
);

AOI321xp33_ASAP7_75t_L g4944 ( 
.A1(n_4854),
.A2(n_590),
.A3(n_592),
.B1(n_586),
.B2(n_588),
.C(n_591),
.Y(n_4944)
);

AOI211xp5_ASAP7_75t_SL g4945 ( 
.A1(n_4877),
.A2(n_596),
.B(n_592),
.C(n_595),
.Y(n_4945)
);

OR2x2_ASAP7_75t_L g4946 ( 
.A(n_4875),
.B(n_596),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4824),
.Y(n_4947)
);

AOI321xp33_ASAP7_75t_L g4948 ( 
.A1(n_4854),
.A2(n_599),
.A3(n_601),
.B1(n_597),
.B2(n_598),
.C(n_600),
.Y(n_4948)
);

O2A1O1Ixp33_ASAP7_75t_L g4949 ( 
.A1(n_4832),
.A2(n_610),
.B(n_618),
.C(n_599),
.Y(n_4949)
);

AOI22xp5_ASAP7_75t_L g4950 ( 
.A1(n_4832),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_4950)
);

INVxp67_ASAP7_75t_L g4951 ( 
.A(n_4825),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4877),
.Y(n_4952)
);

OAI21xp5_ASAP7_75t_L g4953 ( 
.A1(n_4832),
.A2(n_602),
.B(n_603),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4877),
.Y(n_4954)
);

AOI22xp5_ASAP7_75t_L g4955 ( 
.A1(n_4832),
.A2(n_608),
.B1(n_605),
.B2(n_606),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_L g4956 ( 
.A(n_4875),
.B(n_605),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4875),
.B(n_606),
.Y(n_4957)
);

INVxp33_ASAP7_75t_L g4958 ( 
.A(n_4824),
.Y(n_4958)
);

OAI22xp5_ASAP7_75t_L g4959 ( 
.A1(n_4875),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_4959)
);

AOI22xp33_ASAP7_75t_L g4960 ( 
.A1(n_4832),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.Y(n_4960)
);

O2A1O1Ixp33_ASAP7_75t_SL g4961 ( 
.A1(n_4858),
.A2(n_616),
.B(n_614),
.C(n_615),
.Y(n_4961)
);

OAI22xp5_ASAP7_75t_L g4962 ( 
.A1(n_4875),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_4962)
);

OAI221xp5_ASAP7_75t_L g4963 ( 
.A1(n_4875),
.A2(n_619),
.B1(n_617),
.B2(n_618),
.C(n_620),
.Y(n_4963)
);

AOI22x1_ASAP7_75t_L g4964 ( 
.A1(n_4877),
.A2(n_622),
.B1(n_619),
.B2(n_621),
.Y(n_4964)
);

NAND2xp5_ASAP7_75t_L g4965 ( 
.A(n_4875),
.B(n_621),
.Y(n_4965)
);

OAI21xp33_ASAP7_75t_L g4966 ( 
.A1(n_4875),
.A2(n_631),
.B(n_623),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4877),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4906),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4895),
.Y(n_4969)
);

XNOR2xp5_ASAP7_75t_L g4970 ( 
.A(n_4958),
.B(n_623),
.Y(n_4970)
);

NOR2xp33_ASAP7_75t_L g4971 ( 
.A(n_4951),
.B(n_4913),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4914),
.Y(n_4972)
);

XNOR2xp5_ASAP7_75t_L g4973 ( 
.A(n_4879),
.B(n_624),
.Y(n_4973)
);

XNOR2xp5_ASAP7_75t_L g4974 ( 
.A(n_4964),
.B(n_625),
.Y(n_4974)
);

AND2x4_ASAP7_75t_L g4975 ( 
.A(n_4898),
.B(n_625),
.Y(n_4975)
);

OR2x2_ASAP7_75t_L g4976 ( 
.A(n_4946),
.B(n_626),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4939),
.B(n_626),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4945),
.B(n_627),
.Y(n_4978)
);

XOR2x2_ASAP7_75t_L g4979 ( 
.A(n_4900),
.B(n_627),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4884),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4961),
.Y(n_4981)
);

XOR2x2_ASAP7_75t_L g4982 ( 
.A(n_4940),
.B(n_628),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4936),
.B(n_628),
.Y(n_4983)
);

OAI222xp33_ASAP7_75t_L g4984 ( 
.A1(n_4878),
.A2(n_631),
.B1(n_633),
.B2(n_629),
.C1(n_630),
.C2(n_632),
.Y(n_4984)
);

AOI22xp33_ASAP7_75t_L g4985 ( 
.A1(n_4947),
.A2(n_632),
.B1(n_629),
.B2(n_630),
.Y(n_4985)
);

AOI22xp33_ASAP7_75t_SL g4986 ( 
.A1(n_4882),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_4986)
);

INVx2_ASAP7_75t_L g4987 ( 
.A(n_4920),
.Y(n_4987)
);

OAI21xp33_ASAP7_75t_L g4988 ( 
.A1(n_4942),
.A2(n_634),
.B(n_635),
.Y(n_4988)
);

AOI21xp5_ASAP7_75t_L g4989 ( 
.A1(n_4949),
.A2(n_637),
.B(n_638),
.Y(n_4989)
);

BUFx2_ASAP7_75t_L g4990 ( 
.A(n_4894),
.Y(n_4990)
);

INVx4_ASAP7_75t_L g4991 ( 
.A(n_4885),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4881),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4937),
.Y(n_4993)
);

XNOR2x2_ASAP7_75t_L g4994 ( 
.A(n_4953),
.B(n_637),
.Y(n_4994)
);

AOI21xp5_ASAP7_75t_SL g4995 ( 
.A1(n_4956),
.A2(n_4965),
.B(n_4957),
.Y(n_4995)
);

AND2x2_ASAP7_75t_L g4996 ( 
.A(n_4927),
.B(n_638),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4912),
.B(n_639),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4938),
.B(n_639),
.Y(n_4998)
);

NAND2xp5_ASAP7_75t_L g4999 ( 
.A(n_4891),
.B(n_640),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4899),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_4896),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_L g5002 ( 
.A(n_4893),
.B(n_640),
.Y(n_5002)
);

NAND3xp33_ASAP7_75t_L g5003 ( 
.A(n_4960),
.B(n_641),
.C(n_642),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_4926),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_L g5005 ( 
.A(n_4904),
.B(n_641),
.Y(n_5005)
);

NAND2xp5_ASAP7_75t_SL g5006 ( 
.A(n_4944),
.B(n_642),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4889),
.Y(n_5007)
);

NAND3xp33_ASAP7_75t_SL g5008 ( 
.A(n_4880),
.B(n_643),
.C(n_644),
.Y(n_5008)
);

INVx1_ASAP7_75t_SL g5009 ( 
.A(n_4929),
.Y(n_5009)
);

OAI321xp33_ASAP7_75t_L g5010 ( 
.A1(n_4943),
.A2(n_645),
.A3(n_647),
.B1(n_643),
.B2(n_644),
.C(n_646),
.Y(n_5010)
);

XNOR2xp5_ASAP7_75t_L g5011 ( 
.A(n_4910),
.B(n_645),
.Y(n_5011)
);

NAND4xp25_ASAP7_75t_L g5012 ( 
.A(n_4952),
.B(n_648),
.C(n_646),
.D(n_647),
.Y(n_5012)
);

AND2x2_ASAP7_75t_L g5013 ( 
.A(n_4883),
.B(n_648),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_SL g5014 ( 
.A(n_4948),
.B(n_649),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4911),
.Y(n_5015)
);

AOI221x1_ASAP7_75t_SL g5016 ( 
.A1(n_4954),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.C(n_652),
.Y(n_5016)
);

AOI221xp5_ASAP7_75t_L g5017 ( 
.A1(n_4967),
.A2(n_653),
.B1(n_650),
.B2(n_652),
.C(n_654),
.Y(n_5017)
);

NAND2xp33_ASAP7_75t_SL g5018 ( 
.A(n_4888),
.B(n_653),
.Y(n_5018)
);

INVxp67_ASAP7_75t_L g5019 ( 
.A(n_4915),
.Y(n_5019)
);

BUFx2_ASAP7_75t_SL g5020 ( 
.A(n_4892),
.Y(n_5020)
);

NOR2x1_ASAP7_75t_L g5021 ( 
.A(n_4941),
.B(n_654),
.Y(n_5021)
);

INVxp67_ASAP7_75t_L g5022 ( 
.A(n_4924),
.Y(n_5022)
);

OR2x2_ASAP7_75t_L g5023 ( 
.A(n_4918),
.B(n_4922),
.Y(n_5023)
);

NOR2xp33_ASAP7_75t_L g5024 ( 
.A(n_4897),
.B(n_4966),
.Y(n_5024)
);

OR2x2_ASAP7_75t_L g5025 ( 
.A(n_4931),
.B(n_655),
.Y(n_5025)
);

OR2x2_ASAP7_75t_L g5026 ( 
.A(n_4921),
.B(n_655),
.Y(n_5026)
);

A2O1A1Ixp33_ASAP7_75t_L g5027 ( 
.A1(n_4950),
.A2(n_658),
.B(n_656),
.C(n_657),
.Y(n_5027)
);

BUFx3_ASAP7_75t_L g5028 ( 
.A(n_4903),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4925),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_4887),
.B(n_657),
.Y(n_5030)
);

NOR3xp33_ASAP7_75t_L g5031 ( 
.A(n_4908),
.B(n_658),
.C(n_659),
.Y(n_5031)
);

OAI21xp33_ASAP7_75t_L g5032 ( 
.A1(n_4935),
.A2(n_4955),
.B(n_4930),
.Y(n_5032)
);

XNOR2xp5_ASAP7_75t_L g5033 ( 
.A(n_4928),
.B(n_659),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_L g5034 ( 
.A(n_4886),
.B(n_660),
.Y(n_5034)
);

NOR3xp33_ASAP7_75t_L g5035 ( 
.A(n_4933),
.B(n_660),
.C(n_661),
.Y(n_5035)
);

INVx1_ASAP7_75t_SL g5036 ( 
.A(n_4959),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_4890),
.B(n_661),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_4907),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4962),
.Y(n_5039)
);

AND2x2_ASAP7_75t_L g5040 ( 
.A(n_4905),
.B(n_662),
.Y(n_5040)
);

XNOR2xp5_ASAP7_75t_L g5041 ( 
.A(n_4902),
.B(n_662),
.Y(n_5041)
);

INVxp67_ASAP7_75t_L g5042 ( 
.A(n_4963),
.Y(n_5042)
);

INVx1_ASAP7_75t_SL g5043 ( 
.A(n_4901),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4909),
.B(n_663),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4916),
.B(n_664),
.Y(n_5045)
);

OR2x2_ASAP7_75t_L g5046 ( 
.A(n_4919),
.B(n_665),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4934),
.Y(n_5047)
);

NOR4xp75_ASAP7_75t_L g5048 ( 
.A(n_4917),
.B(n_668),
.C(n_665),
.D(n_667),
.Y(n_5048)
);

OR2x2_ASAP7_75t_L g5049 ( 
.A(n_4932),
.B(n_668),
.Y(n_5049)
);

NOR2xp33_ASAP7_75t_L g5050 ( 
.A(n_4923),
.B(n_669),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4906),
.Y(n_5051)
);

BUFx3_ASAP7_75t_L g5052 ( 
.A(n_4914),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4895),
.B(n_670),
.Y(n_5053)
);

AND2x2_ASAP7_75t_L g5054 ( 
.A(n_4895),
.B(n_670),
.Y(n_5054)
);

A2O1A1Ixp33_ASAP7_75t_L g5055 ( 
.A1(n_5016),
.A2(n_673),
.B(n_671),
.C(n_672),
.Y(n_5055)
);

INVxp67_ASAP7_75t_SL g5056 ( 
.A(n_5021),
.Y(n_5056)
);

NOR2xp33_ASAP7_75t_L g5057 ( 
.A(n_4991),
.B(n_671),
.Y(n_5057)
);

NOR2xp33_ASAP7_75t_L g5058 ( 
.A(n_4991),
.B(n_672),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_SL g5059 ( 
.A(n_4981),
.B(n_674),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_5054),
.Y(n_5060)
);

NAND3x1_ASAP7_75t_L g5061 ( 
.A(n_5048),
.B(n_674),
.C(n_675),
.Y(n_5061)
);

AOI22xp5_ASAP7_75t_L g5062 ( 
.A1(n_4971),
.A2(n_679),
.B1(n_677),
.B2(n_678),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_4970),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_4990),
.B(n_679),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4996),
.B(n_680),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_5011),
.Y(n_5066)
);

OAI322xp33_ASAP7_75t_L g5067 ( 
.A1(n_5019),
.A2(n_685),
.A3(n_684),
.B1(n_682),
.B2(n_680),
.C1(n_681),
.C2(n_683),
.Y(n_5067)
);

NAND3xp33_ASAP7_75t_L g5068 ( 
.A(n_5018),
.B(n_682),
.C(n_685),
.Y(n_5068)
);

OAI22xp5_ASAP7_75t_L g5069 ( 
.A1(n_4969),
.A2(n_688),
.B1(n_686),
.B2(n_687),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_4974),
.Y(n_5070)
);

AND2x2_ASAP7_75t_L g5071 ( 
.A(n_4972),
.B(n_687),
.Y(n_5071)
);

O2A1O1Ixp33_ASAP7_75t_SL g5072 ( 
.A1(n_5006),
.A2(n_697),
.B(n_705),
.C(n_689),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4975),
.Y(n_5073)
);

AOI21xp5_ASAP7_75t_L g5074 ( 
.A1(n_4983),
.A2(n_5014),
.B(n_4995),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4975),
.Y(n_5075)
);

INVx1_ASAP7_75t_SL g5076 ( 
.A(n_5020),
.Y(n_5076)
);

AOI22xp5_ASAP7_75t_L g5077 ( 
.A1(n_5036),
.A2(n_691),
.B1(n_689),
.B2(n_690),
.Y(n_5077)
);

NOR2x1_ASAP7_75t_L g5078 ( 
.A(n_5012),
.B(n_690),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4978),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_5013),
.Y(n_5080)
);

BUFx2_ASAP7_75t_L g5081 ( 
.A(n_5052),
.Y(n_5081)
);

INVxp67_ASAP7_75t_L g5082 ( 
.A(n_5050),
.Y(n_5082)
);

XNOR2x2_ASAP7_75t_L g5083 ( 
.A(n_4994),
.B(n_691),
.Y(n_5083)
);

OAI321xp33_ASAP7_75t_L g5084 ( 
.A1(n_5042),
.A2(n_694),
.A3(n_696),
.B1(n_692),
.B2(n_693),
.C(n_695),
.Y(n_5084)
);

AOI222xp33_ASAP7_75t_L g5085 ( 
.A1(n_5032),
.A2(n_698),
.B1(n_700),
.B2(n_694),
.C1(n_696),
.C2(n_699),
.Y(n_5085)
);

INVx2_ASAP7_75t_L g5086 ( 
.A(n_4976),
.Y(n_5086)
);

O2A1O1Ixp33_ASAP7_75t_L g5087 ( 
.A1(n_4984),
.A2(n_701),
.B(n_699),
.C(n_700),
.Y(n_5087)
);

AOI21xp5_ASAP7_75t_L g5088 ( 
.A1(n_4989),
.A2(n_701),
.B(n_702),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4977),
.Y(n_5089)
);

NOR3xp33_ASAP7_75t_L g5090 ( 
.A(n_5024),
.B(n_704),
.C(n_703),
.Y(n_5090)
);

HB1xp67_ASAP7_75t_L g5091 ( 
.A(n_4973),
.Y(n_5091)
);

OR2x2_ASAP7_75t_L g5092 ( 
.A(n_5053),
.B(n_5023),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_5030),
.Y(n_5093)
);

OR2x2_ASAP7_75t_L g5094 ( 
.A(n_4997),
.B(n_702),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_5041),
.Y(n_5095)
);

AOI22xp5_ASAP7_75t_L g5096 ( 
.A1(n_5043),
.A2(n_705),
.B1(n_703),
.B2(n_704),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4968),
.Y(n_5097)
);

NAND2xp5_ASAP7_75t_L g5098 ( 
.A(n_4986),
.B(n_5051),
.Y(n_5098)
);

OR2x2_ASAP7_75t_L g5099 ( 
.A(n_4999),
.B(n_706),
.Y(n_5099)
);

NAND2xp33_ASAP7_75t_L g5100 ( 
.A(n_5035),
.B(n_706),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_5002),
.Y(n_5101)
);

INVx2_ASAP7_75t_L g5102 ( 
.A(n_5025),
.Y(n_5102)
);

AO22x1_ASAP7_75t_L g5103 ( 
.A1(n_5031),
.A2(n_709),
.B1(n_707),
.B2(n_708),
.Y(n_5103)
);

AND2x2_ASAP7_75t_L g5104 ( 
.A(n_4980),
.B(n_707),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5005),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_5033),
.Y(n_5106)
);

OA22x2_ASAP7_75t_L g5107 ( 
.A1(n_5004),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5049),
.Y(n_5108)
);

OAI222xp33_ASAP7_75t_L g5109 ( 
.A1(n_5015),
.A2(n_712),
.B1(n_714),
.B2(n_710),
.C1(n_711),
.C2(n_713),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_5045),
.B(n_713),
.Y(n_5110)
);

AND2x2_ASAP7_75t_L g5111 ( 
.A(n_4987),
.B(n_716),
.Y(n_5111)
);

NAND2xp5_ASAP7_75t_L g5112 ( 
.A(n_5000),
.B(n_717),
.Y(n_5112)
);

AOI322xp5_ASAP7_75t_L g5113 ( 
.A1(n_5039),
.A2(n_722),
.A3(n_721),
.B1(n_719),
.B2(n_717),
.C1(n_718),
.C2(n_720),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5040),
.B(n_718),
.Y(n_5114)
);

OAI21xp5_ASAP7_75t_SL g5115 ( 
.A1(n_5008),
.A2(n_721),
.B(n_723),
.Y(n_5115)
);

OAI221xp5_ASAP7_75t_SL g5116 ( 
.A1(n_5038),
.A2(n_5047),
.B1(n_5009),
.B2(n_5022),
.C(n_4993),
.Y(n_5116)
);

AND2x2_ASAP7_75t_L g5117 ( 
.A(n_5001),
.B(n_724),
.Y(n_5117)
);

OAI22xp5_ASAP7_75t_L g5118 ( 
.A1(n_5003),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.Y(n_5118)
);

AND2x2_ASAP7_75t_L g5119 ( 
.A(n_5028),
.B(n_726),
.Y(n_5119)
);

CKINVDCx16_ASAP7_75t_R g5120 ( 
.A(n_5026),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_4988),
.B(n_728),
.Y(n_5121)
);

OR2x2_ASAP7_75t_L g5122 ( 
.A(n_4998),
.B(n_729),
.Y(n_5122)
);

HB1xp67_ASAP7_75t_L g5123 ( 
.A(n_4982),
.Y(n_5123)
);

AOI22xp33_ASAP7_75t_L g5124 ( 
.A1(n_4992),
.A2(n_731),
.B1(n_729),
.B2(n_730),
.Y(n_5124)
);

AOI222xp33_ASAP7_75t_L g5125 ( 
.A1(n_5007),
.A2(n_732),
.B1(n_734),
.B2(n_730),
.C1(n_731),
.C2(n_733),
.Y(n_5125)
);

AOI221xp5_ASAP7_75t_SL g5126 ( 
.A1(n_5027),
.A2(n_737),
.B1(n_732),
.B2(n_736),
.C(n_738),
.Y(n_5126)
);

AOI221xp5_ASAP7_75t_L g5127 ( 
.A1(n_5010),
.A2(n_739),
.B1(n_736),
.B2(n_738),
.C(n_740),
.Y(n_5127)
);

AND2x2_ASAP7_75t_L g5128 ( 
.A(n_5029),
.B(n_739),
.Y(n_5128)
);

OR2x2_ASAP7_75t_L g5129 ( 
.A(n_5037),
.B(n_740),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_5046),
.Y(n_5130)
);

INVx2_ASAP7_75t_SL g5131 ( 
.A(n_4979),
.Y(n_5131)
);

INVxp67_ASAP7_75t_L g5132 ( 
.A(n_5044),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_5034),
.Y(n_5133)
);

INVx3_ASAP7_75t_L g5134 ( 
.A(n_4985),
.Y(n_5134)
);

OAI21xp5_ASAP7_75t_L g5135 ( 
.A1(n_5017),
.A2(n_746),
.B(n_745),
.Y(n_5135)
);

OA211x2_ASAP7_75t_L g5136 ( 
.A1(n_4988),
.A2(n_748),
.B(n_742),
.C(n_745),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_5054),
.Y(n_5137)
);

AND2x2_ASAP7_75t_L g5138 ( 
.A(n_4990),
.B(n_742),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_5054),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_5054),
.Y(n_5140)
);

XNOR2xp5_ASAP7_75t_L g5141 ( 
.A(n_5048),
.B(n_748),
.Y(n_5141)
);

AOI211x1_ASAP7_75t_SL g5142 ( 
.A1(n_5074),
.A2(n_751),
.B(n_749),
.C(n_750),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_5138),
.Y(n_5143)
);

INVx2_ASAP7_75t_L g5144 ( 
.A(n_5107),
.Y(n_5144)
);

OAI31xp33_ASAP7_75t_L g5145 ( 
.A1(n_5076),
.A2(n_758),
.A3(n_766),
.B(n_750),
.Y(n_5145)
);

OAI321xp33_ASAP7_75t_L g5146 ( 
.A1(n_5116),
.A2(n_753),
.A3(n_755),
.B1(n_751),
.B2(n_752),
.C(n_754),
.Y(n_5146)
);

NAND3xp33_ASAP7_75t_L g5147 ( 
.A(n_5127),
.B(n_752),
.C(n_756),
.Y(n_5147)
);

AOI322xp5_ASAP7_75t_L g5148 ( 
.A1(n_5056),
.A2(n_762),
.A3(n_761),
.B1(n_759),
.B2(n_756),
.C1(n_757),
.C2(n_760),
.Y(n_5148)
);

OAI21xp33_ASAP7_75t_L g5149 ( 
.A1(n_5098),
.A2(n_757),
.B(n_760),
.Y(n_5149)
);

INVx1_ASAP7_75t_SL g5150 ( 
.A(n_5083),
.Y(n_5150)
);

AOI221xp5_ASAP7_75t_L g5151 ( 
.A1(n_5072),
.A2(n_764),
.B1(n_761),
.B2(n_763),
.C(n_765),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5073),
.Y(n_5152)
);

OAI21xp33_ASAP7_75t_L g5153 ( 
.A1(n_5070),
.A2(n_763),
.B(n_764),
.Y(n_5153)
);

XNOR2x1_ASAP7_75t_L g5154 ( 
.A(n_5141),
.B(n_766),
.Y(n_5154)
);

NOR2xp67_ASAP7_75t_L g5155 ( 
.A(n_5068),
.B(n_767),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_5075),
.B(n_767),
.Y(n_5156)
);

INVx2_ASAP7_75t_L g5157 ( 
.A(n_5081),
.Y(n_5157)
);

O2A1O1Ixp33_ASAP7_75t_L g5158 ( 
.A1(n_5055),
.A2(n_770),
.B(n_768),
.C(n_769),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_5064),
.Y(n_5159)
);

AOI22xp5_ASAP7_75t_L g5160 ( 
.A1(n_5120),
.A2(n_774),
.B1(n_770),
.B2(n_772),
.Y(n_5160)
);

INVxp67_ASAP7_75t_L g5161 ( 
.A(n_5057),
.Y(n_5161)
);

AND2x2_ASAP7_75t_L g5162 ( 
.A(n_5060),
.B(n_5137),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_5119),
.Y(n_5163)
);

AOI22x1_ASAP7_75t_L g5164 ( 
.A1(n_5091),
.A2(n_775),
.B1(n_772),
.B2(n_774),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5104),
.Y(n_5165)
);

OAI22xp5_ASAP7_75t_L g5166 ( 
.A1(n_5077),
.A2(n_778),
.B1(n_775),
.B2(n_776),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_5111),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_5071),
.Y(n_5168)
);

XNOR2x1_ASAP7_75t_L g5169 ( 
.A(n_5078),
.B(n_5136),
.Y(n_5169)
);

AOI211xp5_ASAP7_75t_L g5170 ( 
.A1(n_5087),
.A2(n_780),
.B(n_776),
.C(n_779),
.Y(n_5170)
);

OAI222xp33_ASAP7_75t_L g5171 ( 
.A1(n_5082),
.A2(n_782),
.B1(n_784),
.B2(n_780),
.C1(n_781),
.C2(n_783),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_5117),
.Y(n_5172)
);

NOR3xp33_ASAP7_75t_L g5173 ( 
.A(n_5097),
.B(n_781),
.C(n_782),
.Y(n_5173)
);

XNOR2xp5_ASAP7_75t_L g5174 ( 
.A(n_5061),
.B(n_783),
.Y(n_5174)
);

NAND2xp5_ASAP7_75t_L g5175 ( 
.A(n_5103),
.B(n_784),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_5113),
.B(n_785),
.Y(n_5176)
);

INVxp67_ASAP7_75t_L g5177 ( 
.A(n_5058),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_L g5178 ( 
.A(n_5139),
.B(n_785),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_5065),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_5140),
.B(n_786),
.Y(n_5180)
);

INVx1_ASAP7_75t_SL g5181 ( 
.A(n_5128),
.Y(n_5181)
);

A2O1A1Ixp33_ASAP7_75t_L g5182 ( 
.A1(n_5088),
.A2(n_788),
.B(n_786),
.C(n_787),
.Y(n_5182)
);

AOI211xp5_ASAP7_75t_L g5183 ( 
.A1(n_5115),
.A2(n_790),
.B(n_788),
.C(n_789),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_5085),
.B(n_791),
.Y(n_5184)
);

NOR2x1_ASAP7_75t_L g5185 ( 
.A(n_5067),
.B(n_792),
.Y(n_5185)
);

BUFx6f_ASAP7_75t_L g5186 ( 
.A(n_5092),
.Y(n_5186)
);

INVx1_ASAP7_75t_SL g5187 ( 
.A(n_5059),
.Y(n_5187)
);

CKINVDCx8_ASAP7_75t_R g5188 ( 
.A(n_5084),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_5096),
.B(n_792),
.Y(n_5189)
);

INVx2_ASAP7_75t_L g5190 ( 
.A(n_5094),
.Y(n_5190)
);

OR2x2_ASAP7_75t_L g5191 ( 
.A(n_5112),
.B(n_793),
.Y(n_5191)
);

AOI22xp33_ASAP7_75t_L g5192 ( 
.A1(n_5134),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_5192)
);

AOI22xp5_ASAP7_75t_L g5193 ( 
.A1(n_5131),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_5193)
);

XOR2x2_ASAP7_75t_L g5194 ( 
.A(n_5126),
.B(n_798),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5110),
.Y(n_5195)
);

NAND4xp75_ASAP7_75t_L g5196 ( 
.A(n_5108),
.B(n_800),
.C(n_798),
.D(n_799),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_5114),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5121),
.Y(n_5198)
);

O2A1O1Ixp33_ASAP7_75t_L g5199 ( 
.A1(n_5100),
.A2(n_5109),
.B(n_5118),
.C(n_5123),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_5080),
.B(n_800),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_5129),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_5099),
.Y(n_5202)
);

INVx2_ASAP7_75t_L g5203 ( 
.A(n_5122),
.Y(n_5203)
);

XNOR2xp5_ASAP7_75t_L g5204 ( 
.A(n_5063),
.B(n_801),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_5093),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_5086),
.Y(n_5206)
);

AND2x2_ASAP7_75t_L g5207 ( 
.A(n_5102),
.B(n_802),
.Y(n_5207)
);

NOR2xp33_ASAP7_75t_L g5208 ( 
.A(n_5089),
.B(n_803),
.Y(n_5208)
);

OAI21x1_ASAP7_75t_SL g5209 ( 
.A1(n_5135),
.A2(n_804),
.B(n_805),
.Y(n_5209)
);

AOI21xp5_ASAP7_75t_L g5210 ( 
.A1(n_5066),
.A2(n_804),
.B(n_806),
.Y(n_5210)
);

OAI22xp5_ASAP7_75t_L g5211 ( 
.A1(n_5134),
.A2(n_808),
.B1(n_806),
.B2(n_807),
.Y(n_5211)
);

NOR2x1_ASAP7_75t_L g5212 ( 
.A(n_5069),
.B(n_807),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5079),
.Y(n_5213)
);

NAND5xp2_ASAP7_75t_L g5214 ( 
.A(n_5095),
.B(n_811),
.C(n_808),
.D(n_809),
.E(n_812),
.Y(n_5214)
);

AOI22xp33_ASAP7_75t_L g5215 ( 
.A1(n_5130),
.A2(n_817),
.B1(n_814),
.B2(n_816),
.Y(n_5215)
);

AOI22xp5_ASAP7_75t_L g5216 ( 
.A1(n_5090),
.A2(n_817),
.B1(n_814),
.B2(n_816),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_5125),
.B(n_818),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_5062),
.Y(n_5218)
);

NAND2xp5_ASAP7_75t_L g5219 ( 
.A(n_5207),
.B(n_5124),
.Y(n_5219)
);

OAI22xp5_ASAP7_75t_L g5220 ( 
.A1(n_5192),
.A2(n_5132),
.B1(n_5106),
.B2(n_5133),
.Y(n_5220)
);

NOR3xp33_ASAP7_75t_L g5221 ( 
.A(n_5152),
.B(n_5105),
.C(n_5101),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_5164),
.Y(n_5222)
);

NOR2x1_ASAP7_75t_L g5223 ( 
.A(n_5196),
.B(n_818),
.Y(n_5223)
);

NOR3xp33_ASAP7_75t_L g5224 ( 
.A(n_5206),
.B(n_827),
.C(n_819),
.Y(n_5224)
);

NOR2x1p5_ASAP7_75t_SL g5225 ( 
.A(n_5157),
.B(n_819),
.Y(n_5225)
);

NAND5xp2_ASAP7_75t_L g5226 ( 
.A(n_5199),
.B(n_822),
.C(n_820),
.D(n_821),
.E(n_823),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_5150),
.B(n_821),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5174),
.Y(n_5228)
);

NOR2xp33_ASAP7_75t_SL g5229 ( 
.A(n_5171),
.B(n_822),
.Y(n_5229)
);

NOR2x1_ASAP7_75t_L g5230 ( 
.A(n_5214),
.B(n_823),
.Y(n_5230)
);

NAND4xp75_ASAP7_75t_L g5231 ( 
.A(n_5212),
.B(n_826),
.C(n_824),
.D(n_825),
.Y(n_5231)
);

NOR3xp33_ASAP7_75t_L g5232 ( 
.A(n_5205),
.B(n_834),
.C(n_824),
.Y(n_5232)
);

NOR2xp33_ASAP7_75t_L g5233 ( 
.A(n_5153),
.B(n_825),
.Y(n_5233)
);

NOR3xp33_ASAP7_75t_L g5234 ( 
.A(n_5149),
.B(n_837),
.C(n_826),
.Y(n_5234)
);

NAND3xp33_ASAP7_75t_L g5235 ( 
.A(n_5170),
.B(n_827),
.C(n_828),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_5204),
.Y(n_5236)
);

NOR3xp33_ASAP7_75t_L g5237 ( 
.A(n_5146),
.B(n_841),
.C(n_828),
.Y(n_5237)
);

NAND4xp75_ASAP7_75t_L g5238 ( 
.A(n_5185),
.B(n_833),
.C(n_829),
.D(n_832),
.Y(n_5238)
);

AO22x2_ASAP7_75t_L g5239 ( 
.A1(n_5154),
.A2(n_835),
.B1(n_832),
.B2(n_834),
.Y(n_5239)
);

NOR2x1_ASAP7_75t_L g5240 ( 
.A(n_5175),
.B(n_837),
.Y(n_5240)
);

HB1xp67_ASAP7_75t_L g5241 ( 
.A(n_5169),
.Y(n_5241)
);

NOR2x1_ASAP7_75t_L g5242 ( 
.A(n_5156),
.B(n_840),
.Y(n_5242)
);

OA21x2_ASAP7_75t_L g5243 ( 
.A1(n_5143),
.A2(n_841),
.B(n_842),
.Y(n_5243)
);

NOR2x1p5_ASAP7_75t_L g5244 ( 
.A(n_5144),
.B(n_842),
.Y(n_5244)
);

OR2x2_ASAP7_75t_L g5245 ( 
.A(n_5176),
.B(n_843),
.Y(n_5245)
);

NOR2x1_ASAP7_75t_L g5246 ( 
.A(n_5211),
.B(n_844),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_5186),
.Y(n_5247)
);

AND2x2_ASAP7_75t_L g5248 ( 
.A(n_5162),
.B(n_845),
.Y(n_5248)
);

OAI322xp33_ASAP7_75t_L g5249 ( 
.A1(n_5187),
.A2(n_851),
.A3(n_850),
.B1(n_847),
.B2(n_845),
.C1(n_846),
.C2(n_849),
.Y(n_5249)
);

NAND3xp33_ASAP7_75t_L g5250 ( 
.A(n_5145),
.B(n_847),
.C(n_850),
.Y(n_5250)
);

NOR2xp67_ASAP7_75t_L g5251 ( 
.A(n_5210),
.B(n_852),
.Y(n_5251)
);

HB1xp67_ASAP7_75t_L g5252 ( 
.A(n_5186),
.Y(n_5252)
);

NAND3xp33_ASAP7_75t_L g5253 ( 
.A(n_5151),
.B(n_851),
.C(n_852),
.Y(n_5253)
);

NAND3xp33_ASAP7_75t_L g5254 ( 
.A(n_5183),
.B(n_854),
.C(n_855),
.Y(n_5254)
);

NAND3xp33_ASAP7_75t_L g5255 ( 
.A(n_5186),
.B(n_854),
.C(n_855),
.Y(n_5255)
);

NAND4xp25_ASAP7_75t_L g5256 ( 
.A(n_5147),
.B(n_860),
.C(n_856),
.D(n_859),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_5208),
.B(n_856),
.Y(n_5257)
);

INVx2_ASAP7_75t_L g5258 ( 
.A(n_5209),
.Y(n_5258)
);

NAND3xp33_ASAP7_75t_L g5259 ( 
.A(n_5158),
.B(n_859),
.C(n_860),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_5160),
.B(n_861),
.Y(n_5260)
);

A2O1A1Ixp33_ASAP7_75t_L g5261 ( 
.A1(n_5155),
.A2(n_863),
.B(n_861),
.C(n_862),
.Y(n_5261)
);

NAND4xp25_ASAP7_75t_L g5262 ( 
.A(n_5218),
.B(n_868),
.C(n_865),
.D(n_866),
.Y(n_5262)
);

NOR2x1_ASAP7_75t_L g5263 ( 
.A(n_5191),
.B(n_865),
.Y(n_5263)
);

NOR2x1_ASAP7_75t_L g5264 ( 
.A(n_5178),
.B(n_866),
.Y(n_5264)
);

OA22x2_ASAP7_75t_L g5265 ( 
.A1(n_5216),
.A2(n_871),
.B1(n_869),
.B2(n_870),
.Y(n_5265)
);

AND2x2_ASAP7_75t_L g5266 ( 
.A(n_5165),
.B(n_869),
.Y(n_5266)
);

NAND3xp33_ASAP7_75t_L g5267 ( 
.A(n_5182),
.B(n_870),
.C(n_871),
.Y(n_5267)
);

AOI22xp5_ASAP7_75t_L g5268 ( 
.A1(n_5181),
.A2(n_875),
.B1(n_872),
.B2(n_874),
.Y(n_5268)
);

NOR2x1_ASAP7_75t_L g5269 ( 
.A(n_5180),
.B(n_5200),
.Y(n_5269)
);

NOR2x1_ASAP7_75t_L g5270 ( 
.A(n_5163),
.B(n_872),
.Y(n_5270)
);

NOR3xp33_ASAP7_75t_L g5271 ( 
.A(n_5213),
.B(n_882),
.C(n_874),
.Y(n_5271)
);

OAI21xp33_ASAP7_75t_SL g5272 ( 
.A1(n_5184),
.A2(n_875),
.B(n_876),
.Y(n_5272)
);

NOR2x1_ASAP7_75t_SL g5273 ( 
.A(n_5166),
.B(n_876),
.Y(n_5273)
);

AND2x2_ASAP7_75t_L g5274 ( 
.A(n_5168),
.B(n_877),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_5225),
.Y(n_5275)
);

OAI22xp5_ASAP7_75t_L g5276 ( 
.A1(n_5247),
.A2(n_5188),
.B1(n_5217),
.B2(n_5189),
.Y(n_5276)
);

HB1xp67_ASAP7_75t_L g5277 ( 
.A(n_5243),
.Y(n_5277)
);

O2A1O1Ixp33_ASAP7_75t_SL g5278 ( 
.A1(n_5252),
.A2(n_5172),
.B(n_5167),
.C(n_5161),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5239),
.Y(n_5279)
);

INVx2_ASAP7_75t_L g5280 ( 
.A(n_5243),
.Y(n_5280)
);

O2A1O1Ixp5_ASAP7_75t_L g5281 ( 
.A1(n_5227),
.A2(n_5203),
.B(n_5190),
.C(n_5198),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5239),
.Y(n_5282)
);

NAND4xp75_ASAP7_75t_L g5283 ( 
.A(n_5240),
.B(n_5202),
.C(n_5201),
.D(n_5159),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_5248),
.Y(n_5284)
);

CKINVDCx20_ASAP7_75t_R g5285 ( 
.A(n_5241),
.Y(n_5285)
);

INVx1_ASAP7_75t_SL g5286 ( 
.A(n_5231),
.Y(n_5286)
);

NAND2xp5_ASAP7_75t_L g5287 ( 
.A(n_5266),
.B(n_5173),
.Y(n_5287)
);

OR2x2_ASAP7_75t_L g5288 ( 
.A(n_5226),
.B(n_5194),
.Y(n_5288)
);

OAI22xp33_ASAP7_75t_L g5289 ( 
.A1(n_5229),
.A2(n_5193),
.B1(n_5177),
.B2(n_5197),
.Y(n_5289)
);

CKINVDCx16_ASAP7_75t_R g5290 ( 
.A(n_5230),
.Y(n_5290)
);

NOR4xp75_ASAP7_75t_L g5291 ( 
.A(n_5238),
.B(n_5142),
.C(n_5195),
.D(n_5179),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5270),
.Y(n_5292)
);

NAND4xp25_ASAP7_75t_L g5293 ( 
.A(n_5237),
.B(n_5215),
.C(n_5148),
.D(n_879),
.Y(n_5293)
);

NAND3xp33_ASAP7_75t_L g5294 ( 
.A(n_5234),
.B(n_877),
.C(n_878),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5274),
.Y(n_5295)
);

A2O1A1Ixp33_ASAP7_75t_L g5296 ( 
.A1(n_5233),
.A2(n_880),
.B(n_878),
.C(n_879),
.Y(n_5296)
);

CKINVDCx20_ASAP7_75t_R g5297 ( 
.A(n_5228),
.Y(n_5297)
);

NAND3xp33_ASAP7_75t_SL g5298 ( 
.A(n_5261),
.B(n_880),
.C(n_881),
.Y(n_5298)
);

AOI22xp5_ASAP7_75t_L g5299 ( 
.A1(n_5221),
.A2(n_883),
.B1(n_881),
.B2(n_882),
.Y(n_5299)
);

OAI22xp33_ASAP7_75t_L g5300 ( 
.A1(n_5222),
.A2(n_885),
.B1(n_883),
.B2(n_884),
.Y(n_5300)
);

INVx1_ASAP7_75t_SL g5301 ( 
.A(n_5223),
.Y(n_5301)
);

AOI22xp33_ASAP7_75t_L g5302 ( 
.A1(n_5244),
.A2(n_886),
.B1(n_884),
.B2(n_885),
.Y(n_5302)
);

OAI21xp33_ASAP7_75t_SL g5303 ( 
.A1(n_5251),
.A2(n_886),
.B(n_887),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_5265),
.Y(n_5304)
);

CKINVDCx6p67_ASAP7_75t_R g5305 ( 
.A(n_5236),
.Y(n_5305)
);

AOI21x1_ASAP7_75t_L g5306 ( 
.A1(n_5263),
.A2(n_887),
.B(n_888),
.Y(n_5306)
);

OAI31xp33_ASAP7_75t_L g5307 ( 
.A1(n_5250),
.A2(n_891),
.A3(n_889),
.B(n_890),
.Y(n_5307)
);

AOI21xp33_ASAP7_75t_L g5308 ( 
.A1(n_5245),
.A2(n_889),
.B(n_890),
.Y(n_5308)
);

XOR2x2_ASAP7_75t_L g5309 ( 
.A(n_5259),
.B(n_891),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5277),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_L g5311 ( 
.A(n_5275),
.B(n_5232),
.Y(n_5311)
);

NAND3xp33_ASAP7_75t_L g5312 ( 
.A(n_5307),
.B(n_5242),
.C(n_5264),
.Y(n_5312)
);

AND2x4_ASAP7_75t_L g5313 ( 
.A(n_5285),
.B(n_5258),
.Y(n_5313)
);

AND2x2_ASAP7_75t_L g5314 ( 
.A(n_5290),
.B(n_5273),
.Y(n_5314)
);

BUFx2_ASAP7_75t_L g5315 ( 
.A(n_5303),
.Y(n_5315)
);

OAI22xp33_ASAP7_75t_L g5316 ( 
.A1(n_5301),
.A2(n_5256),
.B1(n_5260),
.B2(n_5257),
.Y(n_5316)
);

OR5x1_ASAP7_75t_L g5317 ( 
.A(n_5293),
.B(n_5262),
.C(n_5272),
.D(n_5220),
.E(n_5253),
.Y(n_5317)
);

NOR2xp67_ASAP7_75t_L g5318 ( 
.A(n_5280),
.B(n_5255),
.Y(n_5318)
);

AND2x2_ASAP7_75t_L g5319 ( 
.A(n_5284),
.B(n_5246),
.Y(n_5319)
);

INVxp67_ASAP7_75t_SL g5320 ( 
.A(n_5306),
.Y(n_5320)
);

NAND5xp2_ASAP7_75t_L g5321 ( 
.A(n_5304),
.B(n_5219),
.C(n_5224),
.D(n_5271),
.E(n_5268),
.Y(n_5321)
);

NOR3xp33_ASAP7_75t_SL g5322 ( 
.A(n_5289),
.B(n_5235),
.C(n_5254),
.Y(n_5322)
);

NAND2x1p5_ASAP7_75t_L g5323 ( 
.A(n_5292),
.B(n_5269),
.Y(n_5323)
);

NAND4xp75_ASAP7_75t_L g5324 ( 
.A(n_5281),
.B(n_5267),
.C(n_5249),
.D(n_894),
.Y(n_5324)
);

NAND4xp25_ASAP7_75t_SL g5325 ( 
.A(n_5286),
.B(n_894),
.C(n_892),
.D(n_893),
.Y(n_5325)
);

NOR2xp33_ASAP7_75t_L g5326 ( 
.A(n_5288),
.B(n_892),
.Y(n_5326)
);

NAND2x1p5_ASAP7_75t_SL g5327 ( 
.A(n_5305),
.B(n_895),
.Y(n_5327)
);

OAI221xp5_ASAP7_75t_SL g5328 ( 
.A1(n_5311),
.A2(n_5279),
.B1(n_5282),
.B2(n_5287),
.C(n_5295),
.Y(n_5328)
);

INVxp67_ASAP7_75t_L g5329 ( 
.A(n_5326),
.Y(n_5329)
);

AOI22xp33_ASAP7_75t_L g5330 ( 
.A1(n_5313),
.A2(n_5297),
.B1(n_5298),
.B2(n_5294),
.Y(n_5330)
);

OAI21xp33_ASAP7_75t_SL g5331 ( 
.A1(n_5320),
.A2(n_5283),
.B(n_5308),
.Y(n_5331)
);

NOR4xp25_ASAP7_75t_L g5332 ( 
.A(n_5310),
.B(n_5278),
.C(n_5276),
.D(n_5296),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_SL g5333 ( 
.A(n_5318),
.B(n_5302),
.Y(n_5333)
);

OAI211xp5_ASAP7_75t_SL g5334 ( 
.A1(n_5322),
.A2(n_5291),
.B(n_5299),
.C(n_5309),
.Y(n_5334)
);

AOI22xp5_ASAP7_75t_L g5335 ( 
.A1(n_5314),
.A2(n_5300),
.B1(n_898),
.B2(n_895),
.Y(n_5335)
);

AOI21xp33_ASAP7_75t_SL g5336 ( 
.A1(n_5327),
.A2(n_896),
.B(n_898),
.Y(n_5336)
);

NOR2xp33_ASAP7_75t_L g5337 ( 
.A(n_5315),
.B(n_899),
.Y(n_5337)
);

AOI21xp5_ASAP7_75t_L g5338 ( 
.A1(n_5312),
.A2(n_900),
.B(n_901),
.Y(n_5338)
);

AOI211xp5_ASAP7_75t_SL g5339 ( 
.A1(n_5328),
.A2(n_5316),
.B(n_5319),
.C(n_5317),
.Y(n_5339)
);

NAND4xp75_ASAP7_75t_L g5340 ( 
.A(n_5331),
.B(n_5337),
.C(n_5333),
.D(n_5338),
.Y(n_5340)
);

NOR2x2_ASAP7_75t_L g5341 ( 
.A(n_5336),
.B(n_5324),
.Y(n_5341)
);

NAND5xp2_ASAP7_75t_L g5342 ( 
.A(n_5330),
.B(n_5323),
.C(n_5321),
.D(n_5325),
.E(n_903),
.Y(n_5342)
);

OR2x2_ASAP7_75t_L g5343 ( 
.A(n_5332),
.B(n_900),
.Y(n_5343)
);

OAI221xp5_ASAP7_75t_L g5344 ( 
.A1(n_5335),
.A2(n_905),
.B1(n_902),
.B2(n_904),
.C(n_907),
.Y(n_5344)
);

NOR2x1p5_ASAP7_75t_L g5345 ( 
.A(n_5334),
.B(n_905),
.Y(n_5345)
);

NOR2x1_ASAP7_75t_L g5346 ( 
.A(n_5343),
.B(n_5329),
.Y(n_5346)
);

OR2x2_ASAP7_75t_L g5347 ( 
.A(n_5342),
.B(n_908),
.Y(n_5347)
);

OAI21xp5_ASAP7_75t_L g5348 ( 
.A1(n_5339),
.A2(n_908),
.B(n_909),
.Y(n_5348)
);

OAI22xp5_ASAP7_75t_L g5349 ( 
.A1(n_5344),
.A2(n_912),
.B1(n_910),
.B2(n_911),
.Y(n_5349)
);

OR2x2_ASAP7_75t_L g5350 ( 
.A(n_5345),
.B(n_5340),
.Y(n_5350)
);

XOR2x1_ASAP7_75t_L g5351 ( 
.A(n_5347),
.B(n_5341),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5348),
.Y(n_5352)
);

NAND2x1_ASAP7_75t_L g5353 ( 
.A(n_5352),
.B(n_5346),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5353),
.Y(n_5354)
);

OAI22xp5_ASAP7_75t_SL g5355 ( 
.A1(n_5354),
.A2(n_5350),
.B1(n_5349),
.B2(n_5351),
.Y(n_5355)
);

INVx4_ASAP7_75t_L g5356 ( 
.A(n_5355),
.Y(n_5356)
);

INVxp67_ASAP7_75t_L g5357 ( 
.A(n_5356),
.Y(n_5357)
);

OAI21xp33_ASAP7_75t_SL g5358 ( 
.A1(n_5357),
.A2(n_910),
.B(n_912),
.Y(n_5358)
);

XNOR2xp5_ASAP7_75t_L g5359 ( 
.A(n_5358),
.B(n_913),
.Y(n_5359)
);

AOI22xp5_ASAP7_75t_L g5360 ( 
.A1(n_5359),
.A2(n_915),
.B1(n_913),
.B2(n_914),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5360),
.Y(n_5361)
);

OR2x6_ASAP7_75t_L g5362 ( 
.A(n_5361),
.B(n_915),
.Y(n_5362)
);

AOI22xp33_ASAP7_75t_SL g5363 ( 
.A1(n_5362),
.A2(n_918),
.B1(n_916),
.B2(n_917),
.Y(n_5363)
);

AOI211xp5_ASAP7_75t_L g5364 ( 
.A1(n_5363),
.A2(n_919),
.B(n_917),
.C(n_918),
.Y(n_5364)
);


endmodule