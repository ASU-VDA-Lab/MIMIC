module real_aes_2994_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_0), .B(n_480), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_1), .A2(n_482), .B(n_483), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_2), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_3), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_4), .B(n_241), .Y(n_515) );
INVx1_ASAP7_75t_L g127 ( .A(n_5), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_6), .B(n_146), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_7), .B(n_241), .Y(n_542) );
INVx1_ASAP7_75t_L g210 ( .A(n_8), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g778 ( .A(n_9), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_10), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g504 ( .A(n_11), .B(n_238), .Y(n_504) );
INVx2_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
AOI221x1_ASAP7_75t_L g548 ( .A1(n_13), .A2(n_25), .B1(n_480), .B2(n_482), .C(n_549), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_14), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_15), .B(n_480), .Y(n_500) );
INVx1_ASAP7_75t_L g239 ( .A(n_16), .Y(n_239) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_17), .A2(n_191), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_18), .B(n_150), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_19), .B(n_241), .Y(n_492) );
AO21x1_ASAP7_75t_L g510 ( .A1(n_20), .A2(n_480), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g466 ( .A(n_21), .Y(n_466) );
INVx1_ASAP7_75t_L g236 ( .A(n_22), .Y(n_236) );
INVx1_ASAP7_75t_SL g156 ( .A(n_23), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_24), .B(n_133), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_26), .Y(n_767) );
AOI33xp33_ASAP7_75t_L g196 ( .A1(n_27), .A2(n_53), .A3(n_122), .B1(n_131), .B2(n_197), .B3(n_198), .Y(n_196) );
NAND2x1_ASAP7_75t_L g523 ( .A(n_28), .B(n_241), .Y(n_523) );
NAND2x1_ASAP7_75t_L g541 ( .A(n_29), .B(n_238), .Y(n_541) );
INVx1_ASAP7_75t_L g167 ( .A(n_30), .Y(n_167) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_31), .A2(n_85), .B(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g147 ( .A(n_31), .B(n_85), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_32), .B(n_141), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_33), .B(n_238), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_34), .B(n_241), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_35), .B(n_238), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_36), .A2(n_482), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
AND2x2_ASAP7_75t_L g139 ( .A(n_37), .B(n_127), .Y(n_139) );
AND2x2_ASAP7_75t_L g145 ( .A(n_37), .B(n_124), .Y(n_145) );
OR2x6_ASAP7_75t_L g464 ( .A(n_38), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_39), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_40), .B(n_480), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_41), .B(n_141), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_42), .A2(n_114), .B1(n_146), .B2(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_43), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_44), .B(n_133), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_45), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_46), .B(n_238), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_47), .B(n_191), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_48), .B(n_133), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_49), .A2(n_482), .B(n_540), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_50), .Y(n_223) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_51), .A2(n_100), .B1(n_763), .B2(n_764), .C1(n_767), .C2(n_768), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_51), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_52), .B(n_238), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_54), .B(n_133), .Y(n_186) );
INVx1_ASAP7_75t_L g126 ( .A(n_55), .Y(n_126) );
INVx1_ASAP7_75t_L g135 ( .A(n_55), .Y(n_135) );
AND2x2_ASAP7_75t_L g187 ( .A(n_56), .B(n_150), .Y(n_187) );
AOI221xp5_ASAP7_75t_L g208 ( .A1(n_57), .A2(n_73), .B1(n_119), .B2(n_141), .C(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_58), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_59), .B(n_241), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_60), .B(n_114), .Y(n_177) );
AOI21xp5_ASAP7_75t_SL g118 ( .A1(n_61), .A2(n_119), .B(n_128), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_62), .A2(n_482), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g233 ( .A(n_63), .Y(n_233) );
AO21x1_ASAP7_75t_L g512 ( .A1(n_64), .A2(n_482), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_65), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g185 ( .A(n_66), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_67), .B(n_480), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_68), .A2(n_119), .B(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g534 ( .A(n_69), .B(n_151), .Y(n_534) );
INVx1_ASAP7_75t_L g124 ( .A(n_70), .Y(n_124) );
INVx1_ASAP7_75t_L g137 ( .A(n_70), .Y(n_137) );
AND2x2_ASAP7_75t_L g544 ( .A(n_71), .B(n_113), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_72), .B(n_141), .Y(n_199) );
AND2x2_ASAP7_75t_L g158 ( .A(n_74), .B(n_113), .Y(n_158) );
INVx1_ASAP7_75t_L g234 ( .A(n_75), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_76), .A2(n_119), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_77), .A2(n_119), .B(n_190), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g467 ( .A(n_78), .Y(n_467) );
AND2x2_ASAP7_75t_L g477 ( .A(n_79), .B(n_113), .Y(n_477) );
AND2x2_ASAP7_75t_SL g112 ( .A(n_80), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_81), .B(n_480), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_82), .A2(n_99), .B1(n_772), .B2(n_782), .C1(n_794), .C2(n_798), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g784 ( .A1(n_82), .A2(n_468), .B1(n_785), .B2(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_82), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_83), .A2(n_119), .B1(n_194), .B2(n_195), .Y(n_193) );
AND2x2_ASAP7_75t_L g511 ( .A(n_84), .B(n_146), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_86), .B(n_238), .Y(n_493) );
AND2x2_ASAP7_75t_L g526 ( .A(n_87), .B(n_113), .Y(n_526) );
INVx1_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_89), .B(n_241), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_90), .A2(n_482), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_91), .B(n_238), .Y(n_550) );
AND2x2_ASAP7_75t_L g200 ( .A(n_92), .B(n_113), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_93), .B(n_241), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_94), .A2(n_165), .B(n_166), .C(n_169), .Y(n_164) );
BUFx2_ASAP7_75t_L g779 ( .A(n_95), .Y(n_779) );
BUFx2_ASAP7_75t_SL g802 ( .A(n_95), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_96), .A2(n_482), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_97), .B(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_459), .B1(n_468), .B2(n_761), .Y(n_101) );
AOI22x1_ASAP7_75t_L g768 ( .A1(n_102), .A2(n_460), .B1(n_769), .B2(n_771), .Y(n_768) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
AND3x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_349), .C(n_412), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_313), .Y(n_105) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_254), .C(n_283), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_243), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_159), .B1(n_201), .B2(n_213), .Y(n_108) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_109), .B(n_244), .Y(n_398) );
INVx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_148), .Y(n_110) );
INVx2_ASAP7_75t_L g215 ( .A(n_111), .Y(n_215) );
INVx4_ASAP7_75t_L g259 ( .A(n_111), .Y(n_259) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_111), .Y(n_279) );
AND2x4_ASAP7_75t_L g290 ( .A(n_111), .B(n_258), .Y(n_290) );
AND2x2_ASAP7_75t_L g296 ( .A(n_111), .B(n_218), .Y(n_296) );
NOR2x1_ASAP7_75t_SL g426 ( .A(n_111), .B(n_229), .Y(n_426) );
OR2x6_ASAP7_75t_L g111 ( .A(n_112), .B(n_117), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_113), .A2(n_164), .B1(n_170), .B2(n_171), .Y(n_163) );
INVx3_ASAP7_75t_L g171 ( .A(n_113), .Y(n_171) );
INVx4_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_114), .B(n_174), .Y(n_173) );
INVx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_115), .Y(n_191) );
AND2x4_ASAP7_75t_L g146 ( .A(n_116), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_116), .B(n_147), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_140), .B(n_146), .Y(n_117) );
INVxp67_ASAP7_75t_L g176 ( .A(n_119), .Y(n_176) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_125), .Y(n_119) );
NOR2x1p5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g198 ( .A(n_122), .Y(n_198) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x6_ASAP7_75t_L g130 ( .A(n_123), .B(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_L g238 ( .A(n_124), .B(n_134), .Y(n_238) );
AND2x6_ASAP7_75t_L g482 ( .A(n_125), .B(n_145), .Y(n_482) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
INVx2_ASAP7_75t_L g131 ( .A(n_126), .Y(n_131) );
AND2x4_ASAP7_75t_L g241 ( .A(n_126), .B(n_136), .Y(n_241) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_127), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_132), .C(n_138), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_SL g155 ( .A1(n_130), .A2(n_138), .B(n_156), .C(n_157), .Y(n_155) );
INVxp67_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_130), .A2(n_138), .B(n_185), .C(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_SL g209 ( .A1(n_130), .A2(n_138), .B(n_210), .C(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g228 ( .A(n_130), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_130), .A2(n_168), .B1(n_233), .B2(n_234), .Y(n_232) );
AND2x2_ASAP7_75t_L g142 ( .A(n_131), .B(n_143), .Y(n_142) );
INVxp33_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
INVx1_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
AND2x4_ASAP7_75t_L g480 ( .A(n_133), .B(n_139), .Y(n_480) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g194 ( .A(n_138), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_138), .A2(n_226), .B(n_227), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_138), .B(n_146), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_138), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_138), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_138), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_138), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_138), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_138), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_138), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_138), .A2(n_550), .B(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
INVx1_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_144), .Y(n_222) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_SL g488 ( .A(n_146), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_146), .A2(n_500), .B(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_146), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g262 ( .A(n_148), .Y(n_262) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_148), .Y(n_276) );
INVx1_ASAP7_75t_L g287 ( .A(n_148), .Y(n_287) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_148), .Y(n_299) );
AND2x2_ASAP7_75t_L g331 ( .A(n_148), .B(n_229), .Y(n_331) );
AND2x2_ASAP7_75t_L g363 ( .A(n_148), .B(n_247), .Y(n_363) );
INVx1_ASAP7_75t_L g370 ( .A(n_148), .Y(n_370) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_158), .Y(n_148) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_149), .A2(n_538), .B(n_544), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_150), .A2(n_479), .B(n_481), .Y(n_478) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_150), .A2(n_548), .B(n_552), .Y(n_547) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_150), .A2(n_548), .B(n_552), .Y(n_587) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_179), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g312 ( .A(n_161), .B(n_251), .Y(n_312) );
INVx2_ASAP7_75t_L g386 ( .A(n_161), .Y(n_386) );
AND2x2_ASAP7_75t_L g409 ( .A(n_161), .B(n_179), .Y(n_409) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_162), .B(n_204), .Y(n_250) );
INVx2_ASAP7_75t_L g271 ( .A(n_162), .Y(n_271) );
AND2x4_ASAP7_75t_L g293 ( .A(n_162), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g328 ( .A(n_162), .Y(n_328) );
AND2x2_ASAP7_75t_L g405 ( .A(n_162), .B(n_207), .Y(n_405) );
OR2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_172), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_171), .A2(n_181), .B(n_187), .Y(n_180) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_181), .B(n_187), .Y(n_204) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_171), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_171), .A2(n_528), .B(n_534), .Y(n_527) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_171), .A2(n_520), .B(n_526), .Y(n_555) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_171), .A2(n_528), .B(n_534), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g376 ( .A(n_179), .Y(n_376) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_188), .Y(n_179) );
NOR2xp67_ASAP7_75t_L g301 ( .A(n_180), .B(n_271), .Y(n_301) );
AND2x2_ASAP7_75t_L g306 ( .A(n_180), .B(n_271), .Y(n_306) );
INVx2_ASAP7_75t_L g319 ( .A(n_180), .Y(n_319) );
NOR2x1_ASAP7_75t_L g367 ( .A(n_180), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
AND2x4_ASAP7_75t_L g292 ( .A(n_188), .B(n_203), .Y(n_292) );
AND2x2_ASAP7_75t_L g307 ( .A(n_188), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g360 ( .A(n_188), .Y(n_360) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_189), .B(n_207), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_189), .B(n_204), .Y(n_364) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B(n_200), .Y(n_189) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_190), .A2(n_192), .B(n_200), .Y(n_253) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_191), .A2(n_208), .B(n_212), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_193), .B(n_199), .Y(n_192) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVxp33_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_203), .B(n_205), .Y(n_202) );
INVx3_ASAP7_75t_L g268 ( .A(n_203), .Y(n_268) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
AND2x2_ASAP7_75t_L g435 ( .A(n_204), .B(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g323 ( .A(n_205), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_205), .B(n_360), .Y(n_455) );
BUFx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g270 ( .A(n_206), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g251 ( .A(n_207), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g294 ( .A(n_207), .Y(n_294) );
INVxp67_ASAP7_75t_L g308 ( .A(n_207), .Y(n_308) );
INVx1_ASAP7_75t_L g368 ( .A(n_207), .Y(n_368) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_207), .Y(n_436) );
INVx1_ASAP7_75t_L g420 ( .A(n_213), .Y(n_420) );
NOR2x1_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
NOR2x1_ASAP7_75t_L g340 ( .A(n_214), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g374 ( .A(n_215), .B(n_246), .Y(n_374) );
OR2x2_ASAP7_75t_L g410 ( .A(n_216), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g392 ( .A(n_217), .B(n_370), .Y(n_392) );
AND2x2_ASAP7_75t_L g444 ( .A(n_217), .B(n_279), .Y(n_444) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_229), .Y(n_217) );
AND2x4_ASAP7_75t_L g246 ( .A(n_218), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
INVx2_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_218), .Y(n_453) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_224), .Y(n_218) );
NOR3xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .C(n_223), .Y(n_220) );
INVx3_ASAP7_75t_L g247 ( .A(n_229), .Y(n_247) );
INVx2_ASAP7_75t_L g341 ( .A(n_229), .Y(n_341) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_235), .B(n_242), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_239), .B2(n_240), .Y(n_235) );
INVxp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVxp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_245), .B(n_321), .Y(n_338) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_245), .B(n_259), .Y(n_380) );
INVx4_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_246), .B(n_321), .Y(n_458) );
AND2x2_ASAP7_75t_L g274 ( .A(n_247), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g288 ( .A(n_247), .Y(n_288) );
AOI22xp5_ASAP7_75t_SL g336 ( .A1(n_248), .A2(n_337), .B1(n_338), .B2(n_339), .Y(n_336) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_249), .B(n_307), .Y(n_333) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g394 ( .A(n_250), .B(n_282), .Y(n_394) );
AND2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g300 ( .A(n_251), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g396 ( .A(n_251), .B(n_386), .Y(n_396) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g318 ( .A(n_253), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g344 ( .A(n_253), .Y(n_344) );
AND2x2_ASAP7_75t_L g434 ( .A(n_253), .B(n_271), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_263), .B1(n_267), .B2(n_272), .C(n_277), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g335 ( .A(n_257), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_257), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_257), .B(n_331), .Y(n_450) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NOR2xp67_ASAP7_75t_SL g303 ( .A(n_259), .B(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_259), .Y(n_316) );
OR2x2_ASAP7_75t_L g400 ( .A(n_259), .B(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_259), .B(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g321 ( .A(n_261), .Y(n_321) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_262), .Y(n_411) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI221x1_ASAP7_75t_L g351 ( .A1(n_264), .A2(n_352), .B1(n_354), .B2(n_357), .C(n_361), .Y(n_351) );
AND2x2_ASAP7_75t_L g337 ( .A(n_265), .B(n_293), .Y(n_337) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g280 ( .A(n_268), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_268), .B(n_270), .Y(n_407) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
AND2x2_ASAP7_75t_SL g278 ( .A(n_274), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_274), .B(n_287), .Y(n_304) );
INVx2_ASAP7_75t_L g311 ( .A(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g356 ( .A(n_275), .Y(n_356) );
BUFx2_ASAP7_75t_L g445 ( .A(n_276), .Y(n_445) );
NAND2xp33_ASAP7_75t_SL g277 ( .A(n_278), .B(n_280), .Y(n_277) );
OR2x6_ASAP7_75t_L g310 ( .A(n_279), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g391 ( .A(n_279), .B(n_331), .Y(n_391) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_302), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_291), .B1(n_295), .B2(n_300), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_286), .B(n_290), .Y(n_348) );
AND2x4_ASAP7_75t_L g354 ( .A(n_286), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_SL g286 ( .A(n_287), .B(n_288), .Y(n_286) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_287), .Y(n_379) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_290), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_290), .B(n_321), .Y(n_353) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_290), .Y(n_437) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g384 ( .A(n_292), .B(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g345 ( .A(n_293), .Y(n_345) );
NAND2x1_ASAP7_75t_SL g389 ( .A(n_293), .B(n_344), .Y(n_389) );
AND2x2_ASAP7_75t_L g423 ( .A(n_293), .B(n_318), .Y(n_423) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B1(n_309), .B2(n_312), .Y(n_302) );
BUFx2_ASAP7_75t_L g418 ( .A(n_304), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_305), .A2(n_374), .B1(n_448), .B2(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_306), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_311), .B(n_443), .C(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g346 ( .A(n_312), .Y(n_346) );
AOI211x1_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_322), .B(n_324), .C(n_342), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_317), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g404 ( .A(n_318), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_318), .B(n_385), .Y(n_416) );
AND2x2_ASAP7_75t_L g448 ( .A(n_318), .B(n_386), .Y(n_448) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g429 ( .A(n_321), .Y(n_429) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g358 ( .A(n_323), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_336), .Y(n_324) );
AOI22xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_329), .B1(n_332), .B2(n_334), .Y(n_325) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g366 ( .A(n_328), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g381 ( .A(n_328), .Y(n_381) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_331), .B(n_452), .Y(n_451) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g387 ( .A(n_340), .B(n_370), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .B(n_347), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_344), .B(n_366), .Y(n_441) );
OR2x2_ASAP7_75t_L g419 ( .A(n_345), .B(n_364), .Y(n_419) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND3x1_ASAP7_75t_L g350 ( .A(n_351), .B(n_371), .C(n_395), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_354), .A2(n_384), .B1(n_387), .B2(n_388), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_355), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g428 ( .A(n_355), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_355), .B(n_429), .Y(n_432) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI222xp33_ASAP7_75t_L g415 ( .A1(n_359), .A2(n_416), .B1(n_417), .B2(n_418), .C1(n_419), .C2(n_420), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B1(n_365), .B2(n_369), .Y(n_361) );
INVx1_ASAP7_75t_SL g401 ( .A(n_363), .Y(n_401) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g438 ( .A(n_367), .B(n_434), .Y(n_438) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_372), .B(n_382), .Y(n_371) );
AOI21xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_375), .B(n_381), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_389), .B(n_403), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_392), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_399), .B2(n_402), .C(n_406), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
NAND3x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_439), .C(n_446), .Y(n_413) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_421), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_430), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_425), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_437), .B2(n_438), .Y(n_430) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_440), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_456), .Y(n_446) );
AOI22xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_449), .B1(n_451), .B2(n_454), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
CKINVDCx11_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
OR2x6_ASAP7_75t_SL g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x6_ASAP7_75t_SL g762 ( .A(n_462), .B(n_464), .Y(n_762) );
OR2x2_ASAP7_75t_L g766 ( .A(n_462), .B(n_464), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_462), .B(n_463), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g786 ( .A(n_468), .Y(n_786) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g771 ( .A(n_469), .Y(n_771) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_670), .Y(n_469) );
NOR4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_588), .C(n_614), .D(n_654), .Y(n_470) );
OAI211xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_505), .B(n_535), .C(n_574), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
AND2x2_ASAP7_75t_L g741 ( .A(n_474), .B(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_475), .B(n_486), .Y(n_608) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g536 ( .A(n_476), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_476), .B(n_561), .Y(n_560) );
INVx5_ASAP7_75t_L g594 ( .A(n_476), .Y(n_594) );
NOR2x1_ASAP7_75t_SL g636 ( .A(n_476), .B(n_487), .Y(n_636) );
AND2x2_ASAP7_75t_L g692 ( .A(n_476), .B(n_498), .Y(n_692) );
OR2x6_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_497), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_487), .B(n_498), .Y(n_564) );
AND2x2_ASAP7_75t_L g625 ( .A(n_487), .B(n_594), .Y(n_625) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_495), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_488), .B(n_496), .Y(n_495) );
AO21x2_ASAP7_75t_L g578 ( .A1(n_488), .A2(n_489), .B(n_495), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .Y(n_489) );
AND2x2_ASAP7_75t_L g637 ( .A(n_497), .B(n_561), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_497), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g681 ( .A(n_497), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g714 ( .A(n_497), .B(n_536), .Y(n_714) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g558 ( .A(n_498), .Y(n_558) );
AND2x2_ASAP7_75t_L g591 ( .A(n_498), .B(n_592), .Y(n_591) );
BUFx3_ASAP7_75t_L g626 ( .A(n_498), .Y(n_626) );
OR2x2_ASAP7_75t_L g702 ( .A(n_498), .B(n_561), .Y(n_702) );
INVx1_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
AOI211x1_ASAP7_75t_SL g631 ( .A1(n_507), .A2(n_623), .B(n_632), .C(n_634), .Y(n_631) );
AND2x2_ASAP7_75t_SL g676 ( .A(n_507), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_507), .B(n_674), .Y(n_721) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g571 ( .A(n_508), .Y(n_571) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g546 ( .A(n_509), .Y(n_546) );
OAI21x1_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_512), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_L g517 ( .A(n_511), .Y(n_517) );
AOI322xp5_ASAP7_75t_L g535 ( .A1(n_518), .A2(n_536), .A3(n_545), .B1(n_553), .B2(n_556), .C1(n_562), .C2(n_565), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_518), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
INVx2_ASAP7_75t_L g569 ( .A(n_519), .Y(n_569) );
INVxp67_ASAP7_75t_L g611 ( .A(n_519), .Y(n_611) );
BUFx3_ASAP7_75t_L g675 ( .A(n_519), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
INVx2_ASAP7_75t_L g584 ( .A(n_527), .Y(n_584) );
AND2x2_ASAP7_75t_L g633 ( .A(n_527), .B(n_547), .Y(n_633) );
AND2x2_ASAP7_75t_L g677 ( .A(n_527), .B(n_586), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_533), .Y(n_528) );
AND2x2_ASAP7_75t_L g562 ( .A(n_536), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_536), .B(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_536), .B(n_591), .Y(n_756) );
INVx4_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
AND2x2_ASAP7_75t_L g593 ( .A(n_537), .B(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_537), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_545), .B(n_630), .Y(n_655) );
INVx1_ASAP7_75t_SL g694 ( .A(n_545), .Y(n_694) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x4_ASAP7_75t_L g585 ( .A(n_546), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_546), .B(n_584), .Y(n_653) );
AND2x2_ASAP7_75t_L g705 ( .A(n_546), .B(n_555), .Y(n_705) );
OR2x2_ASAP7_75t_L g729 ( .A(n_546), .B(n_547), .Y(n_729) );
AND2x2_ASAP7_75t_L g553 ( .A(n_547), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g603 ( .A(n_547), .B(n_584), .Y(n_603) );
AND2x2_ASAP7_75t_SL g659 ( .A(n_547), .B(n_571), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_553), .B(n_666), .Y(n_683) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g618 ( .A(n_555), .Y(n_618) );
AND2x4_ASAP7_75t_SL g658 ( .A(n_555), .B(n_572), .Y(n_658) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
OR2x2_ASAP7_75t_L g606 ( .A(n_557), .B(n_560), .Y(n_606) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g575 ( .A(n_558), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g723 ( .A(n_558), .B(n_636), .Y(n_723) );
AND2x2_ASAP7_75t_L g739 ( .A(n_558), .B(n_593), .Y(n_739) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI311xp33_ASAP7_75t_L g709 ( .A1(n_560), .A2(n_648), .A3(n_710), .B(n_712), .C(n_719), .Y(n_709) );
AND2x4_ASAP7_75t_L g576 ( .A(n_561), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g580 ( .A(n_561), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_561), .B(n_594), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_561), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g693 ( .A(n_561), .B(n_680), .Y(n_693) );
AND2x2_ASAP7_75t_L g579 ( .A(n_563), .B(n_580), .Y(n_579) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_564), .Y(n_597) );
OR2x2_ASAP7_75t_L g686 ( .A(n_564), .B(n_650), .Y(n_686) );
INVx1_ASAP7_75t_L g742 ( .A(n_564), .Y(n_742) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g651 ( .A(n_568), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g665 ( .A(n_568), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g740 ( .A(n_568), .B(n_613), .Y(n_740) );
BUFx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g583 ( .A(n_569), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g602 ( .A(n_569), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g664 ( .A(n_570), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_570), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_719) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g613 ( .A(n_571), .B(n_584), .Y(n_613) );
AND2x4_ASAP7_75t_L g666 ( .A(n_571), .B(n_573), .Y(n_666) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI21xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_579), .B(n_581), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_575), .A2(n_661), .B1(n_665), .B2(n_667), .Y(n_660) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_576), .B(n_594), .Y(n_620) );
INVx2_ASAP7_75t_L g682 ( .A(n_576), .Y(n_682) );
AND2x2_ASAP7_75t_L g696 ( .A(n_576), .B(n_692), .Y(n_696) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g592 ( .A(n_578), .Y(n_592) );
INVx1_ASAP7_75t_L g645 ( .A(n_578), .Y(n_645) );
INVx1_ASAP7_75t_L g596 ( .A(n_580), .Y(n_596) );
AND3x2_ASAP7_75t_L g624 ( .A(n_580), .B(n_625), .C(n_626), .Y(n_624) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g688 ( .A(n_583), .Y(n_688) );
AND2x2_ASAP7_75t_L g616 ( .A(n_585), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g687 ( .A(n_585), .B(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_585), .A2(n_699), .B1(n_703), .B2(n_706), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_585), .B(n_733), .Y(n_737) );
BUFx2_ASAP7_75t_L g628 ( .A(n_586), .Y(n_628) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g599 ( .A(n_587), .Y(n_599) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_587), .Y(n_718) );
OAI221xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_598), .B1(n_600), .B2(n_601), .C(n_604), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_595), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g680 ( .A(n_592), .Y(n_680) );
INVx2_ASAP7_75t_SL g669 ( .A(n_593), .Y(n_669) );
AND2x2_ASAP7_75t_L g751 ( .A(n_593), .B(n_618), .Y(n_751) );
INVx4_ASAP7_75t_L g642 ( .A(n_594), .Y(n_642) );
INVx1_ASAP7_75t_L g600 ( .A(n_595), .Y(n_600) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x4_ASAP7_75t_L g711 ( .A(n_599), .B(n_666), .Y(n_711) );
INVx1_ASAP7_75t_SL g750 ( .A(n_599), .Y(n_750) );
AND2x2_ASAP7_75t_L g755 ( .A(n_599), .B(n_658), .Y(n_755) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g697 ( .A(n_603), .Y(n_697) );
OAI21xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g630 ( .A(n_611), .Y(n_630) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g627 ( .A(n_613), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g717 ( .A(n_613), .B(n_718), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_619), .B(n_621), .C(n_638), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g710 ( .A(n_617), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_618), .B(n_633), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_618), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g743 ( .A(n_618), .B(n_666), .Y(n_743) );
OAI221xp5_ASAP7_75t_SL g654 ( .A1(n_619), .A2(n_643), .B1(n_655), .B2(n_656), .C(n_660), .Y(n_654) );
INVx3_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g725 ( .A(n_620), .B(n_626), .Y(n_725) );
OAI32xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_627), .A3(n_629), .B1(n_631), .B2(n_635), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVxp67_ASAP7_75t_SL g715 ( .A(n_625), .Y(n_715) );
INVx2_ASAP7_75t_L g648 ( .A(n_626), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_L g757 ( .A1(n_626), .A2(n_678), .B(n_758), .C(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g663 ( .A(n_628), .Y(n_663) );
OR2x2_ASAP7_75t_L g759 ( .A(n_628), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_632), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g720 ( .A(n_635), .Y(n_720) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g701 ( .A(n_636), .Y(n_701) );
OAI21xp33_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_647), .B(n_651), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
OR2x2_ASAP7_75t_L g678 ( .A(n_641), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_642), .B(n_645), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_644), .A2(n_676), .B1(n_745), .B2(n_748), .C(n_752), .Y(n_744) );
INVx2_ASAP7_75t_L g747 ( .A(n_644), .Y(n_747) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
OR2x2_ASAP7_75t_L g668 ( .A(n_648), .B(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g735 ( .A(n_648), .B(n_693), .Y(n_735) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g733 ( .A(n_658), .Y(n_733) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_666), .B(n_696), .Y(n_753) );
INVx2_ASAP7_75t_L g760 ( .A(n_666), .Y(n_760) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g730 ( .A1(n_668), .A2(n_731), .B1(n_734), .B2(n_736), .C(n_738), .Y(n_730) );
AND5x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_709), .C(n_724), .D(n_744), .E(n_754), .Y(n_670) );
NOR2xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_689), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_678), .B1(n_681), .B2(n_683), .C(n_684), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI221xp5_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_694), .B1(n_695), .B2(n_697), .C(n_698), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_694), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OR2x2_ASAP7_75t_L g707 ( .A(n_702), .B(n_708), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_716), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_730), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_741), .B2(n_743), .Y(n_738) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_740), .A2(n_755), .B(n_756), .C(n_757), .Y(n_754) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g758 ( .A(n_751), .Y(n_758) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
CKINVDCx11_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_762), .Y(n_770) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx3_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
BUFx4f_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_780), .Y(n_773) );
INVxp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_776), .B(n_779), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_SL g797 ( .A(n_777), .B(n_779), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_777), .A2(n_800), .B(n_803), .Y(n_799) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
BUFx3_ASAP7_75t_L g788 ( .A(n_781), .Y(n_788) );
BUFx2_ASAP7_75t_L g804 ( .A(n_781), .Y(n_804) );
INVxp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_787), .B(n_789), .Y(n_783) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_788), .Y(n_792) );
NOR2xp33_ASAP7_75t_SL g789 ( .A(n_790), .B(n_793), .Y(n_789) );
INVx1_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
CKINVDCx11_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
CKINVDCx8_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
endmodule