module fake_jpeg_2961_n_212 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_212);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_33),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_83),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_1),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_58),
.B1(n_65),
.B2(n_70),
.Y(n_93)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_SL g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx2_ASAP7_75t_SL g107 ( 
.A(n_98),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_54),
.B(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_66),
.B1(n_65),
.B2(n_70),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_69),
.B1(n_64),
.B2(n_74),
.Y(n_109)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_63),
.C(n_55),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_120),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_80),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_5),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_118),
.B(n_98),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_71),
.B(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_54),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_57),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_61),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_137),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_143),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_75),
.B1(n_76),
.B2(n_67),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_125),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_76),
.B1(n_99),
.B2(n_91),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_76),
.B(n_20),
.C(n_25),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_17),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_10),
.C(n_12),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_2),
.CI(n_4),
.CON(n_139),
.SN(n_139)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_6),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_31),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_39),
.B(n_50),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_4),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_152),
.C(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_155),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_154),
.A2(n_46),
.B1(n_51),
.B2(n_146),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_162),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_37),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_163),
.C(n_35),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_9),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_40),
.C(n_48),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_15),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_15),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_16),
.B(n_30),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_175),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_152),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_36),
.B(n_41),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_176),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_184),
.B1(n_160),
.B2(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_147),
.B1(n_145),
.B2(n_167),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_145),
.B(n_165),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_171),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_181),
.B1(n_174),
.B2(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_170),
.B1(n_185),
.B2(n_177),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_172),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_189),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_198),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_199),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_189),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_205),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_205),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_208),
.B(n_206),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_202),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_197),
.Y(n_212)
);


endmodule