module fake_jpeg_9863_n_303 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_286;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_273;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_300;
wire n_211;
wire n_294;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_44),
.B(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_34),
.B1(n_30),
.B2(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_33),
.B1(n_20),
.B2(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_63),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_30),
.B1(n_26),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_72),
.B1(n_78),
.B2(n_83),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_85),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_87),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_61),
.B(n_57),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_90),
.B(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_20),
.B1(n_23),
.B2(n_19),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_15),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_20),
.B1(n_23),
.B2(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_84),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_19),
.B1(n_33),
.B2(n_23),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_92),
.B1(n_94),
.B2(n_60),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_20),
.B1(n_19),
.B2(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_27),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_63),
.B1(n_48),
.B2(n_18),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_21),
.B(n_22),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_102),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_60),
.A3(n_41),
.B1(n_54),
.B2(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_108),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_120),
.B1(n_86),
.B2(n_84),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_21),
.B(n_54),
.Y(n_143)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_115),
.Y(n_142)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_41),
.A3(n_54),
.B1(n_64),
.B2(n_53),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_118),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_71),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_27),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_22),
.B1(n_27),
.B2(n_18),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_0),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_21),
.B(n_18),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_82),
.C(n_81),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_21),
.C(n_2),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_82),
.B1(n_81),
.B2(n_40),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_126),
.B1(n_133),
.B2(n_135),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_129),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_40),
.B1(n_75),
.B2(n_76),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_75),
.B1(n_76),
.B2(n_66),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_140),
.B1(n_143),
.B2(n_107),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_18),
.B1(n_27),
.B2(n_79),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_141),
.B(n_1),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_139),
.B(n_3),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_64),
.B(n_54),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_21),
.B1(n_62),
.B2(n_64),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_151),
.B1(n_117),
.B2(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_21),
.B1(n_71),
.B2(n_2),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_158),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_112),
.B(n_103),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_156),
.A2(n_171),
.B(n_176),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_161),
.B1(n_169),
.B2(n_128),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_162),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_96),
.B1(n_113),
.B2(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_71),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_107),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_145),
.B1(n_147),
.B2(n_143),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_128),
.B1(n_138),
.B2(n_143),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_0),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_141),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_4),
.C(n_7),
.Y(n_202)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_3),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_181),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_134),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_189),
.B1(n_200),
.B2(n_178),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_156),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_201),
.C(n_202),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_137),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_153),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_4),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_8),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_174),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_10),
.C(n_11),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_202),
.C(n_204),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_152),
.B(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_203),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_214),
.Y(n_238)
);

OA21x2_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_173),
.B(n_171),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_213),
.B(n_192),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_163),
.B1(n_162),
.B2(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_209),
.B1(n_205),
.B2(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_158),
.Y(n_221)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_175),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_231),
.Y(n_245)
);

OAI221xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_160),
.B1(n_171),
.B2(n_176),
.C(n_157),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_177),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_197),
.B1(n_186),
.B2(n_200),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_233),
.B1(n_187),
.B2(n_197),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_154),
.C(n_12),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_205),
.B1(n_199),
.B2(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_249),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_214),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_186),
.B1(n_154),
.B2(n_199),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_248),
.A2(n_236),
.B(n_246),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_194),
.B1(n_192),
.B2(n_208),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_239),
.B(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_265),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_211),
.C(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_257),
.C(n_258),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_211),
.C(n_228),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_239),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_235),
.A2(n_232),
.B1(n_225),
.B2(n_219),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_221),
.C(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_245),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_244),
.B(n_234),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_217),
.CI(n_218),
.CON(n_265),
.SN(n_265)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_272),
.C(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_271),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_260),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_245),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_275),
.B(n_254),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_243),
.B(n_233),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_240),
.Y(n_276)
);

XNOR2x2_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_285),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_14),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_253),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_284),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_256),
.B(n_265),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_12),
.B(n_14),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_276),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_291),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_277),
.A3(n_272),
.B1(n_274),
.B2(n_15),
.C1(n_16),
.C2(n_14),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_278),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_16),
.C(n_290),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_16),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_299),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_294),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_296),
.B(n_290),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_298),
.Y(n_303)
);


endmodule