module fake_jpeg_24713_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_41),
.Y(n_47)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_15),
.B1(n_26),
.B2(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_24),
.B1(n_21),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_26),
.B1(n_15),
.B2(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_24),
.B1(n_28),
.B2(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_15),
.B1(n_24),
.B2(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_60),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_58),
.B1(n_79),
.B2(n_17),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_72),
.Y(n_107)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_63),
.A2(n_70),
.B1(n_74),
.B2(n_84),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_41),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_37),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_22),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_86),
.B(n_39),
.Y(n_103)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_96),
.B1(n_36),
.B2(n_74),
.Y(n_120)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_37),
.B1(n_41),
.B2(n_40),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_97),
.B1(n_79),
.B2(n_36),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_37),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_108),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_39),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_114),
.B1(n_128),
.B2(n_123),
.Y(n_148)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_127),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_86),
.B1(n_63),
.B2(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_69),
.C(n_40),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_33),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_90),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_104),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_110),
.C(n_2),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_121),
.A2(n_101),
.B1(n_105),
.B2(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_148),
.B1(n_149),
.B2(n_38),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_101),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_151),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_111),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_38),
.B1(n_39),
.B2(n_33),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_33),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_38),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_18),
.B(n_25),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_25),
.B(n_20),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_SL g162 ( 
.A(n_136),
.B(n_131),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_166),
.B1(n_170),
.B2(n_173),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_113),
.C(n_118),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_172),
.C(n_147),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_25),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_20),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_175),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_61),
.B(n_56),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_177),
.B1(n_139),
.B2(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_150),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_23),
.B(n_18),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_145),
.B1(n_138),
.B2(n_144),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_185),
.B1(n_173),
.B2(n_156),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_140),
.C(n_153),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_145),
.B1(n_154),
.B2(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_186),
.B(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_141),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_169),
.C(n_163),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_201),
.C(n_189),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_202),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_169),
.C(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_190),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_185),
.C(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_179),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_210),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_187),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_60),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_191),
.B1(n_196),
.B2(n_199),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_209),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_192),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_216),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_9),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_14),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_217),
.B(n_10),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_12),
.B1(n_10),
.B2(n_3),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_213),
.B1(n_212),
.B2(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_223),
.C(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_220),
.C(n_219),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_1),
.C(n_5),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_230),
.A2(n_231),
.A3(n_1),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_22),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_228),
.A2(n_225),
.B1(n_2),
.B2(n_5),
.Y(n_231)
);

AOI321xp33_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_233),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_29),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_29),
.C(n_22),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_29),
.Y(n_236)
);


endmodule