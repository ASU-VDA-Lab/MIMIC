module fake_jpeg_30460_n_422 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_422);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_422;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_3),
.B(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_21),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_71),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_74),
.Y(n_97)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_12),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_84),
.Y(n_107)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

AND2x4_ASAP7_75t_SL g81 ( 
.A(n_27),
.B(n_30),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_27),
.Y(n_121)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_83),
.Y(n_129)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_10),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_49),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_87),
.Y(n_117)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_89),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_38),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_23),
.B1(n_45),
.B2(n_40),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_102),
.B1(n_125),
.B2(n_31),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_33),
.B1(n_38),
.B2(n_45),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_104),
.B1(n_27),
.B2(n_31),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_23),
.B1(n_45),
.B2(n_40),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_38),
.B1(n_23),
.B2(n_30),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_30),
.B1(n_44),
.B2(n_41),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_115),
.B(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_41),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_131),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_40),
.B1(n_28),
.B2(n_46),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_111),
.A2(n_136),
.B1(n_31),
.B2(n_53),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_44),
.B1(n_28),
.B2(n_46),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_134),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_51),
.A2(n_40),
.B1(n_32),
.B2(n_49),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_88),
.B(n_73),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_46),
.B1(n_39),
.B2(n_36),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx5_ASAP7_75t_SL g193 ( 
.A(n_139),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_140),
.A2(n_145),
.B(n_93),
.C(n_125),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_97),
.A2(n_89),
.B1(n_82),
.B2(n_64),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_162),
.B1(n_170),
.B2(n_108),
.Y(n_174)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_66),
.B1(n_24),
.B2(n_36),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_155),
.B1(n_160),
.B2(n_166),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_149),
.B1(n_106),
.B2(n_134),
.Y(n_176)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_67),
.B1(n_69),
.B2(n_68),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_103),
.A2(n_24),
.B1(n_39),
.B2(n_32),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_83),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_134),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_99),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_103),
.A2(n_53),
.B1(n_15),
.B2(n_21),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_101),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_168),
.Y(n_192)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_83),
.B1(n_14),
.B2(n_15),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_117),
.B1(n_92),
.B2(n_112),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_120),
.B(n_107),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_118),
.C(n_151),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_188),
.B1(n_152),
.B2(n_170),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_160),
.B1(n_149),
.B2(n_147),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_95),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_157),
.C(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_126),
.C(n_119),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_141),
.A2(n_101),
.B1(n_129),
.B2(n_108),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_138),
.B(n_142),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_139),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_191),
.B1(n_133),
.B2(n_108),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_209),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_150),
.C(n_169),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_214),
.C(n_215),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_165),
.CI(n_158),
.CON(n_205),
.SN(n_205)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_220),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_154),
.B(n_118),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_195),
.B(n_182),
.Y(n_231)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_211),
.B1(n_218),
.B2(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_178),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_148),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_183),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_126),
.C(n_119),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_144),
.C(n_168),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_133),
.B1(n_130),
.B2(n_114),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_130),
.B1(n_128),
.B2(n_98),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_191),
.B(n_21),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_192),
.C(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_203),
.C(n_207),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_226),
.Y(n_262)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_236),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_195),
.B(n_182),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_235),
.B(n_237),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_195),
.B(n_198),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_193),
.B1(n_173),
.B2(n_152),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_173),
.B(n_189),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_189),
.B(n_205),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_215),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_243),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_206),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_221),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_253),
.C(n_256),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_242),
.A2(n_200),
.B1(n_210),
.B2(n_211),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_263),
.B1(n_221),
.B2(n_224),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_212),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_222),
.B(n_229),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_239),
.C(n_232),
.Y(n_256)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_205),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_229),
.Y(n_274)
);

AOI32xp33_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_205),
.A3(n_220),
.B1(n_204),
.B2(n_212),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_241),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_214),
.B1(n_201),
.B2(n_185),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_183),
.B1(n_190),
.B2(n_185),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_237),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_227),
.A2(n_226),
.B1(n_223),
.B2(n_228),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_190),
.B1(n_193),
.B2(n_197),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_197),
.C(n_164),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_221),
.C(n_224),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_283),
.Y(n_318)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_277),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_285),
.C(n_287),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_238),
.B1(n_223),
.B2(n_222),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_271),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_247),
.B(n_193),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_288),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_291),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_240),
.B1(n_225),
.B2(n_97),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_256),
.C(n_268),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_254),
.A2(n_97),
.B1(n_92),
.B2(n_112),
.Y(n_286)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_260),
.B(n_175),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_189),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_175),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_290),
.C(n_257),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_187),
.C(n_180),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_162),
.B1(n_196),
.B2(n_180),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_96),
.B(n_175),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_309),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_297),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_269),
.Y(n_297)
);

BUFx12_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_263),
.B1(n_252),
.B2(n_255),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_302),
.B1(n_312),
.B2(n_286),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_267),
.B1(n_264),
.B2(n_246),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_258),
.Y(n_305)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_258),
.Y(n_308)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_272),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_266),
.B1(n_257),
.B2(n_196),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_187),
.Y(n_314)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_17),
.Y(n_315)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_272),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_317),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_284),
.B1(n_281),
.B2(n_283),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_319),
.A2(n_329),
.B1(n_334),
.B2(n_340),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_306),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_SL g351 ( 
.A(n_322),
.B(n_306),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_309),
.C(n_307),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_335),
.C(n_302),
.Y(n_354)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_128),
.B1(n_98),
.B2(n_135),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_330),
.B(n_297),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_329),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_303),
.A2(n_135),
.B(n_152),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_304),
.B(n_316),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_295),
.A2(n_10),
.B1(n_20),
.B2(n_19),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_124),
.C(n_94),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_124),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_312),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_20),
.Y(n_338)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_338),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_308),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_307),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_345),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_318),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_347),
.Y(n_373)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_350),
.C(n_352),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_316),
.B1(n_311),
.B2(n_301),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_352),
.A2(n_323),
.B1(n_340),
.B2(n_339),
.Y(n_367)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_338),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_353),
.B(n_354),
.Y(n_372)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_355),
.A2(n_356),
.B1(n_358),
.B2(n_349),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_326),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_341),
.B(n_304),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_357),
.A2(n_334),
.B(n_333),
.Y(n_368)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_359),
.A2(n_331),
.B(n_321),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_324),
.C(n_328),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_362),
.C(n_363),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_358),
.B(n_349),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_328),
.C(n_322),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_327),
.C(n_336),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_367),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_351),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_369),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_335),
.C(n_298),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_298),
.C(n_124),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_342),
.B1(n_359),
.B2(n_344),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_376),
.A2(n_379),
.B1(n_364),
.B2(n_2),
.Y(n_391)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_377),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_381),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_372),
.A2(n_373),
.B1(n_370),
.B2(n_366),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_360),
.A2(n_298),
.B(n_343),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_380),
.A2(n_379),
.B(n_375),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_383),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_16),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_16),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_384),
.B(n_0),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_361),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_373),
.B1(n_2),
.B2(n_3),
.Y(n_386)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_364),
.C(n_2),
.Y(n_389)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_389),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_385),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_SL g394 ( 
.A(n_377),
.B(n_376),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_394),
.B(n_381),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_375),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_5),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_0),
.B(n_5),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_396),
.B(n_5),
.Y(n_403)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_397),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_399),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_403),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_29),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_404),
.A2(n_392),
.B(n_387),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_406),
.A2(n_410),
.B1(n_405),
.B2(n_398),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_394),
.C(n_389),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_407),
.A2(n_402),
.B(n_397),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_400),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_412),
.A2(n_413),
.B(n_414),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_6),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_6),
.Y(n_415)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g416 ( 
.A1(n_415),
.A2(n_408),
.B(n_9),
.C(n_8),
.D(n_29),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_416),
.B(n_8),
.C(n_9),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_418),
.A2(n_417),
.B(n_9),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_8),
.C(n_9),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_29),
.C(n_398),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_29),
.Y(n_422)
);


endmodule