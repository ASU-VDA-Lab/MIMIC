module fake_jpeg_17961_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_28),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_31),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_32),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_38),
.C(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_15),
.Y(n_74)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_72),
.Y(n_80)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_77),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_45),
.B1(n_56),
.B2(n_16),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_40),
.A3(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_74),
.Y(n_94)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_36),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_20),
.C(n_19),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_R g95 ( 
.A(n_76),
.B(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_57),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_37),
.B1(n_32),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_45),
.B1(n_41),
.B2(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_50),
.C(n_48),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_56),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_95),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_101),
.B1(n_45),
.B2(n_70),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_97),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_37),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_74),
.B(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_73),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_65),
.B1(n_78),
.B2(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_37),
.B1(n_52),
.B2(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_119),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_106),
.B1(n_117),
.B2(n_121),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_65),
.B1(n_75),
.B2(n_70),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_74),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_46),
.B(n_75),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_116),
.B(n_86),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_82),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_84),
.B1(n_98),
.B2(n_42),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_94),
.B(n_83),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_42),
.B1(n_73),
.B2(n_36),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_84),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_52),
.B1(n_34),
.B2(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_93),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_130),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_52),
.B1(n_63),
.B2(n_96),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_137),
.B1(n_111),
.B2(n_30),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_138),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_89),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_133),
.B(n_136),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_113),
.C(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_89),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_140),
.B1(n_105),
.B2(n_120),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_94),
.B(n_99),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_101),
.B1(n_97),
.B2(n_85),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_15),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_142),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_116),
.C(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_104),
.B1(n_115),
.B2(n_109),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_145),
.B1(n_150),
.B2(n_138),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_22),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_152),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_46),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_154),
.B(n_133),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_46),
.C(n_22),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_15),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_30),
.Y(n_169)
);

AOI21x1_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_30),
.B(n_24),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_160),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_139),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_126),
.B1(n_124),
.B2(n_130),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_137),
.C(n_122),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_124),
.B1(n_127),
.B2(n_131),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_146),
.C(n_153),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_149),
.B1(n_156),
.B2(n_148),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_171),
.B1(n_161),
.B2(n_165),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_164),
.A2(n_155),
.B1(n_142),
.B2(n_149),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_173),
.C(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_24),
.C(n_14),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_24),
.C(n_14),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_4),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_8),
.B(n_9),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_169),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_159),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_165),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_167),
.C(n_8),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_187),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_4),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_175),
.B1(n_178),
.B2(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_171),
.B1(n_170),
.B2(n_10),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_9),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_183),
.B1(n_185),
.B2(n_12),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_191),
.C(n_193),
.Y(n_198)
);

AOI211xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_197),
.B(n_191),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_199),
.B(n_194),
.Y(n_202)
);

OAI21x1_ASAP7_75t_SL g201 ( 
.A1(n_200),
.A2(n_195),
.B(n_13),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_202),
.B(n_12),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_13),
.Y(n_204)
);


endmodule