module fake_jpeg_10302_n_128 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_1),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_1),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_2),
.B(n_3),
.Y(n_77)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_59),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_2),
.B1(n_44),
.B2(n_7),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_11),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_92),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_49),
.B1(n_54),
.B2(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_91),
.B1(n_6),
.B2(n_10),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_60),
.B1(n_65),
.B2(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_64),
.B1(n_53),
.B2(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_52),
.C(n_3),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_12),
.C(n_15),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_105)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_109),
.B1(n_103),
.B2(n_100),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_106),
.B(n_107),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_104),
.C(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_102),
.B1(n_105),
.B2(n_101),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_95),
.B1(n_79),
.B2(n_78),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_19),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_20),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_21),
.B(n_22),
.Y(n_122)
);

AO21x1_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_28),
.B(n_30),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_32),
.B(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_34),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_37),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_39),
.B(n_40),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_41),
.Y(n_128)
);


endmodule