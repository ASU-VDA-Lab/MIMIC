module fake_jpeg_14506_n_87 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_87);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_87;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_1),
.B(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_9),
.C(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_35),
.B1(n_36),
.B2(n_30),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_44)
);

FAx1_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_4),
.CI(n_5),
.CON(n_61),
.SN(n_61)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_47),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_10),
.C(n_19),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_59),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_8),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_11),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_46),
.B1(n_45),
.B2(n_48),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_6),
.C(n_7),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_15),
.B(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_48),
.B1(n_16),
.B2(n_17),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_74),
.C(n_61),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_79),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_72),
.C(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_80),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_78),
.B(n_72),
.C(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_75),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_86),
.B(n_27),
.Y(n_87)
);


endmodule