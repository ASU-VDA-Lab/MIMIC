module fake_jpeg_6047_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_8),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_15),
.B1(n_12),
.B2(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_12),
.B1(n_15),
.B2(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_12),
.B1(n_16),
.B2(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_13),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_13),
.B1(n_10),
.B2(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_32),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_18),
.B1(n_17),
.B2(n_23),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_23),
.B1(n_31),
.B2(n_35),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_30),
.B1(n_7),
.B2(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_41),
.B1(n_37),
.B2(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_41),
.B1(n_39),
.B2(n_13),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_24),
.C(n_17),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_24),
.C(n_10),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_62),
.C(n_52),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_44),
.B1(n_49),
.B2(n_46),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_61),
.B(n_55),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_10),
.B(n_2),
.C(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_67),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.C(n_59),
.Y(n_70)
);

OAI321xp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_57),
.A3(n_10),
.B1(n_6),
.B2(n_24),
.C(n_3),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_61),
.B1(n_59),
.B2(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_1),
.B(n_2),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_4),
.Y(n_77)
);


endmodule