module fake_ariane_2772_n_1214 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1214);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1214;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1209;
wire n_1137;
wire n_646;
wire n_1174;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_1029;
wire n_341;
wire n_1187;
wire n_985;
wire n_421;
wire n_245;
wire n_1167;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_1180;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_244;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_1095;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_1200;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_756;
wire n_466;
wire n_940;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_1181;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_162;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_1208;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_1133;
wire n_900;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_899;
wire n_500;
wire n_754;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_903;
wire n_871;
wire n_315;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_167;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_158;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_1201;
wire n_1107;
wire n_173;
wire n_989;
wire n_242;
wire n_645;
wire n_858;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_795;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_770;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_1153;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_222;
wire n_478;
wire n_703;
wire n_1207;
wire n_748;
wire n_1212;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_1074;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_1080;
wire n_576;
wire n_843;
wire n_1148;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_163;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_977;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_1136;
wire n_221;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_1213;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_260;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_1089;
wire n_565;
wire n_236;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_1194;
wire n_907;
wire n_225;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_1210;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_199;
wire n_1135;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1041;
wire n_571;
wire n_680;
wire n_414;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_249;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_171;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_161;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_692;
wire n_216;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_195;
wire n_606;
wire n_1026;
wire n_951;
wire n_938;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_626;
wire n_430;
wire n_493;
wire n_722;
wire n_1206;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_998;
wire n_999;
wire n_1083;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_1211;
wire n_963;
wire n_873;
wire n_1139;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_159;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_434;
wire n_263;
wire n_360;
wire n_1102;
wire n_975;
wire n_1101;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_165;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_470;
wire n_266;
wire n_457;
wire n_1087;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1164;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_1011;
wire n_642;
wire n_978;
wire n_211;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_30),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_112),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_31),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_92),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_84),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_55),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_17),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_97),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_39),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_34),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_14),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_45),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_50),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_43),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_142),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_25),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_154),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_116),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_33),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_4),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_88),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_67),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_39),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_32),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_36),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_26),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_101),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_121),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_13),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_133),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_18),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_48),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_120),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_37),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_33),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_36),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_126),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_130),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_151),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_3),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_77),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_46),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_91),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_110),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_103),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_24),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_107),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_119),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_104),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_137),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_34),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_127),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_144),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_98),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_42),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_35),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_10),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_87),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_53),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_82),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_4),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_83),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_89),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_113),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_63),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_95),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_10),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_60),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_16),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_38),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_139),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_147),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_41),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_122),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_111),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_54),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_134),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_72),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_22),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_156),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_146),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_27),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_68),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_114),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_81),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_125),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_170),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_190),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_161),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_190),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_186),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_179),
.B(n_0),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_158),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_243),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_179),
.Y(n_292)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_172),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_172),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_158),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_206),
.B(n_0),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_174),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_240),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_174),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_187),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_246),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_1),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_187),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_159),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_160),
.B(n_1),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_205),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_193),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_188),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_195),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_193),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_197),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_201),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_208),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_208),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_232),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_232),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_202),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_207),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_238),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_238),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_226),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_246),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_273),
.B(n_2),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_242),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_242),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_255),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_251),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_273),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_189),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_255),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_251),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_176),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_272),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_222),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_189),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_181),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_212),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_161),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_176),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_166),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_222),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_272),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_183),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_184),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_178),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_168),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_203),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_209),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_198),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_258),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_278),
.B(n_2),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_230),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_239),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_254),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_258),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_168),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_257),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_L g370 ( 
.A(n_306),
.B(n_191),
.Y(n_370)
);

OAI21x1_ASAP7_75t_L g371 ( 
.A1(n_305),
.A2(n_277),
.B(n_191),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_173),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_339),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_173),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_285),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_280),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_302),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_335),
.B(n_269),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_292),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_336),
.B(n_269),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_248),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_290),
.B(n_162),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_354),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_292),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_303),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_345),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_279),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_347),
.A2(n_183),
.B1(n_175),
.B2(n_194),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_362),
.B(n_248),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_342),
.B(n_204),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_296),
.B(n_276),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_300),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_364),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_351),
.B(n_248),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_311),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_312),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_282),
.B(n_248),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_314),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_315),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_321),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_353),
.A2(n_289),
.B1(n_297),
.B2(n_295),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_284),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_288),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_325),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_287),
.B(n_307),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_281),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

AND2x2_ASAP7_75t_SL g427 ( 
.A(n_361),
.B(n_248),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_283),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_308),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_344),
.B(n_163),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_309),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_333),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_294),
.B(n_253),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_352),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_424),
.B(n_334),
.Y(n_445)
);

BUFx4f_ASAP7_75t_L g446 ( 
.A(n_427),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_396),
.B(n_356),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_372),
.B(n_318),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

OR2x6_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_326),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_356),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_398),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_373),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_372),
.B(n_349),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_366),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_290),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_399),
.B(n_410),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_399),
.B(n_366),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_372),
.B(n_350),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_427),
.B(n_280),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_427),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_437),
.B(n_286),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_391),
.A2(n_293),
.B1(n_298),
.B2(n_217),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_410),
.B(n_298),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_391),
.A2(n_293),
.B1(n_214),
.B2(n_219),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_394),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_375),
.B(n_355),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_359),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_405),
.A2(n_340),
.B1(n_299),
.B2(n_328),
.Y(n_479)
);

BUFx6f_ASAP7_75t_SL g480 ( 
.A(n_433),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_377),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_391),
.B(n_286),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_413),
.A2(n_241),
.B1(n_224),
.B2(n_245),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_415),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_384),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_375),
.B(n_291),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_291),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_412),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_398),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_395),
.B(n_165),
.C(n_164),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_384),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

AO21x2_ASAP7_75t_L g496 ( 
.A1(n_371),
.A2(n_263),
.B(n_253),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_384),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_386),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_392),
.B(n_299),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_386),
.Y(n_503)
);

AO21x2_ASAP7_75t_L g504 ( 
.A1(n_371),
.A2(n_263),
.B(n_253),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_431),
.B(n_233),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_392),
.B(n_301),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_380),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_379),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_446),
.B(n_437),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_446),
.B(n_437),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_429),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_375),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_461),
.B(n_437),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_446),
.B(n_437),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

NOR3xp33_ASAP7_75t_L g518 ( 
.A(n_459),
.B(n_378),
.C(n_380),
.Y(n_518)
);

O2A1O1Ixp5_ASAP7_75t_L g519 ( 
.A1(n_461),
.A2(n_406),
.B(n_435),
.C(n_434),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_459),
.B(n_378),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_397),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_447),
.B(n_437),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_397),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_446),
.B(n_437),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_466),
.A2(n_405),
.B1(n_406),
.B2(n_401),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_452),
.B(n_397),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_509),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_L g530 ( 
.A1(n_452),
.A2(n_463),
.B(n_458),
.C(n_443),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_458),
.B(n_385),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_440),
.B(n_437),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_463),
.B(n_433),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_442),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_508),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_443),
.B(n_385),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_L g539 ( 
.A(n_466),
.B(n_438),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_480),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_491),
.B(n_434),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_465),
.B(n_438),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_450),
.B(n_435),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_480),
.Y(n_544)
);

AO221x1_ASAP7_75t_L g545 ( 
.A1(n_479),
.A2(n_400),
.B1(n_378),
.B2(n_418),
.C(n_438),
.Y(n_545)
);

AND2x6_ASAP7_75t_SL g546 ( 
.A(n_488),
.B(n_422),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_510),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_490),
.B(n_429),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_440),
.B(n_438),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_462),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_454),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_L g553 ( 
.A(n_501),
.B(n_507),
.C(n_488),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_445),
.B(n_418),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_462),
.Y(n_555)
);

O2A1O1Ixp33_ASAP7_75t_L g556 ( 
.A1(n_476),
.A2(n_412),
.B(n_395),
.C(n_408),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_491),
.B(n_435),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_448),
.B(n_439),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

NOR2xp67_ASAP7_75t_SL g560 ( 
.A(n_510),
.B(n_439),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_477),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_477),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_487),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_450),
.B(n_435),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_466),
.B(n_401),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_471),
.B(n_401),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_471),
.B(n_401),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_487),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_494),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_494),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_457),
.B(n_438),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_480),
.Y(n_572)
);

INVx8_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_497),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_457),
.B(n_438),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_457),
.B(n_438),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_440),
.B(n_468),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_497),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_469),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_476),
.B(n_448),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_448),
.B(n_438),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_465),
.B(n_388),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_509),
.B(n_412),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_488),
.B(n_304),
.C(n_301),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_484),
.B(n_411),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_469),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_498),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_498),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_490),
.B(n_483),
.Y(n_589)
);

NOR3xp33_ASAP7_75t_L g590 ( 
.A(n_479),
.B(n_483),
.C(n_484),
.Y(n_590)
);

CKINVDCx11_ASAP7_75t_R g591 ( 
.A(n_450),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_440),
.B(n_415),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_445),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_445),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_489),
.B(n_388),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_450),
.A2(n_370),
.B1(n_436),
.B2(n_408),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_509),
.B(n_468),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_493),
.B(n_411),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_499),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_440),
.B(n_415),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_464),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_468),
.B(n_415),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_489),
.B(n_450),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_450),
.B(n_412),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_472),
.A2(n_475),
.B1(n_464),
.B2(n_485),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_464),
.A2(n_370),
.B1(n_436),
.B2(n_408),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_412),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_475),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_534),
.B(n_472),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_520),
.B(n_304),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_534),
.B(n_470),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

OAI21xp33_ASAP7_75t_L g613 ( 
.A1(n_514),
.A2(n_470),
.B(n_485),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_524),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_537),
.A2(n_467),
.B(n_486),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_597),
.A2(n_467),
.B(n_486),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_608),
.A2(n_319),
.B1(n_320),
.B2(n_310),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_559),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_521),
.A2(n_486),
.B(n_453),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_561),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_563),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_523),
.A2(n_486),
.B(n_453),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_525),
.A2(n_486),
.B(n_453),
.Y(n_623)
);

NOR2x2_ASAP7_75t_L g624 ( 
.A(n_554),
.B(n_313),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_528),
.A2(n_460),
.B(n_444),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_532),
.B(n_310),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_595),
.B(n_530),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_541),
.A2(n_460),
.B(n_444),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_557),
.A2(n_460),
.B(n_444),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_535),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_548),
.B(n_319),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_595),
.B(n_455),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_SL g633 ( 
.A(n_605),
.B(n_323),
.C(n_320),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_R g634 ( 
.A(n_536),
.B(n_323),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_511),
.A2(n_478),
.B(n_474),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_511),
.A2(n_478),
.B(n_474),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_517),
.B(n_324),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_512),
.A2(n_478),
.B(n_474),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_580),
.B(n_393),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_512),
.A2(n_482),
.B(n_481),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_519),
.A2(n_371),
.B(n_499),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_516),
.A2(n_482),
.B(n_481),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_516),
.A2(n_482),
.B(n_481),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_526),
.A2(n_500),
.B(n_495),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_585),
.B(n_393),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_601),
.B(n_393),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_526),
.A2(n_500),
.B(n_495),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_515),
.A2(n_500),
.B(n_495),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_607),
.B(n_420),
.Y(n_649)
);

NOR2x1_ASAP7_75t_L g650 ( 
.A(n_513),
.B(n_493),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_568),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_531),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_582),
.A2(n_503),
.B(n_449),
.C(n_441),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_579),
.B(n_324),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_573),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_590),
.A2(n_553),
.B1(n_518),
.B2(n_603),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_566),
.A2(n_505),
.B(n_449),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_543),
.A2(n_564),
.B1(n_582),
.B2(n_593),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_567),
.A2(n_505),
.B(n_449),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g660 ( 
.A(n_552),
.B(n_328),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_571),
.B(n_420),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_575),
.A2(n_503),
.B(n_422),
.C(n_425),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_589),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_588),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_539),
.A2(n_505),
.B(n_449),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_586),
.B(n_340),
.Y(n_666)
);

AO21x1_ASAP7_75t_L g667 ( 
.A1(n_542),
.A2(n_376),
.B(n_374),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_543),
.B(n_564),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_420),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_602),
.A2(n_451),
.B(n_441),
.Y(n_670)
);

BUFx4f_ASAP7_75t_L g671 ( 
.A(n_573),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_535),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_594),
.B(n_316),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_542),
.A2(n_441),
.B(n_502),
.C(n_473),
.Y(n_674)
);

AO21x1_ASAP7_75t_L g675 ( 
.A1(n_577),
.A2(n_376),
.B(n_374),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_558),
.B(n_317),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_538),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_602),
.A2(n_451),
.B(n_441),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_581),
.B(n_420),
.Y(n_679)
);

OAI321xp33_ASAP7_75t_L g680 ( 
.A1(n_606),
.A2(n_400),
.A3(n_421),
.B1(n_425),
.B2(n_402),
.C(n_382),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_604),
.A2(n_473),
.B(n_451),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_538),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_546),
.B(n_329),
.Y(n_683)
);

O2A1O1Ixp33_ASAP7_75t_SL g684 ( 
.A1(n_522),
.A2(n_473),
.B(n_451),
.C(n_502),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_583),
.A2(n_502),
.B(n_473),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_560),
.B(n_527),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_549),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_591),
.B(n_502),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_584),
.B(n_421),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_543),
.B(n_402),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_564),
.B(n_509),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_549),
.B(n_390),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_551),
.A2(n_379),
.B1(n_409),
.B2(n_428),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_551),
.A2(n_504),
.B(n_496),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_555),
.B(n_390),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_555),
.A2(n_504),
.B(n_496),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_562),
.A2(n_504),
.B(n_496),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_556),
.A2(n_409),
.B(n_390),
.Y(n_699)
);

AND2x6_ASAP7_75t_L g700 ( 
.A(n_559),
.B(n_509),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_562),
.A2(n_504),
.B(n_496),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_554),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_540),
.B(n_509),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_569),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_SL g705 ( 
.A(n_611),
.B(n_265),
.C(n_237),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_620),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_655),
.B(n_573),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_632),
.B(n_540),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_612),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_626),
.B(n_544),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_609),
.B(n_545),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_613),
.A2(n_547),
.B(n_599),
.C(n_569),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_627),
.A2(n_529),
.B(n_533),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_614),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_654),
.B(n_596),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_676),
.B(n_421),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_639),
.B(n_570),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_R g718 ( 
.A(n_671),
.B(n_544),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_656),
.A2(n_598),
.B(n_533),
.C(n_550),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_660),
.B(n_572),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_645),
.B(n_570),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_663),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_619),
.A2(n_529),
.B(n_550),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_653),
.A2(n_578),
.B(n_574),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_673),
.B(n_572),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_637),
.B(n_415),
.C(n_430),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_672),
.B(n_574),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_621),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_617),
.B(n_578),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_658),
.B(n_529),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_615),
.A2(n_599),
.B(n_587),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_655),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_651),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_657),
.A2(n_529),
.B(n_587),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_659),
.A2(n_577),
.B(n_592),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_610),
.B(n_592),
.Y(n_736)
);

AND2x2_ASAP7_75t_SL g737 ( 
.A(n_671),
.B(n_696),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_623),
.A2(n_600),
.B(n_565),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_625),
.A2(n_600),
.B(n_509),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_631),
.B(n_430),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_655),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_700),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_682),
.B(n_379),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_646),
.B(n_423),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_652),
.B(n_634),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_646),
.B(n_423),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_628),
.A2(n_468),
.B(n_409),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_664),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_690),
.B(n_423),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_629),
.A2(n_622),
.B(n_635),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_633),
.B(n_432),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_686),
.B(n_618),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_668),
.B(n_432),
.Y(n_753)
);

CKINVDCx16_ASAP7_75t_R g754 ( 
.A(n_683),
.Y(n_754)
);

BUFx8_ASAP7_75t_L g755 ( 
.A(n_702),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_650),
.A2(n_436),
.B1(n_415),
.B2(n_403),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_704),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_666),
.A2(n_428),
.B(n_426),
.C(n_419),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_689),
.B(n_409),
.Y(n_759)
);

O2A1O1Ixp5_ASAP7_75t_L g760 ( 
.A1(n_667),
.A2(n_382),
.B(n_383),
.C(n_379),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_636),
.A2(n_468),
.B(n_379),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_688),
.B(n_680),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_630),
.B(n_414),
.Y(n_763)
);

BUFx8_ASAP7_75t_L g764 ( 
.A(n_700),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_618),
.B(n_413),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_638),
.A2(n_468),
.B(n_436),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_700),
.Y(n_768)
);

OAI21xp33_ASAP7_75t_SL g769 ( 
.A1(n_681),
.A2(n_383),
.B(n_413),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_750),
.A2(n_734),
.B(n_739),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_713),
.A2(n_616),
.B(n_694),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_754),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_755),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_715),
.B(n_677),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_722),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_735),
.A2(n_675),
.A3(n_701),
.B(n_698),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_736),
.A2(n_705),
.B(n_745),
.C(n_740),
.Y(n_777)
);

INVx3_ASAP7_75t_SL g778 ( 
.A(n_737),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_721),
.A2(n_697),
.B(n_665),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_706),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_716),
.B(n_687),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_709),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_731),
.A2(n_674),
.B(n_648),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_723),
.A2(n_641),
.B(n_640),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_764),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_725),
.B(n_692),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_741),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_731),
.A2(n_684),
.B(n_693),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_755),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_741),
.Y(n_790)
);

NAND3x1_ASAP7_75t_L g791 ( 
.A(n_762),
.B(n_624),
.C(n_389),
.Y(n_791)
);

AOI21x1_ASAP7_75t_L g792 ( 
.A1(n_747),
.A2(n_703),
.B(n_641),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_729),
.B(n_662),
.C(n_699),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_746),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_738),
.A2(n_643),
.B(n_642),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_717),
.A2(n_724),
.B(n_767),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_SL g797 ( 
.A1(n_751),
.A2(n_699),
.B1(n_695),
.B2(n_692),
.Y(n_797)
);

INVx3_ASAP7_75t_SL g798 ( 
.A(n_741),
.Y(n_798)
);

NOR3xp33_ASAP7_75t_L g799 ( 
.A(n_710),
.B(n_416),
.C(n_413),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_719),
.A2(n_695),
.B(n_649),
.C(n_681),
.Y(n_800)
);

AOI21x1_ASAP7_75t_L g801 ( 
.A1(n_752),
.A2(n_761),
.B(n_708),
.Y(n_801)
);

AOI21xp33_ASAP7_75t_L g802 ( 
.A1(n_711),
.A2(n_693),
.B(n_669),
.Y(n_802)
);

AO31x2_ASAP7_75t_L g803 ( 
.A1(n_727),
.A2(n_644),
.A3(n_647),
.B(n_661),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_744),
.A2(n_691),
.B1(n_679),
.B2(n_416),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_724),
.A2(n_678),
.B(n_670),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_749),
.A2(n_416),
.B(n_417),
.C(n_419),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_728),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_732),
.B(n_700),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_764),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_712),
.A2(n_685),
.B(n_468),
.Y(n_810)
);

BUFx8_ASAP7_75t_L g811 ( 
.A(n_707),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_733),
.B(n_416),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_769),
.A2(n_419),
.B(n_417),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_748),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_757),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_760),
.A2(n_759),
.B(n_743),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_742),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_726),
.A2(n_417),
.B1(n_428),
.B2(n_426),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_742),
.B(n_768),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_753),
.B(n_417),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_732),
.B(n_714),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_720),
.B(n_389),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_727),
.B(n_419),
.Y(n_823)
);

O2A1O1Ixp5_ASAP7_75t_L g824 ( 
.A1(n_765),
.A2(n_428),
.B(n_426),
.C(n_386),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_775),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_797),
.A2(n_730),
.B1(n_756),
.B2(n_387),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_817),
.Y(n_827)
);

BUFx2_ASAP7_75t_R g828 ( 
.A(n_778),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_774),
.B(n_743),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_798),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_SL g831 ( 
.A1(n_797),
.A2(n_742),
.B1(n_718),
.B2(n_765),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_780),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_776),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_SL g834 ( 
.A1(n_793),
.A2(n_707),
.B1(n_766),
.B2(n_436),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_811),
.Y(n_835)
);

OAI22xp33_ASAP7_75t_L g836 ( 
.A1(n_786),
.A2(n_763),
.B1(n_407),
.B2(n_387),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_815),
.B(n_386),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_814),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_793),
.A2(n_791),
.B1(n_781),
.B2(n_809),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_782),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_776),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_807),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_817),
.Y(n_843)
);

CKINVDCx6p67_ASAP7_75t_R g844 ( 
.A(n_807),
.Y(n_844)
);

BUFx2_ASAP7_75t_SL g845 ( 
.A(n_809),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_SL g846 ( 
.A1(n_811),
.A2(n_707),
.B1(n_436),
.B2(n_763),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_794),
.A2(n_404),
.B1(n_387),
.B2(n_407),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_772),
.A2(n_707),
.B1(n_426),
.B2(n_403),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_794),
.B(n_389),
.Y(n_849)
);

OAI22xp33_ASAP7_75t_L g850 ( 
.A1(n_773),
.A2(n_387),
.B1(n_404),
.B2(n_407),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_789),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_787),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_802),
.A2(n_404),
.B1(n_407),
.B2(n_415),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_787),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_803),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_821),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_802),
.A2(n_404),
.B1(n_389),
.B2(n_403),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_785),
.A2(n_707),
.B1(n_403),
.B2(n_253),
.Y(n_858)
);

INVx6_ASAP7_75t_L g859 ( 
.A(n_790),
.Y(n_859)
);

BUFx2_ASAP7_75t_SL g860 ( 
.A(n_787),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_L g861 ( 
.A1(n_812),
.A2(n_777),
.B1(n_820),
.B2(n_823),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_808),
.Y(n_862)
);

INVx6_ASAP7_75t_L g863 ( 
.A(n_790),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_813),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_813),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_808),
.B(n_389),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_800),
.A2(n_758),
.B1(n_403),
.B2(n_414),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_819),
.Y(n_868)
);

CKINVDCx11_ASAP7_75t_R g869 ( 
.A(n_817),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_818),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_818),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_801),
.Y(n_872)
);

CKINVDCx11_ASAP7_75t_R g873 ( 
.A(n_822),
.Y(n_873)
);

INVx6_ASAP7_75t_L g874 ( 
.A(n_799),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_SL g875 ( 
.A1(n_796),
.A2(n_816),
.B1(n_788),
.B2(n_783),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_805),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_803),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_784),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_806),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_816),
.A2(n_403),
.B(n_414),
.Y(n_880)
);

BUFx2_ASAP7_75t_SL g881 ( 
.A(n_779),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_878),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_872),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_832),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_855),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_838),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_826),
.A2(n_804),
.B1(n_263),
.B2(n_253),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_875),
.A2(n_810),
.B(n_771),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_835),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_855),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_877),
.B(n_803),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_877),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_825),
.Y(n_893)
);

HB1xp67_ASAP7_75t_SL g894 ( 
.A(n_835),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_876),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_833),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_833),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_861),
.A2(n_826),
.B(n_834),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_841),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_841),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_876),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_878),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_878),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_878),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_837),
.Y(n_905)
);

INVx3_ASAP7_75t_SL g906 ( 
.A(n_844),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_840),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_842),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_862),
.B(n_770),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_862),
.B(n_795),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_864),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_837),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_865),
.B(n_792),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_881),
.B(n_824),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_856),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_829),
.B(n_3),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_829),
.B(n_5),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_893),
.B(n_839),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_893),
.B(n_868),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_889),
.B(n_851),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_889),
.B(n_851),
.Y(n_921)
);

OA21x2_ASAP7_75t_L g922 ( 
.A1(n_888),
.A2(n_871),
.B(n_870),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_898),
.A2(n_831),
.B1(n_848),
.B2(n_847),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_898),
.A2(n_853),
.B(n_857),
.Y(n_924)
);

AOI221xp5_ASAP7_75t_L g925 ( 
.A1(n_916),
.A2(n_849),
.B1(n_836),
.B2(n_866),
.C(n_867),
.Y(n_925)
);

NOR2x1_ASAP7_75t_SL g926 ( 
.A(n_917),
.B(n_845),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_885),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_884),
.B(n_862),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_884),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_882),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_887),
.A2(n_853),
.B(n_857),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_910),
.B(n_852),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_885),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_886),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_886),
.B(n_854),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_883),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_915),
.B(n_830),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_895),
.B(n_852),
.Y(n_938)
);

OA21x2_ASAP7_75t_L g939 ( 
.A1(n_888),
.A2(n_879),
.B(n_880),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_896),
.A2(n_850),
.B(n_874),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_894),
.Y(n_941)
);

NAND4xp25_ASAP7_75t_L g942 ( 
.A(n_917),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_895),
.B(n_844),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_908),
.Y(n_944)
);

AOI21xp33_ASAP7_75t_SL g945 ( 
.A1(n_906),
.A2(n_6),
.B(n_7),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_883),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_SL g947 ( 
.A1(n_917),
.A2(n_828),
.B(n_869),
.C(n_11),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_901),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_887),
.A2(n_907),
.B1(n_915),
.B2(n_905),
.Y(n_949)
);

AO21x1_ASAP7_75t_L g950 ( 
.A1(n_916),
.A2(n_8),
.B(n_9),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_915),
.B(n_827),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_SL g952 ( 
.A1(n_889),
.A2(n_874),
.B1(n_843),
.B2(n_827),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_908),
.B(n_827),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_911),
.B(n_827),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_885),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_882),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_905),
.B(n_843),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_932),
.B(n_901),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_922),
.B(n_928),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_929),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_923),
.A2(n_894),
.B1(n_874),
.B2(n_912),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_922),
.B(n_928),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_924),
.A2(n_907),
.B1(n_912),
.B2(n_902),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_944),
.B(n_911),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_944),
.B(n_911),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_936),
.B(n_913),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_927),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_948),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_922),
.B(n_913),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_929),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_934),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_932),
.B(n_904),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_930),
.B(n_909),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_948),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_922),
.B(n_913),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_932),
.B(n_904),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_936),
.B(n_891),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_927),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_932),
.B(n_909),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_930),
.B(n_909),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_930),
.B(n_909),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_927),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_979),
.B(n_938),
.Y(n_983)
);

OAI21xp33_ASAP7_75t_L g984 ( 
.A1(n_969),
.A2(n_942),
.B(n_918),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_961),
.A2(n_950),
.B1(n_942),
.B2(n_924),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_SL g986 ( 
.A(n_961),
.B(n_950),
.C(n_945),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_968),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_979),
.B(n_938),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_974),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_969),
.A2(n_947),
.B1(n_945),
.B2(n_923),
.C(n_931),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_960),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_979),
.B(n_943),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_977),
.B(n_964),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_960),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_958),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_959),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_958),
.B(n_943),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_977),
.B(n_964),
.Y(n_998)
);

OAI33xp33_ASAP7_75t_L g999 ( 
.A1(n_966),
.A2(n_919),
.A3(n_937),
.B1(n_934),
.B2(n_946),
.B3(n_957),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_969),
.B(n_946),
.Y(n_1000)
);

AOI31xp33_ASAP7_75t_L g1001 ( 
.A1(n_975),
.A2(n_941),
.A3(n_921),
.B(n_920),
.Y(n_1001)
);

BUFx2_ASAP7_75t_SL g1002 ( 
.A(n_959),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_959),
.B(n_937),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_1002),
.B(n_962),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_987),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_1002),
.B(n_962),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_995),
.B(n_962),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_993),
.B(n_966),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_989),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_995),
.B(n_976),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_996),
.B(n_973),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_983),
.B(n_976),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_993),
.B(n_965),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_991),
.Y(n_1014)
);

NOR2x1p5_ASAP7_75t_L g1015 ( 
.A(n_1009),
.B(n_986),
.Y(n_1015)
);

NAND4xp25_ASAP7_75t_L g1016 ( 
.A(n_1004),
.B(n_990),
.C(n_984),
.D(n_985),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_1008),
.B(n_998),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_1010),
.B(n_992),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1010),
.B(n_992),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1012),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1008),
.B(n_998),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1018),
.B(n_1007),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1019),
.B(n_1007),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1017),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_984),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_1025),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1022),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_1024),
.B(n_1015),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1022),
.B(n_1016),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_1023),
.B(n_1021),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1023),
.B(n_1014),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1024),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_1025),
.A2(n_990),
.B(n_1001),
.C(n_986),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1024),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_1025),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1024),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1035),
.B(n_1020),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1026),
.B(n_1005),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_1032),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1033),
.A2(n_1029),
.B(n_1028),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1027),
.B(n_1014),
.Y(n_1041)
);

NAND2x1_ASAP7_75t_L g1042 ( 
.A(n_1028),
.B(n_1004),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1030),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_SL g1044 ( 
.A(n_1029),
.B(n_1036),
.C(n_1034),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1031),
.B(n_1006),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1031),
.A2(n_999),
.B1(n_975),
.B2(n_1006),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_1035),
.A2(n_1001),
.B(n_1013),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_1035),
.B(n_989),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1033),
.A2(n_996),
.B1(n_1011),
.B2(n_1013),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1030),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1030),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1033),
.A2(n_975),
.B(n_996),
.Y(n_1052)
);

AOI22x1_ASAP7_75t_L g1053 ( 
.A1(n_1048),
.A2(n_1040),
.B1(n_1050),
.B2(n_1043),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1044),
.A2(n_1011),
.B(n_1000),
.Y(n_1054)
);

OAI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1046),
.A2(n_1052),
.B1(n_1049),
.B2(n_1047),
.Y(n_1055)
);

AND2x2_ASAP7_75t_SL g1056 ( 
.A(n_1038),
.B(n_906),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1051),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1037),
.Y(n_1058)
);

OAI31xp33_ASAP7_75t_L g1059 ( 
.A1(n_1039),
.A2(n_1003),
.A3(n_1000),
.B(n_989),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1041),
.Y(n_1060)
);

AOI21xp33_ASAP7_75t_SL g1061 ( 
.A1(n_1045),
.A2(n_906),
.B(n_987),
.Y(n_1061)
);

AOI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1046),
.A2(n_963),
.B1(n_1003),
.B2(n_925),
.C(n_931),
.Y(n_1062)
);

OAI211xp5_ASAP7_75t_L g1063 ( 
.A1(n_1042),
.A2(n_869),
.B(n_873),
.C(n_1012),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1048),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1043),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1044),
.A2(n_994),
.B1(n_991),
.B2(n_1011),
.C(n_949),
.Y(n_1066)
);

AOI222xp33_ASAP7_75t_L g1067 ( 
.A1(n_1044),
.A2(n_926),
.B1(n_965),
.B2(n_994),
.C1(n_906),
.C2(n_1011),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1043),
.B(n_997),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1043),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1043),
.Y(n_1070)
);

AO22x2_ASAP7_75t_L g1071 ( 
.A1(n_1044),
.A2(n_997),
.B1(n_988),
.B2(n_983),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_1057),
.B(n_953),
.C(n_970),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1053),
.A2(n_926),
.B(n_939),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_1063),
.B(n_11),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1068),
.B(n_988),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1060),
.B(n_970),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1056),
.B(n_980),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1064),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1058),
.B(n_873),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1055),
.A2(n_1062),
.B1(n_1071),
.B2(n_1069),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1065),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1070),
.B(n_971),
.Y(n_1082)
);

NAND5xp2_ASAP7_75t_L g1083 ( 
.A(n_1067),
.B(n_952),
.C(n_846),
.D(n_858),
.E(n_980),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1071),
.Y(n_1084)
);

NAND4xp25_ASAP7_75t_L g1085 ( 
.A(n_1067),
.B(n_981),
.C(n_980),
.D(n_973),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1054),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1066),
.B(n_971),
.Y(n_1087)
);

NOR3x1_ASAP7_75t_L g1088 ( 
.A(n_1061),
.B(n_12),
.C(n_13),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1080),
.A2(n_1059),
.B(n_939),
.Y(n_1089)
);

XOR2x2_ASAP7_75t_L g1090 ( 
.A(n_1074),
.B(n_1059),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_SL g1091 ( 
.A(n_1078),
.B(n_859),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1081),
.B(n_935),
.Y(n_1092)
);

OAI21xp33_ASAP7_75t_L g1093 ( 
.A1(n_1083),
.A2(n_981),
.B(n_973),
.Y(n_1093)
);

AOI211xp5_ASAP7_75t_SL g1094 ( 
.A1(n_1084),
.A2(n_12),
.B(n_15),
.C(n_16),
.Y(n_1094)
);

AOI211xp5_ASAP7_75t_L g1095 ( 
.A1(n_1079),
.A2(n_976),
.B(n_972),
.C(n_981),
.Y(n_1095)
);

AOI32xp33_ASAP7_75t_L g1096 ( 
.A1(n_1086),
.A2(n_1087),
.A3(n_1088),
.B1(n_1077),
.B2(n_1082),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_1073),
.B(n_1076),
.C(n_1072),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1083),
.A2(n_939),
.B(n_17),
.C(n_18),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1075),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_SL g1100 ( 
.A(n_1085),
.B(n_15),
.C(n_19),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_1078),
.B(n_859),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1078),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1084),
.A2(n_940),
.B1(n_935),
.B2(n_902),
.C(n_954),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1078),
.B(n_19),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1074),
.A2(n_939),
.B(n_973),
.Y(n_1105)
);

AOI221xp5_ASAP7_75t_L g1106 ( 
.A1(n_1084),
.A2(n_940),
.B1(n_902),
.B2(n_954),
.C(n_263),
.Y(n_1106)
);

OAI211xp5_ASAP7_75t_L g1107 ( 
.A1(n_1080),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_SL g1108 ( 
.A(n_1080),
.B(n_847),
.C(n_169),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1074),
.A2(n_973),
.B(n_972),
.Y(n_1109)
);

OAI221xp5_ASAP7_75t_SL g1110 ( 
.A1(n_1080),
.A2(n_914),
.B1(n_951),
.B2(n_930),
.C(n_956),
.Y(n_1110)
);

NAND4xp25_ASAP7_75t_L g1111 ( 
.A(n_1080),
.B(n_956),
.C(n_21),
.D(n_23),
.Y(n_1111)
);

AOI222xp33_ASAP7_75t_L g1112 ( 
.A1(n_1084),
.A2(n_982),
.B1(n_978),
.B2(n_967),
.C1(n_907),
.C2(n_263),
.Y(n_1112)
);

XNOR2xp5_ASAP7_75t_L g1113 ( 
.A(n_1090),
.B(n_20),
.Y(n_1113)
);

AOI211xp5_ASAP7_75t_L g1114 ( 
.A1(n_1102),
.A2(n_23),
.B(n_24),
.C(n_27),
.Y(n_1114)
);

AOI321xp33_ASAP7_75t_L g1115 ( 
.A1(n_1110),
.A2(n_891),
.A3(n_951),
.B1(n_967),
.B2(n_978),
.C(n_982),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1099),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_SL g1117 ( 
.A(n_1107),
.B(n_171),
.C(n_167),
.Y(n_1117)
);

NAND4xp25_ASAP7_75t_SL g1118 ( 
.A(n_1096),
.B(n_1097),
.C(n_1098),
.D(n_1095),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_1089),
.A2(n_940),
.B1(n_177),
.B2(n_231),
.C(n_180),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1104),
.Y(n_1120)
);

AOI211xp5_ASAP7_75t_L g1121 ( 
.A1(n_1111),
.A2(n_1108),
.B(n_1091),
.C(n_1101),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1094),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_1092),
.B(n_28),
.Y(n_1123)
);

OAI211xp5_ASAP7_75t_L g1124 ( 
.A1(n_1100),
.A2(n_1093),
.B(n_1105),
.C(n_1106),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1112),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1109),
.A2(n_956),
.B1(n_903),
.B2(n_863),
.Y(n_1126)
);

NAND2x1_ASAP7_75t_SL g1127 ( 
.A(n_1103),
.B(n_29),
.Y(n_1127)
);

OAI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_1100),
.A2(n_956),
.B(n_903),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1107),
.A2(n_859),
.B1(n_863),
.B2(n_882),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_1089),
.A2(n_234),
.B1(n_185),
.B2(n_192),
.C(n_196),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1089),
.A2(n_882),
.B1(n_903),
.B2(n_891),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1089),
.A2(n_236),
.B1(n_199),
.B2(n_200),
.C(n_210),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1102),
.Y(n_1133)
);

BUFx2_ASAP7_75t_R g1134 ( 
.A(n_1102),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1090),
.A2(n_32),
.B(n_35),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1107),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_1136)
);

NAND4xp75_ASAP7_75t_L g1137 ( 
.A(n_1135),
.B(n_40),
.C(n_41),
.D(n_42),
.Y(n_1137)
);

NOR4xp75_ASAP7_75t_L g1138 ( 
.A(n_1127),
.B(n_43),
.C(n_44),
.D(n_45),
.Y(n_1138)
);

NAND4xp75_ASAP7_75t_L g1139 ( 
.A(n_1120),
.B(n_1133),
.C(n_1123),
.D(n_1130),
.Y(n_1139)
);

NAND4xp75_ASAP7_75t_L g1140 ( 
.A(n_1132),
.B(n_44),
.C(n_863),
.D(n_860),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1116),
.B(n_909),
.Y(n_1141)
);

NAND4xp75_ASAP7_75t_L g1142 ( 
.A(n_1119),
.B(n_982),
.C(n_978),
.D(n_967),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1134),
.B(n_910),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1122),
.B(n_843),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1113),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1136),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1114),
.B(n_910),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1121),
.B(n_910),
.Y(n_1148)
);

OAI322xp33_ASAP7_75t_L g1149 ( 
.A1(n_1125),
.A2(n_266),
.A3(n_211),
.B1(n_213),
.B2(n_216),
.C1(n_220),
.C2(n_221),
.Y(n_1149)
);

AO22x2_ASAP7_75t_L g1150 ( 
.A1(n_1117),
.A2(n_910),
.B1(n_903),
.B2(n_955),
.Y(n_1150)
);

AND2x2_ASAP7_75t_SL g1151 ( 
.A(n_1131),
.B(n_843),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1126),
.A2(n_882),
.B1(n_914),
.B2(n_933),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1124),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1118),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1129),
.B(n_914),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1128),
.B(n_882),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1115),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1116),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1158),
.B(n_182),
.Y(n_1159)
);

OAI322xp33_ASAP7_75t_L g1160 ( 
.A1(n_1153),
.A2(n_270),
.A3(n_225),
.B1(n_227),
.B2(n_228),
.C1(n_229),
.C2(n_235),
.Y(n_1160)
);

XNOR2x1_ASAP7_75t_L g1161 ( 
.A(n_1138),
.B(n_223),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1154),
.B(n_914),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_L g1163 ( 
.A(n_1145),
.B(n_275),
.C(n_268),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_L g1164 ( 
.A(n_1139),
.B(n_260),
.C(n_256),
.Y(n_1164)
);

NAND4xp75_ASAP7_75t_L g1165 ( 
.A(n_1146),
.B(n_1143),
.C(n_1144),
.D(n_1157),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1141),
.B(n_244),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1148),
.A2(n_1149),
.B1(n_1147),
.B2(n_1156),
.C(n_1152),
.Y(n_1167)
);

OAI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1150),
.A2(n_914),
.B1(n_250),
.B2(n_249),
.C(n_882),
.Y(n_1168)
);

OAI211xp5_ASAP7_75t_L g1169 ( 
.A1(n_1140),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_1169)
);

AOI211xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1141),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_1170)
);

AOI221x1_ASAP7_75t_L g1171 ( 
.A1(n_1150),
.A2(n_896),
.B1(n_61),
.B2(n_62),
.C(n_64),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1137),
.A2(n_914),
.B(n_65),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1155),
.B(n_1142),
.Y(n_1173)
);

AOI211xp5_ASAP7_75t_L g1174 ( 
.A1(n_1163),
.A2(n_1155),
.B(n_1151),
.C(n_955),
.Y(n_1174)
);

XNOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1161),
.B(n_59),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1165),
.Y(n_1176)
);

XNOR2xp5_ASAP7_75t_L g1177 ( 
.A(n_1169),
.B(n_1164),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1162),
.Y(n_1178)
);

AO22x2_ASAP7_75t_L g1179 ( 
.A1(n_1173),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1159),
.A2(n_955),
.B1(n_933),
.B2(n_890),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1166),
.Y(n_1181)
);

XNOR2x1_ASAP7_75t_L g1182 ( 
.A(n_1172),
.B(n_71),
.Y(n_1182)
);

NAND5xp2_ASAP7_75t_L g1183 ( 
.A(n_1167),
.B(n_73),
.C(n_74),
.D(n_76),
.E(n_78),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1170),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1160),
.B(n_933),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1168),
.A2(n_892),
.B1(n_890),
.B2(n_897),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1171),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1159),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1176),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1187),
.A2(n_892),
.B1(n_890),
.B2(n_897),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1184),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1178),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1179),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1175),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1179),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1185),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1182),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1181),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1192),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1198),
.A2(n_1177),
.B(n_1188),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_1191),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1189),
.A2(n_1183),
.B(n_1174),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1196),
.A2(n_1194),
.B1(n_1197),
.B2(n_1195),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1193),
.A2(n_1186),
.B1(n_1180),
.B2(n_892),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1201),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1199),
.A2(n_1194),
.B1(n_1190),
.B2(n_900),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1202),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1203),
.A2(n_900),
.B1(n_899),
.B2(n_897),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1207),
.A2(n_1200),
.B1(n_1204),
.B2(n_90),
.C(n_93),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1209),
.A2(n_1205),
.B(n_1206),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1210),
.A2(n_1208),
.B(n_85),
.Y(n_1211)
);

NOR2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1211),
.B(n_80),
.Y(n_1212)
);

OAI221xp5_ASAP7_75t_R g1213 ( 
.A1(n_1212),
.A2(n_96),
.B1(n_100),
.B2(n_102),
.C(n_105),
.Y(n_1213)
);

AOI211xp5_ASAP7_75t_L g1214 ( 
.A1(n_1213),
.A2(n_106),
.B(n_108),
.C(n_109),
.Y(n_1214)
);


endmodule