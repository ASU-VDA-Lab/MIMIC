module real_jpeg_23543_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_70),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_70),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_73),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx8_ASAP7_75t_SL g48 ( 
.A(n_6),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_8),
.B(n_52),
.C(n_64),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_79),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_119),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_57),
.B1(n_101),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_9),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_11),
.A2(n_26),
.B1(n_106),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_26),
.B1(n_52),
.B2(n_53),
.Y(n_159)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_20),
.B(n_87),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_61),
.C(n_75),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_21),
.A2(n_22),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_43),
.C(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_32),
.B2(n_39),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_25),
.A2(n_31),
.B1(n_78),
.B2(n_119),
.Y(n_178)
);

INVx5_ASAP7_75t_SL g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_29),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_27),
.B(n_79),
.CON(n_78),
.SN(n_78)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_27),
.B(n_34),
.C(n_37),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_27),
.A2(n_47),
.B(n_92),
.C(n_95),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_48),
.C(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_31),
.A2(n_40),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_32)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_33),
.A2(n_35),
.B(n_78),
.C(n_80),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_35),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_35),
.B(n_133),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_60),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_105),
.B1(n_109),
.B2(n_113),
.Y(n_104)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_46),
.B(n_110),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_47),
.A2(n_48),
.B1(n_96),
.B2(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_56),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_55),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_53),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_54),
.A2(n_84),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_55),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_57),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_57),
.A2(n_86),
.B1(n_152),
.B2(n_159),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_61),
.A2(n_75),
.B1(n_76),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_61),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_68),
.B(n_71),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_62),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_62),
.A2(n_67),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_62),
.A2(n_67),
.B1(n_137),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_67),
.B(n_79),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_69),
.A2(n_74),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_74),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_77),
.A2(n_81),
.B1(n_82),
.B2(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_77),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_93),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_92),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_79),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_102),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_103),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_181),
.B(n_187),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_170),
.B(n_180),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_148),
.B(n_169),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_156),
.B(n_168),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_154),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_164),
.B(n_167),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_166),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_179),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_175),
.C(n_178),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_182),
.B(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);


endmodule