module fake_jpeg_16798_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_5),
.B(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_26),
.B1(n_24),
.B2(n_28),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_33),
.Y(n_59)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_66),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_69),
.B1(n_73),
.B2(n_42),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_36),
.B1(n_32),
.B2(n_40),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_36),
.B1(n_21),
.B2(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_21),
.B1(n_32),
.B2(n_31),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_79),
.Y(n_111)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_34),
.C(n_55),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_95),
.B(n_16),
.Y(n_127)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_43),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_43),
.Y(n_124)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_96),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_25),
.B(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_29),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_107),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_64),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_110),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_49),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_112),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_60),
.A2(n_23),
.B(n_31),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_118),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_101),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_70),
.B1(n_78),
.B2(n_77),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_83),
.B1(n_44),
.B2(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_70),
.Y(n_118)
);

BUFx16f_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_126),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_33),
.B1(n_43),
.B2(n_49),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_108),
.B1(n_99),
.B2(n_109),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_130),
.B(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_29),
.Y(n_126)
);

AOI22x1_ASAP7_75t_R g141 ( 
.A1(n_127),
.A2(n_101),
.B1(n_110),
.B2(n_97),
.Y(n_141)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_53),
.B1(n_79),
.B2(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_137),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_15),
.B(n_1),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_93),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_99),
.B1(n_109),
.B2(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_53),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_44),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_105),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_144),
.C(n_165),
.Y(n_187)
);

XNOR2x2_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_15),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_75),
.B1(n_102),
.B2(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_149),
.B1(n_152),
.B2(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_44),
.B1(n_111),
.B2(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_161),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_124),
.B1(n_132),
.B2(n_115),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_167),
.Y(n_178)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_116),
.A3(n_122),
.B1(n_139),
.B2(n_135),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_126),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_83),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_16),
.B1(n_24),
.B2(n_12),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_15),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_115),
.A2(n_30),
.B1(n_27),
.B2(n_18),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_130),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_119),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_137),
.B1(n_138),
.B2(n_130),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_22),
.B1(n_15),
.B2(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_181),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_184),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_177),
.B(n_182),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_121),
.A3(n_120),
.B1(n_119),
.B2(n_30),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_128),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_133),
.B(n_128),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_143),
.A2(n_125),
.B1(n_30),
.B2(n_27),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_188),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_142),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_125),
.B1(n_30),
.B2(n_133),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_195),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_22),
.B1(n_15),
.B2(n_2),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_18),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_22),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_151),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_151),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_140),
.B(n_6),
.C(n_11),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_144),
.C(n_162),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_208),
.C(n_225),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_205),
.B(n_217),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_170),
.Y(n_208)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_215),
.B1(n_219),
.B2(n_173),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_157),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_181),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_180),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_177),
.B1(n_195),
.B2(n_191),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_157),
.B1(n_168),
.B2(n_152),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_224),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_168),
.C(n_165),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_182),
.B1(n_218),
.B2(n_172),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_234),
.B1(n_207),
.B2(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_228),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_238),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_172),
.B1(n_197),
.B2(n_177),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_192),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_179),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_188),
.B1(n_216),
.B2(n_185),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_201),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_175),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_194),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_8),
.B1(n_11),
.B2(n_3),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_208),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_252),
.C(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_262),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_230),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_213),
.B1(n_216),
.B2(n_225),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_253),
.B1(n_255),
.B2(n_236),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_243),
.C(n_235),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_226),
.B1(n_242),
.B2(n_231),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_234),
.A2(n_203),
.B1(n_190),
.B2(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_227),
.B(n_171),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_239),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_171),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_261),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_270),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_241),
.B(n_227),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_268),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_273),
.C(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_211),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_274),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_236),
.B(n_230),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_254),
.B(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_184),
.C(n_1),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_184),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_0),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_283),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_248),
.B1(n_249),
.B2(n_255),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_282),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_4),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_287),
.Y(n_292)
);

OAI21x1_ASAP7_75t_SL g285 ( 
.A1(n_273),
.A2(n_4),
.B(n_6),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_9),
.B(n_10),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_6),
.B(n_8),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_14),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_293),
.Y(n_299)
);

HAxp5_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_263),
.CON(n_293),
.SN(n_293)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_295),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_9),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_290),
.B(n_293),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_284),
.C(n_281),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_303),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_14),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_304),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_296),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_308),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_294),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_305),
.B(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_307),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_312),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_306),
.Y(n_315)
);


endmodule