module fake_jpeg_13048_n_567 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_567);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_567;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_54),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_55),
.Y(n_155)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_70),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx2_ASAP7_75t_SL g161 ( 
.A(n_62),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_18),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_9),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_49),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_9),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_83),
.Y(n_129)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_10),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_10),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g162 ( 
.A(n_106),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_52),
.B1(n_21),
.B2(n_23),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_115),
.A2(n_121),
.B1(n_125),
.B2(n_132),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_30),
.B1(n_21),
.B2(n_44),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_34),
.B1(n_43),
.B2(n_20),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_23),
.B1(n_31),
.B2(n_41),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_127),
.A2(n_137),
.B1(n_145),
.B2(n_149),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_48),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_20),
.B1(n_24),
.B2(n_33),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_43),
.B1(n_34),
.B2(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_33),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_140),
.B(n_165),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_60),
.A2(n_43),
.B1(n_34),
.B2(n_42),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_72),
.A2(n_43),
.B1(n_34),
.B2(n_42),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_72),
.A2(n_43),
.B1(n_34),
.B2(n_41),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_154),
.B1(n_104),
.B2(n_100),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_49),
.B1(n_31),
.B2(n_36),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_129),
.B1(n_162),
.B2(n_147),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_74),
.A2(n_77),
.B1(n_65),
.B2(n_85),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_53),
.B(n_36),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_54),
.B(n_11),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_168),
.B(n_48),
.Y(n_215)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_172),
.A2(n_121),
.B1(n_150),
.B2(n_125),
.Y(n_239)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_173),
.Y(n_250)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g274 ( 
.A(n_174),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_179),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_180),
.Y(n_280)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_186),
.Y(n_265)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_124),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_108),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_187),
.B(n_200),
.Y(n_287)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_190),
.Y(n_276)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_77),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_193),
.B(n_195),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_194),
.A2(n_207),
.B1(n_210),
.B2(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_74),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_196),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_111),
.B(n_112),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_197),
.B(n_198),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_119),
.B(n_0),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_202),
.B(n_214),
.Y(n_281)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_133),
.Y(n_203)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_120),
.B(n_48),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_208),
.Y(n_252)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_211),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_127),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_123),
.B(n_0),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_138),
.B(n_26),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_118),
.B(n_48),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_216),
.B(n_220),
.Y(n_285)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_219),
.Y(n_273)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_111),
.B(n_17),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_112),
.B(n_1),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_222),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_156),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_226),
.Y(n_279)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_128),
.B(n_1),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_158),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_228),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_169),
.B(n_88),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_230),
.B(n_221),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_137),
.A2(n_145),
.B(n_149),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_152),
.B(n_62),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_232),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_239),
.B(n_278),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_175),
.A2(n_212),
.B1(n_232),
.B2(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_240),
.A2(n_216),
.B1(n_208),
.B2(n_190),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_166),
.B(n_164),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_177),
.B(n_203),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_191),
.A2(n_134),
.B1(n_159),
.B2(n_141),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_243),
.A2(n_268),
.B1(n_186),
.B2(n_187),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_191),
.A2(n_148),
.B1(n_152),
.B2(n_138),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_244),
.A2(n_259),
.B1(n_226),
.B2(n_184),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_249),
.A2(n_282),
.B(n_27),
.Y(n_329)
);

AO22x2_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_134),
.B1(n_159),
.B2(n_141),
.Y(n_251)
);

AO22x1_ASAP7_75t_SL g314 ( 
.A1(n_251),
.A2(n_209),
.B1(n_218),
.B2(n_199),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_201),
.B(n_213),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_261),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_175),
.A2(n_156),
.B1(n_143),
.B2(n_163),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_143),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_267),
.B(n_2),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_202),
.A2(n_167),
.B1(n_87),
.B2(n_86),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_220),
.B(n_167),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_228),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_202),
.A2(n_59),
.B(n_27),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_174),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_198),
.Y(n_297)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_296),
.Y(n_365)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_216),
.A3(n_189),
.B1(n_173),
.B2(n_225),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_291),
.B(n_282),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_271),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g350 ( 
.A1(n_293),
.A2(n_234),
.B(n_256),
.Y(n_350)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_287),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_305),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_243),
.A2(n_68),
.B1(n_79),
.B2(n_217),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_297),
.B(n_304),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_192),
.C(n_208),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_299),
.B(n_327),
.C(n_333),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_240),
.A2(n_171),
.B1(n_200),
.B2(n_196),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_300),
.A2(n_308),
.B1(n_330),
.B2(n_233),
.Y(n_361)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_302),
.Y(n_341)
);

AO22x1_ASAP7_75t_L g344 ( 
.A1(n_303),
.A2(n_314),
.B1(n_286),
.B2(n_257),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_269),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_239),
.A2(n_183),
.B1(n_206),
.B2(n_222),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_238),
.A2(n_188),
.B1(n_207),
.B2(n_176),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_309),
.A2(n_313),
.B1(n_331),
.B2(n_337),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_251),
.A2(n_181),
.B1(n_205),
.B2(n_224),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_310),
.A2(n_263),
.B1(n_245),
.B2(n_253),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_317),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_238),
.A2(n_229),
.B1(n_185),
.B2(n_210),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_211),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_236),
.B(n_1),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_318),
.B(n_334),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_284),
.A2(n_11),
.B1(n_18),
.B2(n_4),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_319),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_265),
.B(n_11),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_320),
.B(n_323),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_249),
.A2(n_10),
.B(n_17),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_321),
.A2(n_324),
.B(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_322),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_281),
.A2(n_252),
.B1(n_269),
.B2(n_251),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_242),
.A2(n_3),
.B(n_27),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_326),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_27),
.C(n_3),
.Y(n_327)
);

OAI21x1_ASAP7_75t_SL g328 ( 
.A1(n_237),
.A2(n_27),
.B(n_4),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_329),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_12),
.B1(n_4),
.B2(n_6),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_241),
.A2(n_237),
.B1(n_273),
.B2(n_251),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_332),
.B(n_336),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_258),
.B(n_12),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_261),
.B(n_277),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_264),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_254),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_267),
.B(n_3),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_251),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_317),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_342),
.B(n_346),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_324),
.A2(n_252),
.B1(n_268),
.B2(n_275),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_348),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_344),
.A2(n_350),
.B(n_363),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_309),
.Y(n_346)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_336),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_275),
.B1(n_279),
.B2(n_254),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_280),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_355),
.C(n_358),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_260),
.Y(n_355)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_270),
.C(n_283),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_334),
.A2(n_270),
.B1(n_233),
.B2(n_272),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_369),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_318),
.B(n_274),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_360),
.B(n_362),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_361),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_295),
.B(n_274),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_290),
.A2(n_300),
.B(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_305),
.A2(n_255),
.B1(n_247),
.B2(n_253),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_283),
.C(n_235),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_380),
.C(n_294),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_235),
.C(n_274),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_382),
.B(n_388),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_L g383 ( 
.A1(n_370),
.A2(n_290),
.B(n_291),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_383),
.B(n_341),
.C(n_340),
.Y(n_449)
);

AOI322xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_289),
.A3(n_337),
.B1(n_321),
.B2(n_313),
.C1(n_314),
.C2(n_328),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_329),
.B(n_303),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_343),
.B(n_351),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_375),
.A2(n_312),
.B1(n_314),
.B2(n_325),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_392),
.A2(n_402),
.B1(n_407),
.B2(n_411),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_393),
.B(n_353),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_353),
.Y(n_429)
);

AO22x1_ASAP7_75t_SL g395 ( 
.A1(n_377),
.A2(n_322),
.B1(n_332),
.B2(n_301),
.Y(n_395)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_395),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_377),
.A2(n_315),
.B(n_326),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_396),
.A2(n_403),
.B(n_405),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_302),
.C(n_306),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_410),
.C(n_412),
.Y(n_428)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_398),
.Y(n_447)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_400),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_288),
.B1(n_296),
.B2(n_330),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_374),
.A2(n_307),
.B(n_274),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_344),
.A2(n_292),
.B(n_335),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_339),
.Y(n_406)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_406),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_365),
.A2(n_255),
.B1(n_316),
.B2(n_247),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_338),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_414),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_348),
.A2(n_264),
.B1(n_248),
.B2(n_245),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_409),
.A2(n_376),
.B1(n_346),
.B2(n_345),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_355),
.B(n_248),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_365),
.A2(n_255),
.B1(n_247),
.B2(n_263),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_354),
.B(n_347),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_381),
.B(n_263),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_413),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_357),
.B(n_17),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_357),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_416),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_359),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_8),
.Y(n_417)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_369),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_419),
.Y(n_425)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_420),
.B(n_438),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_426),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_404),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_397),
.C(n_410),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_433),
.B1(n_436),
.B2(n_441),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_391),
.A2(n_376),
.B(n_344),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_444),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_405),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_385),
.A2(n_363),
.B1(n_368),
.B2(n_360),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_385),
.A2(n_363),
.B1(n_350),
.B2(n_367),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_412),
.B(n_371),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_408),
.A2(n_373),
.B1(n_366),
.B2(n_378),
.Y(n_439)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_384),
.B(n_380),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_448),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_416),
.A2(n_366),
.B1(n_361),
.B2(n_372),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_384),
.B(n_378),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_446),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_404),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_393),
.B(n_372),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_394),
.B(n_341),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_401),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_399),
.A2(n_349),
.B1(n_352),
.B2(n_345),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_451),
.A2(n_452),
.B1(n_418),
.B2(n_419),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_392),
.A2(n_349),
.B1(n_352),
.B2(n_379),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_456),
.C(n_474),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_450),
.Y(n_454)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_454),
.Y(n_489)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_447),
.Y(n_455)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_403),
.C(n_396),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_458),
.A2(n_424),
.B1(n_421),
.B2(n_436),
.Y(n_484)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_386),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_461),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_386),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_469),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_441),
.A2(n_415),
.B1(n_402),
.B2(n_407),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_463),
.A2(n_445),
.B1(n_452),
.B2(n_421),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_387),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_472),
.Y(n_494)
);

NOR3xp33_ASAP7_75t_SL g469 ( 
.A(n_437),
.B(n_417),
.C(n_414),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_470),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_413),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_429),
.B(n_401),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_476),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_395),
.C(n_390),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_409),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_480),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_423),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_395),
.C(n_390),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_478),
.C(n_422),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_420),
.B(n_395),
.C(n_406),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_435),
.B(n_433),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_479),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_400),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_481),
.A2(n_493),
.B1(n_500),
.B2(n_470),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_471),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_492),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_456),
.A2(n_432),
.B1(n_431),
.B2(n_443),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_460),
.A2(n_445),
.B1(n_425),
.B2(n_451),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_443),
.C(n_434),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_499),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_468),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_501),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_434),
.C(n_427),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_460),
.A2(n_389),
.B1(n_427),
.B2(n_447),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_467),
.B(n_411),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_389),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_480),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_464),
.A2(n_398),
.B1(n_379),
.B2(n_16),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_503),
.B(n_455),
.Y(n_516)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_504),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_512),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_490),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_510),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_485),
.B(n_457),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_509),
.B(n_516),
.Y(n_530)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_491),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_482),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_511),
.B(n_515),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_495),
.B(n_465),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_513),
.B(n_519),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_493),
.A2(n_475),
.B1(n_477),
.B2(n_478),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_514),
.Y(n_527)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_500),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_517),
.B(n_520),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_486),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_496),
.B(n_466),
.C(n_465),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_466),
.C(n_483),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_513),
.A2(n_481),
.B1(n_487),
.B2(n_488),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_522),
.A2(n_533),
.B1(n_514),
.B2(n_527),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_525),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_483),
.C(n_499),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_506),
.A2(n_492),
.B(n_502),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_526),
.A2(n_529),
.B(n_524),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_498),
.C(n_494),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_505),
.A2(n_484),
.B(n_463),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_532),
.A2(n_521),
.B1(n_507),
.B2(n_512),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_520),
.A2(n_495),
.B1(n_501),
.B2(n_469),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_530),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_541),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_538),
.Y(n_552)
);

INVxp33_ASAP7_75t_SL g550 ( 
.A(n_540),
.Y(n_550)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_534),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_542),
.B(n_543),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_507),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_532),
.A2(n_528),
.B1(n_523),
.B2(n_531),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_544),
.B(n_545),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_519),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_529),
.A2(n_494),
.B(n_15),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_547),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_535),
.B(n_13),
.Y(n_547)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_539),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_549),
.B(n_551),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_555),
.B(n_556),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_554),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_550),
.B(n_544),
.C(n_543),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_557),
.A2(n_558),
.B(n_553),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_552),
.A2(n_536),
.B(n_540),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_559),
.A2(n_561),
.B(n_548),
.Y(n_562)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g561 ( 
.A1(n_558),
.A2(n_532),
.B(n_553),
.C(n_533),
.D(n_528),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_562),
.B(n_563),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_560),
.B(n_13),
.C(n_15),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_13),
.B(n_15),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_565),
.A2(n_13),
.B(n_15),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_566),
.B(n_16),
.Y(n_567)
);


endmodule