module fake_jpeg_3232_n_576 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_576);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_576;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_58),
.B(n_74),
.Y(n_140)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_59),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_61),
.B(n_68),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_0),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_70),
.B(n_77),
.Y(n_154)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_75),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_33),
.B(n_2),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_79),
.B(n_91),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_20),
.B(n_4),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_80),
.B(n_84),
.Y(n_157)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_86),
.B(n_90),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_27),
.B(n_4),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_102),
.Y(n_163)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_95),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_20),
.B(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_96),
.B(n_97),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_22),
.B(n_6),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_98),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_100),
.B(n_110),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_40),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_40),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_103),
.B(n_104),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_6),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_23),
.B(n_6),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

BUFx16f_ASAP7_75t_L g120 ( 
.A(n_19),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_57),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_124),
.Y(n_171)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_19),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_39),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_52),
.B1(n_32),
.B2(n_29),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_128),
.A2(n_132),
.B1(n_164),
.B2(n_188),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_49),
.B1(n_125),
.B2(n_123),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_66),
.A2(n_113),
.B1(n_112),
.B2(n_111),
.Y(n_132)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g267 ( 
.A(n_141),
.Y(n_267)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_63),
.A2(n_49),
.B1(n_25),
.B2(n_29),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_150),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_76),
.A2(n_21),
.B1(n_55),
.B2(n_54),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_151),
.B(n_130),
.Y(n_285)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_152),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_75),
.A2(n_49),
.B1(n_25),
.B2(n_44),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_73),
.B(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_159),
.B(n_162),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_82),
.A2(n_32),
.B1(n_44),
.B2(n_21),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_85),
.A2(n_32),
.B1(n_44),
.B2(n_54),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_166),
.A2(n_182),
.B(n_207),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_104),
.A2(n_26),
.B1(n_55),
.B2(n_51),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_167),
.A2(n_172),
.B1(n_193),
.B2(n_194),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_67),
.A2(n_23),
.B1(n_51),
.B2(n_39),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_174),
.B(n_178),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_92),
.B(n_38),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_176),
.B(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_71),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_38),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_185),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_59),
.A2(n_37),
.B1(n_35),
.B2(n_28),
.Y(n_182)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_69),
.B(n_37),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_64),
.A2(n_35),
.B1(n_26),
.B2(n_56),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_89),
.A2(n_56),
.B1(n_46),
.B2(n_9),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_65),
.A2(n_56),
.B1(n_8),
.B2(n_9),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_93),
.B(n_7),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_105),
.A2(n_56),
.B1(n_8),
.B2(n_9),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_198),
.A2(n_206),
.B1(n_14),
.B2(n_15),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_94),
.B(n_7),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_200),
.B(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_201),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_119),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_106),
.B(n_116),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_114),
.C(n_108),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_215),
.B(n_218),
.C(n_235),
.Y(n_326)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_217),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_62),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_149),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_219),
.B(n_232),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_72),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_227),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_149),
.A2(n_98),
.B(n_109),
.C(n_107),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_221),
.A2(n_284),
.B(n_191),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g224 ( 
.A(n_163),
.B(n_117),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_224),
.A2(n_252),
.B(n_271),
.Y(n_311)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_225),
.Y(n_325)
);

AO22x2_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_117),
.B1(n_87),
.B2(n_83),
.Y(n_226)
);

AO21x2_ASAP7_75t_L g314 ( 
.A1(n_226),
.A2(n_212),
.B(n_222),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_87),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_11),
.C(n_13),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_228),
.B(n_262),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_229),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_69),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_231),
.B(n_248),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_171),
.Y(n_232)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_234),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_143),
.B(n_83),
.C(n_14),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_157),
.B(n_11),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_161),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_239),
.B(n_242),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_241),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_204),
.Y(n_242)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_133),
.Y(n_245)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_245),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_188),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_246),
.A2(n_258),
.B1(n_250),
.B2(n_233),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_247),
.A2(n_276),
.B1(n_222),
.B2(n_277),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_14),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_140),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_249),
.B(n_257),
.Y(n_320)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_128),
.Y(n_250)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_127),
.Y(n_251)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

OAI32xp33_ASAP7_75t_L g252 ( 
.A1(n_142),
.A2(n_189),
.A3(n_146),
.B1(n_137),
.B2(n_134),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_158),
.Y(n_255)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_255),
.Y(n_331)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_256),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_156),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_132),
.A2(n_155),
.B1(n_164),
.B2(n_206),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_175),
.B(n_195),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_259),
.B(n_273),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_187),
.Y(n_260)
);

INVx11_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

BUFx12f_ASAP7_75t_SL g317 ( 
.A(n_261),
.Y(n_317)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_186),
.B(n_196),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_265),
.B(n_272),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_145),
.B(n_213),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_269),
.B(n_283),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_270),
.Y(n_327)
);

OR2x4_ASAP7_75t_L g271 ( 
.A(n_182),
.B(n_131),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_145),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_169),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_208),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_274),
.B(n_286),
.Y(n_308)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_275),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_166),
.A2(n_150),
.B1(n_153),
.B2(n_207),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_278),
.B(n_285),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_199),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_212),
.B1(n_240),
.B2(n_260),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_129),
.B(n_135),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_130),
.A2(n_135),
.B(n_129),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_199),
.B(n_127),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_199),
.B(n_191),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_287),
.B(n_288),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_148),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_291),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_148),
.B1(n_138),
.B2(n_168),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_294),
.B(n_334),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g295 ( 
.A1(n_230),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_233),
.A2(n_282),
.B1(n_280),
.B2(n_277),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_136),
.B1(n_139),
.B2(n_147),
.Y(n_297)
);

OAI21x1_ASAP7_75t_SL g360 ( 
.A1(n_300),
.A2(n_283),
.B(n_221),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_230),
.A2(n_168),
.B(n_183),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_304),
.A2(n_260),
.B(n_253),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_183),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_312),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_321),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_218),
.B(n_203),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_227),
.B(n_203),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_342),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_328),
.B1(n_226),
.B2(n_284),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_241),
.Y(n_321)
);

OAI32xp33_ASAP7_75t_L g334 ( 
.A1(n_220),
.A2(n_252),
.A3(n_280),
.B1(n_268),
.B2(n_285),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g337 ( 
.A1(n_243),
.A2(n_238),
.A3(n_236),
.B1(n_224),
.B2(n_248),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_343),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_269),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_338),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_269),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_283),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_248),
.B(n_224),
.Y(n_342)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_215),
.A2(n_244),
.A3(n_276),
.B1(n_226),
.B2(n_235),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_237),
.C(n_231),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_354),
.C(n_362),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_348),
.A2(n_350),
.B1(n_377),
.B2(n_295),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_328),
.A2(n_226),
.B1(n_247),
.B2(n_267),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_351),
.Y(n_411)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_279),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_291),
.A2(n_267),
.B1(n_217),
.B2(n_234),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_358),
.B1(n_374),
.B2(n_375),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_296),
.A2(n_231),
.B1(n_216),
.B2(n_223),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_360),
.A2(n_324),
.B(n_341),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_299),
.C(n_311),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_290),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_369),
.Y(n_400)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_299),
.B(n_279),
.C(n_245),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_289),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_366),
.A2(n_370),
.B(n_300),
.Y(n_396)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_310),
.Y(n_367)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_303),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_342),
.A2(n_253),
.B1(n_281),
.B2(n_275),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_323),
.B(n_278),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

AND2x2_ASAP7_75t_SL g372 ( 
.A(n_289),
.B(n_262),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_381),
.Y(n_394)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_314),
.A2(n_223),
.B1(n_266),
.B2(n_255),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_314),
.A2(n_266),
.B1(n_256),
.B2(n_265),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_311),
.B(n_272),
.C(n_281),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_340),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_314),
.A2(n_270),
.B1(n_251),
.B2(n_225),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_314),
.A2(n_261),
.B1(n_297),
.B2(n_313),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_378),
.A2(n_294),
.B1(n_304),
.B2(n_338),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_320),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_382),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_308),
.B(n_306),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_383),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_305),
.B(n_307),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_305),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_354),
.B(n_337),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_387),
.B(n_391),
.Y(n_427)
);

AO22x1_ASAP7_75t_L g389 ( 
.A1(n_344),
.A2(n_359),
.B1(n_350),
.B2(n_377),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_395),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_335),
.B(n_334),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_393),
.A2(n_396),
.B(n_403),
.Y(n_448)
);

XOR2x1_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_324),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_412),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_343),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_413),
.C(n_376),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_408),
.B1(n_414),
.B2(n_349),
.Y(n_431)
);

NAND2x1_ASAP7_75t_SL g405 ( 
.A(n_379),
.B(n_317),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_405),
.A2(n_416),
.B(n_403),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_355),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_355),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_344),
.A2(n_348),
.B1(n_378),
.B2(n_347),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_346),
.B(n_289),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_347),
.A2(n_316),
.B1(n_327),
.B2(n_330),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_419),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_344),
.A2(n_327),
.B1(n_298),
.B2(n_301),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_420),
.Y(n_434)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_368),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_422),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_414),
.A2(n_374),
.B1(n_375),
.B2(n_384),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_423),
.A2(n_431),
.B1(n_443),
.B2(n_399),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_357),
.Y(n_424)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_415),
.Y(n_425)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_400),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_430),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_397),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_384),
.C(n_364),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_444),
.C(n_446),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_373),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_435),
.B(n_438),
.Y(n_461)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_332),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_345),
.Y(n_439)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_352),
.Y(n_440)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_440),
.Y(n_467)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_351),
.Y(n_442)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_442),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_408),
.A2(n_366),
.B1(n_358),
.B2(n_360),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_401),
.B(n_372),
.C(n_370),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_398),
.C(n_387),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_332),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_447),
.B(n_410),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_372),
.C(n_380),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_405),
.C(n_404),
.Y(n_477)
);

XOR2x1_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_394),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_396),
.A2(n_365),
.B(n_367),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_405),
.B(n_420),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_427),
.B(n_391),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_454),
.B(n_430),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_435),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_474),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_468),
.C(n_433),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_424),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_393),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_464),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_427),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_409),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_465),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_434),
.A2(n_389),
.B1(n_399),
.B2(n_416),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_466),
.A2(n_471),
.B(n_436),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_389),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_472),
.A2(n_426),
.B1(n_442),
.B2(n_356),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_422),
.B(n_392),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_475),
.A2(n_451),
.B(n_448),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_449),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_394),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_SL g486 ( 
.A(n_478),
.B(n_450),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_482),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_475),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_488),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_431),
.B1(n_429),
.B2(n_443),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_484),
.A2(n_489),
.B1(n_490),
.B2(n_494),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_446),
.C(n_448),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_487),
.C(n_464),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_491),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_460),
.C(n_478),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_461),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_429),
.B1(n_423),
.B2(n_434),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_467),
.A2(n_434),
.B1(n_440),
.B2(n_426),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_438),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_492),
.B(n_497),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_493),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_458),
.A2(n_426),
.B1(n_439),
.B2(n_390),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_394),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_495),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_496),
.A2(n_499),
.B1(n_469),
.B2(n_456),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_473),
.B(n_447),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_452),
.B(n_441),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_501),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_477),
.B(n_437),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_503),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_498),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_484),
.A2(n_458),
.B1(n_457),
.B2(n_476),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_508),
.A2(n_511),
.B1(n_519),
.B2(n_407),
.Y(n_534)
);

A2O1A1Ixp33_ASAP7_75t_L g510 ( 
.A1(n_503),
.A2(n_457),
.B(n_471),
.C(n_476),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_495),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_470),
.C(n_468),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_512),
.B(n_514),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_454),
.C(n_469),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_456),
.C(n_453),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_518),
.B(n_491),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_494),
.A2(n_453),
.B1(n_479),
.B2(n_459),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g521 ( 
.A(n_500),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_496),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_502),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_336),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_506),
.A2(n_489),
.B1(n_490),
.B2(n_483),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_524),
.A2(n_532),
.B1(n_519),
.B2(n_504),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_525),
.A2(n_512),
.B(n_516),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_527),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_498),
.C(n_485),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_529),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_495),
.C(n_493),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_531),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_520),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_515),
.A2(n_481),
.B1(n_425),
.B2(n_421),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_508),
.A2(n_407),
.B1(n_404),
.B2(n_417),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_533),
.A2(n_534),
.B1(n_510),
.B2(n_520),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_509),
.B(n_381),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_411),
.Y(n_541)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_536),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_541),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_524),
.A2(n_513),
.B1(n_517),
.B2(n_505),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_539),
.A2(n_365),
.B1(n_329),
.B2(n_292),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_525),
.A2(n_411),
.B1(n_417),
.B2(n_514),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_540),
.A2(n_523),
.B1(n_301),
.B2(n_298),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_505),
.Y(n_543)
);

XNOR2x1_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_544),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_507),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_545),
.B(n_547),
.Y(n_552)
);

AO22x1_ASAP7_75t_L g549 ( 
.A1(n_537),
.A2(n_533),
.B1(n_522),
.B2(n_528),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_556),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_550),
.B(n_547),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_546),
.A2(n_526),
.B(n_353),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_554),
.B(n_555),
.Y(n_560)
);

AND2x4_ASAP7_75t_SL g555 ( 
.A(n_539),
.B(n_329),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_542),
.A2(n_331),
.B(n_333),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_538),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_561),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_544),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_562),
.A2(n_563),
.B(n_553),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_552),
.B(n_551),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_SL g564 ( 
.A1(n_555),
.A2(n_543),
.B(n_333),
.C(n_318),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_564),
.A2(n_556),
.B(n_325),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_558),
.A2(n_560),
.B(n_553),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_565),
.B(n_566),
.Y(n_572)
);

BUFx24_ASAP7_75t_SL g566 ( 
.A(n_560),
.Y(n_566)
);

INVxp33_ASAP7_75t_L g571 ( 
.A(n_567),
.Y(n_571)
);

A2O1A1O1Ixp25_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_549),
.B(n_555),
.C(n_319),
.D(n_293),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_570),
.A2(n_568),
.B1(n_318),
.B2(n_325),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_571),
.B(n_572),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_319),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_293),
.Y(n_576)
);


endmodule