module fake_netlist_6_2411_n_1625 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1625);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1625;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_77),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_59),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_127),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_26),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_13),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_53),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_81),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_28),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_10),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_108),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_72),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_35),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_35),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_13),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_40),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_7),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_73),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_60),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_8),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_116),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_69),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_58),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_18),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_48),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_18),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_90),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_12),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_3),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_135),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_99),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_67),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_78),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_40),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_42),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_38),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_130),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_79),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_113),
.Y(n_211)
);

BUFx2_ASAP7_75t_SL g212 ( 
.A(n_9),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_86),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_101),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_17),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_76),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_10),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_37),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_37),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_45),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_26),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_65),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_47),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_46),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_22),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_32),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_83),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_54),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_43),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_3),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_94),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_1),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_0),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_21),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_22),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_100),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_109),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_97),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_85),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_32),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_47),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_89),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_133),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_98),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_20),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_15),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_44),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_57),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_129),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_51),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_16),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_15),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_24),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_46),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_50),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_55),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_111),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_42),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_56),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_33),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_61),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_80),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_145),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_27),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_5),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_52),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_2),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_39),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_68),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_92),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_1),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_75),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_93),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_33),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_95),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_96),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_82),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_120),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_125),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_25),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_7),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_122),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_104),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_74),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_64),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_14),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_63),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_110),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_138),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_146),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_21),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_38),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_161),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_182),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

INVxp33_ASAP7_75t_SL g310 ( 
.A(n_156),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_242),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_232),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_156),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_180),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_265),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_153),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_215),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_217),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_164),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_215),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_209),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_153),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_215),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_183),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_215),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_217),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_215),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_175),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_158),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_218),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_184),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_218),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_185),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_248),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_186),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_187),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_188),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_190),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_191),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_218),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_195),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_218),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_218),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_198),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_229),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_229),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_199),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_200),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_240),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_203),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_229),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_229),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_174),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_240),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_240),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_171),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_204),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_158),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_171),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_283),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_205),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_168),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_281),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_211),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_178),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_320),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_310),
.B(n_213),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_213),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_303),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_323),
.B(n_168),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_306),
.A2(n_260),
.B1(n_192),
.B2(n_233),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_281),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_293),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_286),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_286),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_312),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_293),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_202),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_150),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_303),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_319),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_304),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_305),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_327),
.B(n_150),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_329),
.B(n_332),
.Y(n_403)
);

CKINVDCx11_ASAP7_75t_R g404 ( 
.A(n_331),
.Y(n_404)
);

BUFx8_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_202),
.Y(n_407)
);

OAI22x1_ASAP7_75t_SL g408 ( 
.A1(n_334),
.A2(n_290),
.B1(n_196),
.B2(n_302),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_226),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_330),
.B(n_241),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_318),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_305),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_316),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_325),
.B(n_241),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_308),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_308),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_339),
.B(n_313),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_309),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_309),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_330),
.B(n_272),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_315),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_311),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_348),
.B(n_272),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_348),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_307),
.A2(n_291),
.B1(n_302),
.B2(n_315),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_349),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_418),
.B(n_325),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_328),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_338),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_378),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

INVx4_ASAP7_75t_SL g444 ( 
.A(n_398),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g445 ( 
.A1(n_390),
.A2(n_314),
.B(n_311),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

CKINVDCx6p67_ASAP7_75t_R g447 ( 
.A(n_427),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_342),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_314),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_418),
.B(n_344),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_378),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_345),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_404),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_378),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_397),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_375),
.B(n_347),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_398),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_401),
.Y(n_458)
);

BUFx6f_ASAP7_75t_SL g459 ( 
.A(n_418),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_350),
.Y(n_460)
);

AO22x2_ASAP7_75t_L g461 ( 
.A1(n_376),
.A2(n_307),
.B1(n_212),
.B2(n_282),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_419),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_401),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_411),
.B(n_354),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_376),
.A2(n_269),
.B1(n_274),
.B2(n_193),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g469 ( 
.A(n_385),
.B(n_317),
.C(n_352),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_411),
.B(n_357),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_382),
.B(n_369),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_414),
.B(n_364),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_419),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_416),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_432),
.A2(n_221),
.B1(n_223),
.B2(n_291),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_422),
.B(n_368),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_377),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_416),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_394),
.B(n_340),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_422),
.B(n_371),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_385),
.B(n_372),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_424),
.B(n_282),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_421),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_382),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_382),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_380),
.B(n_333),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_416),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_404),
.Y(n_495)
);

INVxp33_ASAP7_75t_SL g496 ( 
.A(n_381),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_412),
.A2(n_425),
.B1(n_388),
.B2(n_407),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_429),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_424),
.B(n_353),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_389),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_412),
.A2(n_251),
.B1(n_206),
.B2(n_267),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_405),
.B(n_336),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_432),
.A2(n_208),
.B1(n_179),
.B2(n_181),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_429),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_380),
.B(n_343),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_394),
.B(n_340),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_392),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_417),
.A2(n_355),
.B1(n_238),
.B2(n_225),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_405),
.B(n_341),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_398),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_406),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_377),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_396),
.B(n_358),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_377),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_406),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_377),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_409),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_396),
.B(n_358),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_409),
.Y(n_527)
);

BUFx8_ASAP7_75t_SL g528 ( 
.A(n_389),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_412),
.A2(n_197),
.B1(n_194),
.B2(n_207),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_410),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_394),
.B(n_363),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_399),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_413),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_413),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_388),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_402),
.B(n_359),
.Y(n_539)
);

NOR2x1p5_ASAP7_75t_L g540 ( 
.A(n_425),
.B(n_219),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_400),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_400),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_402),
.A2(n_257),
.B(n_157),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_420),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_405),
.B(n_165),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_388),
.B(n_317),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_407),
.B(n_154),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_426),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_387),
.B(n_400),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_387),
.B(n_155),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_400),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_400),
.Y(n_555)
);

BUFx6f_ASAP7_75t_SL g556 ( 
.A(n_430),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_428),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_405),
.B(n_425),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_431),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_400),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_433),
.Y(n_563)
);

INVx8_ASAP7_75t_L g564 ( 
.A(n_400),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_434),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_434),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_399),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_435),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_400),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_387),
.B(n_360),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_405),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_435),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_436),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_407),
.A2(n_288),
.B1(n_258),
.B2(n_227),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_436),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_423),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_423),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_437),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_430),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_430),
.Y(n_582)
);

AND2x6_ASAP7_75t_SL g583 ( 
.A(n_456),
.B(n_234),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_440),
.B(n_151),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_449),
.B(n_423),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_448),
.B(n_151),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_482),
.B(n_423),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_487),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_498),
.B(n_423),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_508),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_521),
.B(n_526),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_452),
.B(n_460),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_531),
.Y(n_594)
);

BUFx12f_ASAP7_75t_L g595 ( 
.A(n_453),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_L g596 ( 
.A(n_483),
.B(n_214),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_539),
.B(n_423),
.Y(n_597)
);

AND2x2_ASAP7_75t_SL g598 ( 
.A(n_504),
.B(n_153),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_449),
.B(n_423),
.Y(n_599)
);

O2A1O1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_439),
.A2(n_390),
.B(n_301),
.C(n_237),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_449),
.B(n_423),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_509),
.B(n_153),
.Y(n_602)
);

BUFx6f_ASAP7_75t_SL g603 ( 
.A(n_487),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_550),
.A2(n_430),
.B1(n_201),
.B2(n_216),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_531),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_581),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_552),
.B(n_153),
.Y(n_607)
);

OAI22x1_ASAP7_75t_R g608 ( 
.A1(n_453),
.A2(n_236),
.B1(n_224),
.B2(n_220),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_571),
.B(n_553),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_483),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_520),
.B(n_403),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_513),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_520),
.B(n_403),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_480),
.B(n_512),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_513),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_522),
.B(n_162),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_550),
.A2(n_278),
.B1(n_271),
.B2(n_268),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_514),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_514),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_438),
.B(n_381),
.C(n_373),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_548),
.B(n_189),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_450),
.B(n_152),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_522),
.B(n_176),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_480),
.B(n_512),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_517),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_517),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_471),
.B(n_373),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_488),
.B(n_186),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_459),
.A2(n_249),
.B1(n_254),
.B2(n_177),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_572),
.B(n_246),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_477),
.B(n_152),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_488),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_524),
.B(n_264),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_582),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_481),
.B(n_159),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_465),
.B(n_470),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_540),
.Y(n_639)
);

INVxp33_ASAP7_75t_L g640 ( 
.A(n_485),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_547),
.A2(n_300),
.B1(n_297),
.B2(n_256),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_529),
.B(n_159),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_550),
.A2(n_189),
.B1(n_262),
.B2(n_280),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_524),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_537),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_529),
.B(n_160),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_572),
.B(n_160),
.Y(n_647)
);

INVx8_ASAP7_75t_L g648 ( 
.A(n_459),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_472),
.B(n_163),
.Y(n_649)
);

INVx8_ASAP7_75t_L g650 ( 
.A(n_459),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_580),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_525),
.B(n_374),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_550),
.A2(n_222),
.B(n_230),
.C(n_231),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_525),
.B(n_527),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_580),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_515),
.B(n_163),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_537),
.B(n_166),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_537),
.B(n_166),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_540),
.A2(n_167),
.B1(n_279),
.B2(n_284),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_533),
.B(n_374),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_519),
.Y(n_661)
);

NOR2x1p5_ASAP7_75t_SL g662 ( 
.A(n_442),
.B(n_379),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_537),
.B(n_509),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_535),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_510),
.B(n_189),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_478),
.B(n_363),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_374),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_528),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_536),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_559),
.B(n_167),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_478),
.B(n_366),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_510),
.B(n_189),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_538),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_538),
.B(n_170),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_503),
.A2(n_170),
.B1(n_172),
.B2(n_279),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_542),
.B(n_391),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_542),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_546),
.B(n_391),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_505),
.B(n_511),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_505),
.B(n_172),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_502),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_546),
.B(n_391),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_549),
.B(n_561),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_469),
.B(n_549),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_519),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_561),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_563),
.Y(n_688)
);

INVxp33_ASAP7_75t_SL g689 ( 
.A(n_502),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_545),
.A2(n_189),
.B1(n_287),
.B2(n_169),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_563),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_461),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_575),
.B(n_284),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_565),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_545),
.A2(n_165),
.B1(n_169),
.B2(n_173),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_565),
.B(n_285),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_566),
.A2(n_299),
.B1(n_289),
.B2(n_292),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_566),
.B(n_285),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_567),
.B(n_391),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_534),
.B(n_239),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_567),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_523),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_574),
.B(n_289),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_492),
.B(n_263),
.C(n_250),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_574),
.B(n_391),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_516),
.B(n_534),
.C(n_532),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_469),
.A2(n_298),
.B1(n_292),
.B2(n_294),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_523),
.B(n_235),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_530),
.B(n_70),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_545),
.B(n_384),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_530),
.B(n_243),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_543),
.B(n_384),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_543),
.B(n_384),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_551),
.B(n_384),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_461),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_557),
.B(n_71),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_557),
.B(n_294),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_558),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_532),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_558),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_560),
.B(n_295),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_467),
.B(n_295),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_560),
.B(n_384),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_476),
.B(n_245),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_569),
.B(n_298),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_569),
.B(n_247),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_573),
.B(n_244),
.Y(n_727)
);

AND2x2_ASAP7_75t_SL g728 ( 
.A(n_476),
.B(n_408),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_556),
.A2(n_299),
.B1(n_255),
.B2(n_259),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_573),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_576),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_461),
.A2(n_483),
.B1(n_578),
.B2(n_576),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_578),
.B(n_457),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_442),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_457),
.B(n_386),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_568),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_445),
.B(n_253),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_445),
.B(n_277),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_474),
.B(n_386),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_568),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_474),
.B(n_386),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_483),
.Y(n_742)
);

NOR2x1p5_ASAP7_75t_L g743 ( 
.A(n_447),
.B(n_252),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_483),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_606),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_593),
.B(n_441),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_614),
.B(n_626),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_592),
.B(n_443),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_609),
.B(n_496),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_617),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_636),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_590),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_584),
.B(n_455),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_588),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_584),
.B(n_455),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_638),
.B(n_474),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_590),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_591),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_586),
.B(n_462),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_621),
.B(n_408),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_680),
.B(n_447),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_591),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_612),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_589),
.A2(n_564),
.B(n_577),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_648),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_586),
.B(n_462),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_633),
.A2(n_556),
.B1(n_483),
.B2(n_461),
.Y(n_767)
);

BUFx4f_ASAP7_75t_L g768 ( 
.A(n_648),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_634),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_648),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_663),
.B(n_464),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_650),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_650),
.B(n_595),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_692),
.A2(n_715),
.B1(n_685),
.B2(n_594),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_640),
.Y(n_775)
);

OR2x2_ASAP7_75t_SL g776 ( 
.A(n_682),
.B(n_495),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_615),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_619),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_619),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_633),
.A2(n_489),
.B1(n_494),
.B2(n_562),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_620),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_650),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_665),
.B(n_670),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_605),
.B(n_489),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_674),
.B(n_464),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_669),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_630),
.B(n_495),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_587),
.A2(n_564),
.B(n_577),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_685),
.Y(n_789)
);

AOI21xp33_ASAP7_75t_L g790 ( 
.A1(n_637),
.A2(n_624),
.B(n_649),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_637),
.A2(n_554),
.B1(n_494),
.B2(n_518),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_620),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_627),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_627),
.Y(n_794)
);

INVxp33_ASAP7_75t_L g795 ( 
.A(n_629),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_624),
.B(n_494),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_736),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_628),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_681),
.B(n_518),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_645),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_SL g801 ( 
.A(n_642),
.B(n_261),
.C(n_273),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_651),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_651),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_655),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_SL g805 ( 
.A(n_649),
.B(n_276),
.C(n_275),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_SL g806 ( 
.A(n_646),
.B(n_266),
.C(n_500),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_610),
.B(n_541),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_595),
.B(n_564),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_SL g809 ( 
.A(n_719),
.B(n_165),
.C(n_169),
.Y(n_809)
);

INVx3_ASAP7_75t_SL g810 ( 
.A(n_740),
.Y(n_810)
);

INVx5_ASAP7_75t_L g811 ( 
.A(n_610),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_661),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_678),
.B(n_473),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_709),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_709),
.B(n_716),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_687),
.B(n_688),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_691),
.B(n_473),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_724),
.A2(n_484),
.B1(n_490),
.B2(n_491),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_686),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_694),
.B(n_484),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_701),
.B(n_490),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_689),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_686),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_732),
.B(n_570),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_700),
.B(n_554),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_702),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_742),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_702),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_742),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_667),
.B(n_173),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_716),
.B(n_555),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_598),
.B(n_555),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_654),
.B(n_499),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_720),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_718),
.Y(n_835)
);

INVx5_ASAP7_75t_L g836 ( 
.A(n_602),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_684),
.B(n_499),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_737),
.A2(n_562),
.B1(n_555),
.B2(n_507),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_744),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_667),
.B(n_287),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_730),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_730),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_656),
.B(n_562),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_720),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_675),
.B(n_703),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_731),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_734),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_SL g848 ( 
.A(n_598),
.B(n_287),
.Y(n_848)
);

O2A1O1Ixp5_ASAP7_75t_L g849 ( 
.A1(n_607),
.A2(n_501),
.B(n_507),
.C(n_451),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_734),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_744),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_737),
.A2(n_501),
.B1(n_577),
.B2(n_486),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_644),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_639),
.B(n_444),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_672),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_672),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_672),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_733),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_632),
.B(n_444),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_675),
.B(n_703),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_599),
.B(n_570),
.Y(n_861)
);

AOI22x1_ASAP7_75t_L g862 ( 
.A1(n_743),
.A2(n_466),
.B1(n_446),
.B2(n_451),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_712),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_717),
.B(n_468),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_717),
.B(n_468),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_738),
.A2(n_579),
.B1(n_486),
.B2(n_497),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_632),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_601),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_708),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_632),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_622),
.B(n_444),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_713),
.Y(n_872)
);

INVx5_ASAP7_75t_L g873 ( 
.A(n_602),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_585),
.B(n_570),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_708),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_608),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_602),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_721),
.B(n_466),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_690),
.A2(n_475),
.B1(n_479),
.B2(n_446),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_721),
.B(n_725),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_585),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_671),
.B(n_579),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_SL g883 ( 
.A(n_603),
.B(n_570),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_603),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_444),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_714),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_696),
.B(n_579),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_725),
.B(n_475),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_641),
.B(n_486),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_706),
.B(n_497),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_597),
.B(n_710),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_611),
.B(n_497),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_613),
.B(n_458),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_728),
.A2(n_458),
.B1(n_454),
.B2(n_506),
.Y(n_894)
);

INVx5_ASAP7_75t_L g895 ( 
.A(n_602),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_664),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_711),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_652),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_618),
.B(n_463),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_659),
.B(n_506),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_604),
.B(n_454),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_711),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_723),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_660),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_698),
.B(n_697),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_668),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_664),
.B(n_493),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_811),
.A2(n_564),
.B(n_596),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_789),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_790),
.B(n_728),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_749),
.A2(n_647),
.B1(n_658),
.B2(n_657),
.Y(n_911)
);

BUFx2_ASAP7_75t_SL g912 ( 
.A(n_786),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_845),
.A2(n_695),
.B(n_676),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_860),
.B(n_631),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_811),
.A2(n_564),
.B(n_739),
.Y(n_915)
);

BUFx2_ASAP7_75t_SL g916 ( 
.A(n_765),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_880),
.A2(n_600),
.B(n_726),
.C(n_727),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_811),
.A2(n_741),
.B(n_735),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_795),
.B(n_583),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_SL g920 ( 
.A1(n_848),
.A2(n_707),
.B1(n_729),
.B2(n_722),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_747),
.B(n_643),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_891),
.A2(n_607),
.B(n_623),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_749),
.A2(n_727),
.B(n_726),
.C(n_653),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_SL g924 ( 
.A(n_760),
.B(n_693),
.C(n_673),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_815),
.A2(n_662),
.B(n_635),
.C(n_616),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_761),
.A2(n_625),
.B1(n_699),
.B2(n_683),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_795),
.B(n_705),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_789),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_805),
.A2(n_666),
.B(n_673),
.C(n_677),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_775),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_746),
.B(n_679),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_SL g932 ( 
.A(n_814),
.B(n_602),
.Y(n_932)
);

OA21x2_ASAP7_75t_L g933 ( 
.A1(n_891),
.A2(n_666),
.B(n_479),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_815),
.B(n_493),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_SL g935 ( 
.A(n_760),
.B(n_0),
.C(n_4),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_800),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_814),
.B(n_544),
.Y(n_937)
);

AO22x1_ASAP7_75t_L g938 ( 
.A1(n_787),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_822),
.B(n_149),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_754),
.B(n_11),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_754),
.B(n_12),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_748),
.B(n_393),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_800),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_847),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_797),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_830),
.B(n_14),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_847),
.Y(n_947)
);

O2A1O1Ixp5_ASAP7_75t_L g948 ( 
.A1(n_796),
.A2(n_393),
.B(n_379),
.C(n_148),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_857),
.B(n_144),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_745),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_850),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_831),
.A2(n_384),
.B(n_142),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_765),
.B(n_139),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_769),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_R g955 ( 
.A(n_768),
.B(n_126),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_831),
.A2(n_119),
.B(n_118),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_761),
.B(n_106),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_840),
.B(n_769),
.Y(n_958)
);

CKINVDCx16_ASAP7_75t_R g959 ( 
.A(n_773),
.Y(n_959)
);

BUFx2_ASAP7_75t_SL g960 ( 
.A(n_770),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_810),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_774),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_892),
.A2(n_102),
.B(n_88),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_800),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_869),
.B(n_23),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_774),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_905),
.B(n_28),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_750),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_800),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_768),
.B(n_29),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_770),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_772),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_875),
.B(n_29),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_751),
.B(n_30),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_850),
.Y(n_975)
);

OAI21xp33_ASAP7_75t_L g976 ( 
.A1(n_783),
.A2(n_31),
.B(n_34),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_892),
.A2(n_31),
.B(n_34),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_816),
.B(n_36),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_810),
.B(n_36),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_L g980 ( 
.A(n_867),
.B(n_39),
.C(n_41),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_R g981 ( 
.A(n_883),
.B(n_49),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_855),
.B(n_43),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_788),
.A2(n_824),
.B(n_893),
.Y(n_983)
);

CKINVDCx8_ASAP7_75t_R g984 ( 
.A(n_773),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_853),
.B(n_44),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_825),
.B(n_49),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_757),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_772),
.B(n_782),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_897),
.B(n_902),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_757),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_782),
.B(n_876),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_881),
.B(n_896),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_870),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_773),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_832),
.A2(n_756),
.B(n_766),
.C(n_753),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_825),
.B(n_755),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_799),
.A2(n_843),
.B(n_887),
.C(n_882),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_752),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_764),
.A2(n_837),
.B(n_833),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_864),
.A2(n_878),
.B(n_865),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_888),
.A2(n_759),
.B(n_861),
.Y(n_1001)
);

NOR2xp67_ASAP7_75t_SL g1002 ( 
.A(n_836),
.B(n_873),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_SL g1003 ( 
.A1(n_889),
.A2(n_874),
.B(n_907),
.C(n_807),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_858),
.B(n_898),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_881),
.B(n_896),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_758),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_763),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_881),
.A2(n_818),
.B1(n_839),
.B2(n_829),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_808),
.B(n_856),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_896),
.B(n_890),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_904),
.B(n_906),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_778),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_868),
.B(n_863),
.Y(n_1013)
);

NAND2x1p5_ASAP7_75t_L g1014 ( 
.A(n_827),
.B(n_829),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_808),
.Y(n_1015)
);

BUFx5_ASAP7_75t_L g1016 ( 
.A(n_854),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_827),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_870),
.B(n_884),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_900),
.A2(n_801),
.B(n_817),
.C(n_785),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_781),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_896),
.B(n_827),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_849),
.A2(n_818),
.B(n_903),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_827),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_890),
.A2(n_799),
.B1(n_871),
.B2(n_887),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_901),
.A2(n_882),
.B(n_866),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_829),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_872),
.B(n_886),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_871),
.A2(n_801),
.B1(n_784),
.B2(n_843),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_894),
.A2(n_767),
.B1(n_839),
.B2(n_829),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_798),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_784),
.B(n_834),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_919),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_945),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_999),
.A2(n_852),
.B(n_907),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_914),
.B(n_820),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_1025),
.A2(n_899),
.B(n_821),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_913),
.A2(n_806),
.B(n_889),
.C(n_885),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_950),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_944),
.Y(n_1039)
);

NOR2xp67_ASAP7_75t_SL g1040 ( 
.A(n_984),
.B(n_912),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_910),
.A2(n_967),
.B(n_965),
.C(n_966),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1004),
.B(n_839),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_908),
.A2(n_819),
.B(n_763),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_996),
.A2(n_894),
.B1(n_839),
.B2(n_851),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_930),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_1023),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_997),
.A2(n_838),
.B(n_791),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1000),
.A2(n_813),
.B(n_771),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1009),
.B(n_808),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1001),
.A2(n_780),
.B(n_879),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_958),
.B(n_776),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_961),
.B(n_851),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_927),
.B(n_834),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_911),
.B(n_851),
.Y(n_1054)
);

INVx8_ASAP7_75t_L g1055 ( 
.A(n_936),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_968),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_954),
.Y(n_1057)
);

AND2x6_ASAP7_75t_L g1058 ( 
.A(n_1017),
.B(n_851),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_936),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_971),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_986),
.A2(n_885),
.B(n_826),
.C(n_803),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_915),
.A2(n_792),
.B(n_777),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_1023),
.B(n_844),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_946),
.B(n_806),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_920),
.B(n_809),
.C(n_862),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_998),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_993),
.Y(n_1067)
);

CKINVDCx8_ASAP7_75t_R g1068 ( 
.A(n_916),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_991),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_925),
.A2(n_779),
.A3(n_846),
.B(n_828),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_931),
.A2(n_895),
.B(n_873),
.Y(n_1071)
);

BUFx4_ASAP7_75t_SL g1072 ( 
.A(n_979),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1011),
.B(n_842),
.Y(n_1073)
);

OAI22x1_ASAP7_75t_L g1074 ( 
.A1(n_1028),
.A2(n_859),
.B1(n_809),
.B2(n_812),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_1017),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_995),
.A2(n_895),
.B(n_836),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_909),
.B(n_762),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_962),
.A2(n_804),
.B(n_793),
.C(n_794),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_989),
.B(n_859),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1027),
.B(n_802),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_928),
.B(n_823),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_1018),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_978),
.B(n_835),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1006),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_1017),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1003),
.A2(n_836),
.B(n_873),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_1021),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_943),
.B(n_841),
.Y(n_1088)
);

AO31x2_ASAP7_75t_L g1089 ( 
.A1(n_1029),
.A2(n_879),
.A3(n_877),
.B(n_873),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1013),
.B(n_854),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_943),
.B(n_877),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1022),
.A2(n_922),
.B(n_917),
.Y(n_1092)
);

AO21x2_ASAP7_75t_L g1093 ( 
.A1(n_1022),
.A2(n_1024),
.B(n_1010),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_923),
.A2(n_924),
.B(n_1019),
.C(n_973),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_1029),
.A2(n_1008),
.A3(n_977),
.B(n_966),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_921),
.B(n_1012),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_962),
.A2(n_1030),
.B1(n_1020),
.B2(n_974),
.Y(n_1097)
);

NOR4xp25_ASAP7_75t_L g1098 ( 
.A(n_976),
.B(n_957),
.C(n_985),
.D(n_929),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1031),
.B(n_982),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_963),
.A2(n_952),
.A3(n_942),
.B(n_934),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_932),
.A2(n_926),
.B(n_992),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1005),
.B(n_941),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_948),
.A2(n_933),
.B(n_947),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_959),
.B(n_1015),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_951),
.B(n_1007),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_1026),
.Y(n_1106)
);

AOI221x1_ASAP7_75t_L g1107 ( 
.A1(n_980),
.A2(n_956),
.B1(n_940),
.B2(n_1009),
.C(n_949),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_SL g1108 ( 
.A1(n_975),
.A2(n_987),
.B(n_990),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_SL g1109 ( 
.A(n_936),
.B(n_964),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_949),
.B(n_972),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_935),
.B(n_953),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_932),
.A2(n_937),
.B(n_1014),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_960),
.B(n_972),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_988),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_939),
.A2(n_953),
.B(n_938),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_971),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1002),
.A2(n_1026),
.B(n_964),
.C(n_969),
.Y(n_1117)
);

BUFx2_ASAP7_75t_SL g1118 ( 
.A(n_971),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1026),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1016),
.B(n_964),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1016),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_969),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1016),
.B(n_969),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_981),
.A2(n_1016),
.A3(n_970),
.B(n_955),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1016),
.A2(n_972),
.B(n_994),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_983),
.A2(n_918),
.B(n_908),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_997),
.A2(n_790),
.B(n_1025),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1004),
.B(n_593),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_983),
.A2(n_918),
.B(n_908),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_944),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_971),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_983),
.A2(n_918),
.B(n_908),
.Y(n_1132)
);

INVx5_ASAP7_75t_L g1133 ( 
.A(n_936),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1004),
.B(n_593),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_945),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_914),
.B(n_593),
.Y(n_1136)
);

NOR2x1_ASAP7_75t_SL g1137 ( 
.A(n_1008),
.B(n_814),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1004),
.B(n_593),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_950),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1009),
.B(n_765),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_997),
.A2(n_790),
.B(n_1025),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_914),
.B(n_593),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_945),
.Y(n_1143)
);

CKINVDCx8_ASAP7_75t_R g1144 ( 
.A(n_912),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_911),
.B(n_790),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_997),
.A2(n_1025),
.A3(n_983),
.B(n_925),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_914),
.B(n_593),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_SL g1148 ( 
.A1(n_962),
.A2(n_790),
.B(n_680),
.C(n_547),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_983),
.A2(n_918),
.B(n_908),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1004),
.B(n_593),
.Y(n_1150)
);

NAND3x1_ASAP7_75t_L g1151 ( 
.A(n_910),
.B(n_476),
.C(n_505),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_914),
.B(n_593),
.Y(n_1152)
);

INVx8_ASAP7_75t_L g1153 ( 
.A(n_1055),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1043),
.A2(n_1062),
.B(n_1126),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1129),
.A2(n_1149),
.B(n_1132),
.Y(n_1155)
);

OAI211xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1145),
.A2(n_1136),
.B(n_1152),
.C(n_1147),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1142),
.A2(n_1127),
.B1(n_1141),
.B2(n_1035),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1064),
.A2(n_1127),
.B1(n_1141),
.B2(n_1111),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1039),
.Y(n_1159)
);

OA21x2_ASAP7_75t_L g1160 ( 
.A1(n_1092),
.A2(n_1034),
.B(n_1103),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1094),
.A2(n_1041),
.B(n_1150),
.C(n_1138),
.Y(n_1161)
);

AOI221x1_ASAP7_75t_L g1162 ( 
.A1(n_1065),
.A2(n_1074),
.B1(n_1037),
.B2(n_1101),
.C(n_1097),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1130),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1148),
.A2(n_1047),
.B(n_1098),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_1057),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1065),
.A2(n_1134),
.B(n_1128),
.C(n_1138),
.Y(n_1166)
);

INVx6_ASAP7_75t_L g1167 ( 
.A(n_1059),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1048),
.A2(n_1036),
.B(n_1050),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1102),
.B(n_1099),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1033),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_1135),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_1054),
.B(n_1125),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1051),
.A2(n_1032),
.B1(n_1115),
.B2(n_1150),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1060),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1128),
.A2(n_1134),
.B(n_1097),
.C(n_1098),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1056),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_1049),
.B(n_1112),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1096),
.B(n_1042),
.Y(n_1178)
);

INVx8_ASAP7_75t_L g1179 ( 
.A(n_1055),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1139),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1137),
.A2(n_1076),
.A3(n_1086),
.B(n_1044),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1050),
.A2(n_1061),
.B(n_1078),
.C(n_1110),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1032),
.A2(n_1115),
.B1(n_1093),
.B2(n_1143),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1096),
.B(n_1042),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1053),
.B(n_1073),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1066),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1083),
.A2(n_1107),
.B(n_1071),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_1045),
.Y(n_1188)
);

AOI21xp33_ASAP7_75t_L g1189 ( 
.A1(n_1151),
.A2(n_1093),
.B(n_1044),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1082),
.B(n_1135),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1067),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1144),
.B(n_1068),
.Y(n_1192)
);

OAI211xp5_ASAP7_75t_L g1193 ( 
.A1(n_1079),
.A2(n_1104),
.B(n_1084),
.C(n_1114),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1040),
.A2(n_1080),
.B1(n_1081),
.B2(n_1140),
.C(n_1087),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1080),
.A2(n_1105),
.B(n_1108),
.Y(n_1195)
);

AND2x6_ASAP7_75t_L g1196 ( 
.A(n_1121),
.B(n_1063),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1077),
.A2(n_1117),
.B1(n_1090),
.B2(n_1113),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1059),
.A2(n_1133),
.B1(n_1118),
.B2(n_1105),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1124),
.B(n_1085),
.Y(n_1199)
);

AO22x2_ASAP7_75t_L g1200 ( 
.A1(n_1095),
.A2(n_1146),
.B1(n_1119),
.B2(n_1122),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_SL g1201 ( 
.A1(n_1109),
.A2(n_1123),
.B(n_1120),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1088),
.A2(n_1046),
.B(n_1091),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1059),
.A2(n_1133),
.B1(n_1116),
.B2(n_1060),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1052),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1069),
.A2(n_1095),
.B1(n_1058),
.B2(n_1124),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1133),
.A2(n_1116),
.B1(n_1131),
.B2(n_1060),
.Y(n_1206)
);

AOI21xp33_ASAP7_75t_L g1207 ( 
.A1(n_1146),
.A2(n_1046),
.B(n_1088),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1058),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1070),
.A2(n_1091),
.B(n_1089),
.Y(n_1209)
);

AOI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1075),
.A2(n_1106),
.B1(n_1131),
.B2(n_1116),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1058),
.A2(n_1100),
.B(n_1075),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1106),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1131),
.A2(n_1055),
.B1(n_1072),
.B2(n_1124),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1136),
.B(n_306),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1043),
.A2(n_1062),
.B(n_1126),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1060),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1145),
.A2(n_790),
.B1(n_910),
.B2(n_680),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1136),
.A2(n_910),
.B1(n_312),
.B2(n_319),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1136),
.A2(n_910),
.B1(n_312),
.B2(n_319),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1092),
.A2(n_1141),
.B(n_1127),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1057),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1136),
.B(n_306),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1043),
.A2(n_1062),
.B(n_1126),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1059),
.B(n_814),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1038),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_L g1226 ( 
.A(n_1045),
.B(n_930),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1135),
.B(n_1033),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1060),
.Y(n_1228)
);

CKINVDCx8_ASAP7_75t_R g1229 ( 
.A(n_1118),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1136),
.B(n_1152),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1136),
.A2(n_1142),
.B1(n_1152),
.B2(n_1147),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1038),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1092),
.A2(n_1141),
.B(n_1127),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1058),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1145),
.A2(n_790),
.B1(n_910),
.B2(n_680),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1127),
.A2(n_1141),
.B(n_1092),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_L g1237 ( 
.A1(n_1136),
.A2(n_790),
.B1(n_1147),
.B2(n_1142),
.C(n_1152),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1136),
.A2(n_910),
.B1(n_312),
.B2(n_319),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1135),
.B(n_1033),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1136),
.A2(n_1147),
.B1(n_1152),
.B2(n_1142),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1145),
.A2(n_790),
.B1(n_910),
.B2(n_680),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1136),
.A2(n_1147),
.B1(n_1152),
.B2(n_1142),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1033),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1102),
.B(n_747),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1059),
.B(n_814),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1069),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1054),
.B(n_1010),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1054),
.B(n_1010),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1136),
.A2(n_1147),
.B1(n_1152),
.B2(n_1142),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1135),
.B(n_1033),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1136),
.A2(n_790),
.B(n_1147),
.C(n_1142),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1057),
.Y(n_1252)
);

AOI21xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1051),
.A2(n_689),
.B(n_810),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1038),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1044),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1102),
.B(n_747),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1217),
.A2(n_1241),
.B1(n_1235),
.B2(n_1231),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1227),
.B(n_1239),
.Y(n_1258)
);

OA22x2_ASAP7_75t_L g1259 ( 
.A1(n_1193),
.A2(n_1213),
.B1(n_1162),
.B2(n_1169),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1231),
.A2(n_1238),
.B1(n_1219),
.B2(n_1218),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1249),
.B(n_1240),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1251),
.A2(n_1161),
.B(n_1166),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1156),
.A2(n_1249),
.B(n_1161),
.C(n_1242),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1250),
.B(n_1171),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1171),
.B(n_1158),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1182),
.A2(n_1175),
.B(n_1245),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1165),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1178),
.B(n_1184),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1156),
.A2(n_1240),
.B(n_1242),
.C(n_1175),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1164),
.A2(n_1230),
.B(n_1190),
.C(n_1189),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1237),
.B(n_1178),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1170),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1236),
.B(n_1220),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1191),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1204),
.A2(n_1173),
.B1(n_1214),
.B2(n_1222),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1184),
.B(n_1185),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1220),
.B(n_1233),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1224),
.A2(n_1203),
.B(n_1198),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1167),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1233),
.B(n_1255),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1168),
.A2(n_1223),
.B(n_1154),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1244),
.B(n_1256),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1157),
.B(n_1165),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1255),
.B(n_1157),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1243),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1199),
.B(n_1189),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1226),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1197),
.A2(n_1253),
.B(n_1193),
.C(n_1221),
.Y(n_1288)
);

AOI211xp5_ASAP7_75t_L g1289 ( 
.A1(n_1194),
.A2(n_1197),
.B(n_1192),
.C(n_1252),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1176),
.B(n_1180),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1252),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1211),
.A2(n_1177),
.B(n_1206),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1177),
.B(n_1172),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1186),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1188),
.A2(n_1247),
.B(n_1248),
.C(n_1172),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1225),
.B(n_1254),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1232),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1159),
.B(n_1163),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1188),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1247),
.Y(n_1300)
);

BUFx4f_ASAP7_75t_SL g1301 ( 
.A(n_1204),
.Y(n_1301)
);

NOR2xp67_ASAP7_75t_L g1302 ( 
.A(n_1246),
.B(n_1212),
.Y(n_1302)
);

O2A1O1Ixp5_ASAP7_75t_L g1303 ( 
.A1(n_1207),
.A2(n_1206),
.B(n_1208),
.C(n_1234),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1229),
.Y(n_1304)
);

AOI31xp33_ASAP7_75t_L g1305 ( 
.A1(n_1205),
.A2(n_1183),
.A3(n_1216),
.B(n_1228),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1205),
.B(n_1187),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1195),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1195),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1248),
.A2(n_1172),
.B(n_1201),
.C(n_1187),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1167),
.A2(n_1234),
.B1(n_1210),
.B2(n_1153),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1202),
.B(n_1209),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1160),
.B(n_1181),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1174),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1153),
.A2(n_1179),
.B1(n_1174),
.B2(n_1196),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1181),
.B(n_1215),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1179),
.A2(n_1155),
.B1(n_1142),
.B2(n_1136),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1217),
.A2(n_910),
.B1(n_728),
.B2(n_496),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1249),
.B(n_1169),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1217),
.A2(n_1136),
.B1(n_1147),
.B2(n_1142),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1200),
.B(n_1236),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1249),
.B(n_1169),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1191),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1200),
.B(n_1236),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1200),
.B(n_1236),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1217),
.A2(n_1136),
.B1(n_1147),
.B2(n_1142),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1249),
.B(n_1169),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1249),
.B(n_1169),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1200),
.B(n_1236),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1227),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1229),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1293),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1307),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1294),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1308),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1261),
.B(n_1284),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1277),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1293),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1273),
.B(n_1280),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1273),
.B(n_1280),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1312),
.A2(n_1315),
.B(n_1320),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1284),
.B(n_1271),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1297),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1320),
.B(n_1323),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1323),
.B(n_1324),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1311),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1324),
.B(n_1328),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1296),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1268),
.B(n_1276),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1328),
.Y(n_1349)
);

AO21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1283),
.A2(n_1327),
.B(n_1321),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1306),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1266),
.A2(n_1262),
.B(n_1309),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1329),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1306),
.B(n_1286),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1286),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1300),
.B(n_1290),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1281),
.B(n_1292),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1303),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1316),
.A2(n_1257),
.B(n_1259),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1266),
.A2(n_1292),
.B(n_1269),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1298),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1265),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1305),
.A2(n_1270),
.B(n_1263),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1334),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1336),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1331),
.B(n_1278),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1343),
.B(n_1264),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1350),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1334),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1345),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1343),
.B(n_1258),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1359),
.A2(n_1260),
.B1(n_1326),
.B2(n_1318),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1338),
.B(n_1339),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1332),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1341),
.B(n_1291),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1352),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1343),
.B(n_1267),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1332),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1355),
.B(n_1325),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1335),
.B(n_1363),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1352),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1339),
.B(n_1346),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1344),
.B(n_1322),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1362),
.B(n_1319),
.Y(n_1384)
);

AOI33xp33_ASAP7_75t_L g1385 ( 
.A1(n_1353),
.A2(n_1289),
.A3(n_1288),
.B1(n_1272),
.B2(n_1295),
.B3(n_1317),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1346),
.B(n_1274),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1362),
.B(n_1299),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1340),
.B(n_1349),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1340),
.B(n_1282),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1333),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1362),
.B(n_1313),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1350),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1340),
.B(n_1285),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1350),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1375),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1365),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1371),
.B(n_1344),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1364),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1371),
.B(n_1344),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1371),
.B(n_1351),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_SL g1401 ( 
.A(n_1385),
.B(n_1363),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1364),
.Y(n_1402)
);

OAI31xp33_ASAP7_75t_L g1403 ( 
.A1(n_1372),
.A2(n_1275),
.A3(n_1358),
.B(n_1357),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1380),
.B(n_1354),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1386),
.B(n_1351),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1372),
.A2(n_1363),
.B1(n_1360),
.B2(n_1352),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1384),
.A2(n_1363),
.B1(n_1360),
.B2(n_1352),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1369),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1367),
.B(n_1354),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1366),
.B(n_1337),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1375),
.B(n_1363),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1385),
.B(n_1352),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1379),
.B(n_1335),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1379),
.A2(n_1353),
.B1(n_1358),
.B2(n_1342),
.C(n_1348),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1384),
.A2(n_1358),
.B1(n_1342),
.B2(n_1348),
.C(n_1347),
.Y(n_1415)
);

OAI33xp33_ASAP7_75t_L g1416 ( 
.A1(n_1387),
.A2(n_1377),
.A3(n_1374),
.B1(n_1378),
.B2(n_1383),
.B3(n_1347),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1391),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1370),
.Y(n_1418)
);

OAI211xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1368),
.A2(n_1392),
.B(n_1394),
.C(n_1287),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1390),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1368),
.B(n_1359),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1390),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1387),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1366),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1388),
.A2(n_1349),
.B1(n_1354),
.B2(n_1356),
.C(n_1361),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1374),
.Y(n_1426)
);

OAI31xp33_ASAP7_75t_L g1427 ( 
.A1(n_1392),
.A2(n_1357),
.A3(n_1310),
.B(n_1361),
.Y(n_1427)
);

INVxp33_ASAP7_75t_SL g1428 ( 
.A(n_1386),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1383),
.B(n_1360),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1366),
.B(n_1337),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1378),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1420),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1422),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1398),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1402),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1396),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1408),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1410),
.B(n_1388),
.Y(n_1438)
);

NOR2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1404),
.B(n_1359),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1411),
.B(n_1413),
.Y(n_1440)
);

INVx4_ASAP7_75t_SL g1441 ( 
.A(n_1424),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1426),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1401),
.B(n_1412),
.C(n_1403),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1431),
.Y(n_1444)
);

NOR2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1424),
.B(n_1304),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1411),
.B(n_1389),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1410),
.B(n_1388),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1418),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1410),
.B(n_1366),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1397),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1401),
.A2(n_1360),
.B(n_1381),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1399),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1405),
.B(n_1382),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1406),
.A2(n_1376),
.B(n_1381),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1430),
.B(n_1366),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1400),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1423),
.Y(n_1457)
);

AND2x6_ASAP7_75t_L g1458 ( 
.A(n_1424),
.B(n_1337),
.Y(n_1458)
);

NOR3xp33_ASAP7_75t_L g1459 ( 
.A(n_1443),
.B(n_1419),
.C(n_1429),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1456),
.B(n_1409),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1456),
.B(n_1395),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1432),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1432),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1441),
.B(n_1438),
.Y(n_1464)
);

OAI21xp33_ASAP7_75t_L g1465 ( 
.A1(n_1443),
.A2(n_1406),
.B(n_1407),
.Y(n_1465)
);

NAND4xp25_ASAP7_75t_SL g1466 ( 
.A(n_1440),
.B(n_1407),
.C(n_1414),
.D(n_1415),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1441),
.B(n_1393),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1440),
.B(n_1413),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1439),
.B(n_1389),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1441),
.B(n_1393),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1458),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1441),
.B(n_1373),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1441),
.B(n_1430),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1433),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1445),
.B(n_1424),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1433),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1434),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1434),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1435),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1457),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1439),
.B(n_1421),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1435),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1458),
.Y(n_1483)
);

AND3x1_ASAP7_75t_SL g1484 ( 
.A(n_1445),
.B(n_1425),
.C(n_1427),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1436),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1450),
.B(n_1377),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1457),
.B(n_1421),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1448),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1458),
.A2(n_1394),
.B1(n_1455),
.B2(n_1449),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1448),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1436),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1458),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1457),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1437),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1468),
.B(n_1465),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1438),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1493),
.B(n_1452),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1478),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1493),
.B(n_1452),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1464),
.B(n_1447),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1481),
.B(n_1446),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1478),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1490),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1473),
.B(n_1447),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1471),
.B(n_1483),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1494),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1466),
.A2(n_1458),
.B1(n_1381),
.B2(n_1376),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1494),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1490),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1471),
.B(n_1449),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1488),
.B(n_1428),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1487),
.B(n_1446),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1459),
.B(n_1417),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1485),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1488),
.B(n_1453),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1480),
.B(n_1453),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1461),
.B(n_1442),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1461),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1462),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1471),
.B(n_1483),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1460),
.B(n_1442),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1463),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1476),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1460),
.B(n_1444),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1505),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1496),
.B(n_1473),
.Y(n_1531)
);

AOI222xp33_ASAP7_75t_L g1532 ( 
.A1(n_1495),
.A2(n_1469),
.B1(n_1416),
.B2(n_1467),
.C1(n_1470),
.C2(n_1475),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1495),
.A2(n_1475),
.B1(n_1451),
.B2(n_1492),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1496),
.B(n_1492),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1520),
.B(n_1477),
.Y(n_1535)
);

NAND2xp33_ASAP7_75t_SL g1536 ( 
.A(n_1515),
.B(n_1475),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1498),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1519),
.B(n_1479),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1498),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1509),
.A2(n_1484),
.B1(n_1489),
.B2(n_1458),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_1482),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_1492),
.Y(n_1542)
);

INVxp67_ASAP7_75t_SL g1543 ( 
.A(n_1513),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1504),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1467),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1504),
.Y(n_1546)
);

INVx4_ASAP7_75t_L g1547 ( 
.A(n_1505),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1517),
.B(n_1486),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1522),
.B(n_1470),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1522),
.B(n_1501),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1508),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1508),
.Y(n_1553)
);

INVx4_ASAP7_75t_L g1554 ( 
.A(n_1511),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1530),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1543),
.B(n_1511),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1530),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1550),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1550),
.Y(n_1559)
);

XNOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1540),
.B(n_1302),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1537),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1537),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1544),
.Y(n_1563)
);

AOI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1544),
.A2(n_1511),
.B(n_1516),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1536),
.B(n_1497),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1500),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1532),
.A2(n_1503),
.B1(n_1451),
.B2(n_1514),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1547),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1551),
.B(n_1499),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1533),
.A2(n_1500),
.B1(n_1506),
.B2(n_1526),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1551),
.B(n_1521),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1531),
.B(n_1547),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1556),
.B(n_1535),
.Y(n_1574)
);

OAI222xp33_ASAP7_75t_L g1575 ( 
.A1(n_1567),
.A2(n_1542),
.B1(n_1534),
.B2(n_1545),
.C1(n_1549),
.C2(n_1554),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1565),
.B(n_1536),
.Y(n_1576)
);

OAI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1567),
.A2(n_1554),
.B1(n_1547),
.B2(n_1535),
.C(n_1553),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1558),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1566),
.B(n_1545),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1571),
.B(n_1518),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1573),
.B(n_1549),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1558),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1573),
.B(n_1554),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1555),
.B(n_1539),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1576),
.A2(n_1570),
.B1(n_1565),
.B2(n_1534),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1577),
.A2(n_1572),
.B1(n_1569),
.B2(n_1560),
.C(n_1559),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_SL g1587 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1578),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1577),
.A2(n_1568),
.B(n_1562),
.Y(n_1589)
);

NOR4xp25_ASAP7_75t_L g1590 ( 
.A(n_1582),
.B(n_1568),
.C(n_1563),
.D(n_1561),
.Y(n_1590)
);

OAI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1574),
.A2(n_1564),
.B(n_1552),
.C(n_1546),
.Y(n_1591)
);

AOI21xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1581),
.A2(n_1542),
.B(n_1541),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1579),
.B(n_1583),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1580),
.B(n_1500),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1583),
.A2(n_1500),
.B1(n_1506),
.B2(n_1542),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1588),
.Y(n_1596)
);

OAI21xp33_ASAP7_75t_L g1597 ( 
.A1(n_1587),
.A2(n_1584),
.B(n_1524),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1593),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1585),
.A2(n_1526),
.B1(n_1506),
.B2(n_1584),
.Y(n_1599)
);

NOR3xp33_ASAP7_75t_L g1600 ( 
.A(n_1586),
.B(n_1541),
.C(n_1538),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1599),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1598),
.Y(n_1602)
);

NAND2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1596),
.B(n_1595),
.Y(n_1603)
);

CKINVDCx14_ASAP7_75t_R g1604 ( 
.A(n_1597),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1600),
.B(n_1594),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1599),
.B(n_1592),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1605),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1603),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1602),
.Y(n_1609)
);

AOI222xp33_ASAP7_75t_L g1610 ( 
.A1(n_1601),
.A2(n_1591),
.B1(n_1590),
.B2(n_1589),
.C1(n_1527),
.C2(n_1525),
.Y(n_1610)
);

AOI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1604),
.A2(n_1528),
.B1(n_1527),
.B2(n_1525),
.C(n_1510),
.Y(n_1611)
);

NOR4xp75_ASAP7_75t_SL g1612 ( 
.A(n_1610),
.B(n_1604),
.C(n_1606),
.D(n_1506),
.Y(n_1612)
);

NAND4xp25_ASAP7_75t_L g1613 ( 
.A(n_1608),
.B(n_1330),
.C(n_1304),
.D(n_1538),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1607),
.B(n_1330),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1613),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1615),
.A2(n_1614),
.B1(n_1609),
.B2(n_1611),
.Y(n_1616)
);

OR3x1_ASAP7_75t_L g1617 ( 
.A(n_1616),
.B(n_1612),
.C(n_1510),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1617),
.B(n_1528),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1618),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1619),
.A2(n_1516),
.B1(n_1512),
.B2(n_1524),
.C(n_1529),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1620),
.A2(n_1516),
.B1(n_1526),
.B2(n_1512),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1621),
.A2(n_1529),
.B1(n_1523),
.B2(n_1502),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1622),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1623),
.A2(n_1491),
.B1(n_1485),
.B2(n_1301),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1314),
.B(n_1454),
.C(n_1279),
.Y(n_1625)
);


endmodule