module fake_jpeg_14883_n_301 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_47),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_22),
.B(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_22),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_53),
.Y(n_96)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_62),
.Y(n_100)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_0),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_68),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_70),
.Y(n_108)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_15),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_30),
.B1(n_39),
.B2(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_84),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_83),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_30),
.B1(n_35),
.B2(n_31),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_19),
.B1(n_38),
.B2(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_23),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_39),
.B1(n_35),
.B2(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_18),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_91),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_18),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_114),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_SL g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_45),
.A2(n_38),
.B1(n_29),
.B2(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_97),
.A2(n_111),
.B1(n_4),
.B2(n_85),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_40),
.B(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_113),
.Y(n_136)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_42),
.A2(n_71),
.B1(n_23),
.B2(n_17),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_67),
.B1(n_15),
.B2(n_36),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_25),
.Y(n_110)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_54),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_20),
.Y(n_112)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_19),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_14),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_48),
.B(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_125),
.B1(n_147),
.B2(n_148),
.Y(n_166)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_49),
.A3(n_43),
.B1(n_62),
.B2(n_60),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_127),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_130),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_73),
.B(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_160),
.Y(n_163)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_37),
.B1(n_15),
.B2(n_44),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_145),
.B1(n_152),
.B2(n_161),
.Y(n_169)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_73),
.A2(n_44),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_135),
.A2(n_146),
.B1(n_156),
.B2(n_157),
.Y(n_193)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

CKINVDCx6p67_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_37),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_37),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_95),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_155),
.C(n_143),
.Y(n_181)
);

OAI22x1_ASAP7_75t_R g144 ( 
.A1(n_104),
.A2(n_62),
.B1(n_1),
.B2(n_3),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_114),
.B(n_116),
.C(n_135),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_88),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_85),
.A2(n_3),
.B1(n_4),
.B2(n_105),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_107),
.B1(n_81),
.B2(n_79),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_156),
.Y(n_185)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_92),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_76),
.A2(n_89),
.B1(n_102),
.B2(n_80),
.Y(n_152)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_119),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_94),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_126),
.Y(n_178)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_100),
.A2(n_89),
.B(n_94),
.C(n_99),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_81),
.A2(n_115),
.B1(n_107),
.B2(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_115),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_182),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_99),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_167),
.A2(n_172),
.B(n_164),
.Y(n_212)
);

NAND2x1_ASAP7_75t_SL g216 ( 
.A(n_170),
.B(n_190),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_127),
.B(n_133),
.C(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_136),
.B(n_154),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_173),
.B(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_121),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_121),
.B(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_139),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_120),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_187),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_175),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_125),
.B1(n_145),
.B2(n_122),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_193),
.B1(n_169),
.B2(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_152),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_148),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_131),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_128),
.B(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_198),
.B(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_188),
.A2(n_189),
.B1(n_187),
.B2(n_169),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_212),
.B1(n_213),
.B2(n_224),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_172),
.A2(n_166),
.B1(n_170),
.B2(n_167),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_221),
.B(n_168),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_176),
.B(n_174),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_179),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_171),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_170),
.B(n_171),
.C(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_170),
.A2(n_167),
.B1(n_181),
.B2(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_183),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_170),
.C(n_182),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_238),
.C(n_199),
.Y(n_253)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_206),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_243),
.B(n_206),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_168),
.C(n_165),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_207),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_221),
.B1(n_205),
.B2(n_208),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_203),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_221),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_221),
.B1(n_216),
.B2(n_202),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_260),
.B1(n_264),
.B2(n_240),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_224),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_253),
.C(n_254),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_246),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_261),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_199),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_219),
.C(n_209),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_257),
.C(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_214),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_221),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_234),
.A2(n_229),
.B1(n_235),
.B2(n_226),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_232),
.B1(n_228),
.B2(n_229),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_235),
.B1(n_225),
.B2(n_239),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_227),
.B(n_242),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_240),
.B1(n_236),
.B2(n_231),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_265),
.B1(n_271),
.B2(n_276),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_247),
.B(n_250),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_256),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_254),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_270),
.Y(n_286)
);

XOR2x2_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_253),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_281),
.B(n_282),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_249),
.B(n_255),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_275),
.B(n_267),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_278),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_272),
.B(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_291),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.C(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_290),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_296),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_297),
.Y(n_301)
);


endmodule