module real_jpeg_5436_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVxp33_ASAP7_75t_L g510 ( 
.A(n_0),
.Y(n_510)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_1),
.A2(n_51),
.B1(n_147),
.B2(n_247),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_1),
.A2(n_51),
.B1(n_289),
.B2(n_298),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_1),
.A2(n_51),
.B1(n_67),
.B2(n_436),
.Y(n_435)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_2),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_2),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_2),
.Y(n_330)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_2),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_2),
.Y(n_453)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_3),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g411 ( 
.A(n_3),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_3),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_138),
.B1(n_165),
.B2(n_169),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_4),
.A2(n_138),
.B1(n_195),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_5),
.A2(n_209),
.B1(n_210),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_5),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_5),
.A2(n_252),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_5),
.A2(n_252),
.B1(n_265),
.B2(n_342),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_5),
.A2(n_252),
.B1(n_431),
.B2(n_433),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_6),
.A2(n_265),
.B1(n_266),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_6),
.B(n_278),
.C(n_281),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_6),
.B(n_115),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_6),
.B(n_235),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_6),
.B(n_91),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_6),
.B(n_348),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_7),
.A2(n_34),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_7),
.A2(n_61),
.B1(n_113),
.B2(n_176),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_7),
.A2(n_61),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_7),
.A2(n_61),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_8),
.A2(n_265),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_8),
.A2(n_288),
.B1(n_296),
.B2(n_303),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_8),
.A2(n_303),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_8),
.A2(n_303),
.B1(n_457),
.B2(n_459),
.Y(n_456)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_10),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_13),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_13),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_14),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_14),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_14),
.A2(n_97),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_97),
.B1(n_190),
.B2(n_194),
.Y(n_189)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_16),
.A2(n_122),
.B1(n_127),
.B2(n_128),
.Y(n_121)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_16),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_16),
.A2(n_127),
.B1(n_151),
.B2(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_16),
.A2(n_127),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_16),
.A2(n_127),
.B1(n_296),
.B2(n_417),
.Y(n_416)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_18),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_18),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_18),
.A2(n_95),
.B1(n_208),
.B2(n_272),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_18),
.A2(n_208),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_18),
.A2(n_208),
.B1(n_353),
.B2(n_355),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_505),
.B(n_508),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_215),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_214),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_158),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_24),
.B(n_158),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_139),
.B2(n_140),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_62),
.C(n_98),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_27),
.A2(n_141),
.B1(n_142),
.B2(n_157),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_27),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_27),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_28),
.A2(n_56),
.B1(n_58),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_28),
.A2(n_251),
.B(n_253),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_28),
.A2(n_39),
.B1(n_251),
.B2(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_29),
.B(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_29),
.A2(n_425),
.B(n_427),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_39),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_34),
.A2(n_404),
.A3(n_405),
.B1(n_406),
.B2(n_408),
.Y(n_403)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_37),
.Y(n_405)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_38),
.Y(n_407)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_39),
.B(n_269),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_39)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_41),
.Y(n_432)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_42),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_43),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_43),
.Y(n_404)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_44),
.Y(n_132)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_44),
.Y(n_177)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g363 ( 
.A(n_46),
.Y(n_363)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_50),
.B(n_57),
.Y(n_205)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_56),
.A2(n_206),
.B(n_456),
.Y(n_475)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_57),
.B(n_207),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_59),
.Y(n_213)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_59),
.Y(n_460)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_60),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_62),
.A2(n_63),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_62),
.A2(n_63),
.B1(n_98),
.B2(n_99),
.Y(n_160)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_90),
.B(n_92),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_64),
.A2(n_264),
.B(n_270),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_64),
.A2(n_90),
.B1(n_302),
.B2(n_341),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_64),
.A2(n_270),
.B(n_341),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_64),
.A2(n_90),
.B1(n_435),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_65),
.A2(n_91),
.B1(n_164),
.B2(n_171),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_65),
.A2(n_91),
.B1(n_164),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_65),
.A2(n_91),
.B1(n_199),
.B2(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_65),
.B(n_271),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_80),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_73),
.B2(n_77),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_69),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_69),
.Y(n_265)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_69),
.Y(n_274)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_79),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_79),
.Y(n_436)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_80),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_82),
.Y(n_280)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_85),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_86),
.Y(n_197)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g391 ( 
.A(n_88),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_90),
.A2(n_305),
.B(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_91),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_92),
.Y(n_171)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_93),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_120),
.B1(n_133),
.B2(n_134),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_133),
.B1(n_134),
.B2(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_100),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_100),
.A2(n_133),
.B1(n_175),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_100),
.A2(n_133),
.B1(n_376),
.B2(n_430),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_107),
.B1(n_108),
.B2(n_112),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_112),
.B(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g345 ( 
.A1(n_113),
.A2(n_269),
.B(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_114),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_115),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_115),
.A2(n_121),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22x1_ASAP7_75t_L g461 ( 
.A1(n_115),
.A2(n_173),
.B1(n_383),
.B2(n_462),
.Y(n_461)
);

AOI32xp33_ASAP7_75t_L g362 ( 
.A1(n_118),
.A2(n_265),
.A3(n_347),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_119),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_132),
.Y(n_350)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_132),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_133),
.B(n_352),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_133),
.A2(n_376),
.B(n_382),
.Y(n_375)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_178),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_159),
.B(n_162),
.CI(n_178),
.CON(n_217),
.SN(n_217)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_162),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_172),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_168),
.Y(n_268)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_173),
.A2(n_345),
.B(n_351),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_173),
.B(n_383),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_173),
.A2(n_351),
.B(n_478),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_177),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B(n_204),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_198),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_180),
.A2(n_204),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_180),
.A2(n_198),
.B1(n_223),
.B2(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_188),
.B(n_189),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_181),
.A2(n_189),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_181),
.A2(n_287),
.B(n_293),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_181),
.A2(n_269),
.B(n_293),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_181),
.A2(n_361),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_182),
.B(n_295),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_182),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_182),
.A2(n_360),
.B1(n_387),
.B2(n_392),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_182),
.A2(n_416),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_193),
.Y(n_418)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_194),
.Y(n_288)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_197),
.Y(n_284)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_197),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_198),
.Y(n_445)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_203),
.Y(n_304)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_254),
.B(n_504),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_217),
.B(n_218),
.Y(n_504)
);

BUFx24_ASAP7_75t_SL g511 ( 
.A(n_217),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.C(n_227),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_224),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_227),
.B(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_245),
.C(n_250),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_228),
.B(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_229),
.B(n_236),
.Y(n_472)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_230),
.Y(n_451)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_237),
.Y(n_449)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_245),
.B(n_250),
.Y(n_443)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_246),
.Y(n_462)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g354 ( 
.A(n_249),
.Y(n_354)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_253),
.Y(n_427)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI311xp33_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_439),
.A3(n_480),
.B1(n_498),
.C1(n_499),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_397),
.B(n_438),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_367),
.B(n_396),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_335),
.B(n_366),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_308),
.B(n_334),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_285),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_262),
.B(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_275),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_263),
.A2(n_275),
.B1(n_276),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_269),
.B(n_409),
.Y(n_408)
);

OAI21xp33_ASAP7_75t_SL g425 ( 
.A1(n_269),
.A2(n_408),
.B(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_299),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_300),
.C(n_307),
.Y(n_336)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_298),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_306),
.B2(n_307),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp33_ASAP7_75t_SL g364 ( 
.A(n_304),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_325),
.B(n_333),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_318),
.B(n_324),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_317),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_323),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B(n_322),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_359),
.B(n_361),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_331),
.Y(n_333)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_329),
.Y(n_361)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_337),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_357),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_343),
.B2(n_344),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_343),
.C(n_357),
.Y(n_368)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_362),
.Y(n_373)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_368),
.B(n_369),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_374),
.B2(n_395),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_373),
.C(n_395),
.Y(n_398)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_384),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_385),
.C(n_386),
.Y(n_419)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_377),
.Y(n_433)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_398),
.B(n_399),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_422),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_400)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_412),
.B2(n_413),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_403),
.B(n_412),
.Y(n_476)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_419),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_419),
.B(n_420),
.C(n_422),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_428),
.B2(n_437),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_423),
.B(n_429),
.C(n_434),
.Y(n_489)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_434),
.Y(n_428)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_430),
.Y(n_478)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_466),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_SL g499 ( 
.A1(n_440),
.A2(n_466),
.B(n_500),
.C(n_503),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_463),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_463),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.C(n_446),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_442),
.B(n_444),
.CI(n_446),
.CON(n_479),
.SN(n_479)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_454),
.C(n_461),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_450),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_450),
.Y(n_488)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_454),
.A2(n_455),
.B1(n_461),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_461),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_479),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_467),
.B(n_479),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_472),
.C(n_473),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_468),
.A2(n_469),
.B1(n_472),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.C(n_477),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_474),
.A2(n_475),
.B1(n_477),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_477),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_479),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_493),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_482),
.A2(n_501),
.B(n_502),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_490),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_490),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.C(n_489),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_496),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_487),
.A2(n_488),
.B1(n_489),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_489),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_495),
.Y(n_501)
);

BUFx4f_ASAP7_75t_SL g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_506),
.Y(n_509)
);

INVx13_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_510),
.Y(n_508)
);


endmodule