module fake_netlist_6_1755_n_49 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_11, n_8, n_10, n_49);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_49;

wire n_41;
wire n_16;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_21;
wire n_18;
wire n_24;
wire n_37;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_38;
wire n_39;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_13;
wire n_35;
wire n_28;
wire n_23;
wire n_17;
wire n_12;
wire n_20;
wire n_30;
wire n_43;
wire n_19;
wire n_47;
wire n_48;
wire n_29;
wire n_31;
wire n_25;
wire n_40;
wire n_44;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_19),
.B1(n_14),
.B2(n_21),
.Y(n_25)
);

AND2x6_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_9),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_1),
.B1(n_3),
.B2(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_15),
.Y(n_30)
);

OAI21x1_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_20),
.B(n_18),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

OAI21x1_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_13),
.B(n_15),
.Y(n_34)
);

OA21x2_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_24),
.B(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_32),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_33),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_43),
.C(n_37),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_46),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_35),
.B(n_38),
.Y(n_49)
);


endmodule