module real_aes_6418_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_713;
wire n_728;
wire n_598;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_762;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_0), .B(n_112), .C(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g459 ( .A(n_0), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_1), .A2(n_138), .B(n_142), .C(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_2), .A2(n_172), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g516 ( .A(n_3), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_4), .B(n_239), .Y(n_258) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_5), .A2(n_172), .B(n_482), .Y(n_481) );
AND2x6_ASAP7_75t_L g138 ( .A(n_6), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g213 ( .A(n_7), .Y(n_213) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_8), .B(n_41), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_9), .A2(n_171), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_10), .B(n_150), .Y(n_225) );
INVx1_ASAP7_75t_L g486 ( .A(n_11), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_12), .B(n_253), .Y(n_541) );
INVx1_ASAP7_75t_L g158 ( .A(n_13), .Y(n_158) );
INVx1_ASAP7_75t_L g553 ( .A(n_14), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_15), .A2(n_148), .B(n_235), .C(n_237), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_16), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_17), .B(n_504), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_18), .B(n_172), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_19), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_20), .A2(n_253), .B(n_268), .C(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_21), .B(n_239), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_22), .B(n_150), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_23), .A2(n_180), .B(n_237), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_24), .B(n_150), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_25), .Y(n_189) );
INVx1_ASAP7_75t_L g146 ( .A(n_26), .Y(n_146) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_28), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_29), .B(n_150), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_30), .A2(n_31), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_30), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_31), .Y(n_751) );
INVx1_ASAP7_75t_L g178 ( .A(n_32), .Y(n_178) );
INVx1_ASAP7_75t_L g495 ( .A(n_33), .Y(n_495) );
INVx2_ASAP7_75t_L g136 ( .A(n_34), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_35), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_36), .A2(n_253), .B(n_254), .C(n_256), .Y(n_252) );
INVxp67_ASAP7_75t_L g179 ( .A(n_37), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_38), .A2(n_142), .B(n_145), .C(n_153), .Y(n_141) );
CKINVDCx14_ASAP7_75t_R g251 ( .A(n_39), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_40), .A2(n_138), .B(n_142), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_41), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g494 ( .A(n_42), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_43), .A2(n_197), .B(n_211), .C(n_212), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_44), .B(n_150), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_45), .A2(n_749), .B1(n_750), .B2(n_753), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_45), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_46), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_47), .Y(n_174) );
INVx1_ASAP7_75t_L g266 ( .A(n_48), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_49), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_50), .B(n_172), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_51), .B(n_462), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_52), .A2(n_142), .B1(n_270), .B2(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_53), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_54), .Y(n_513) );
CKINVDCx14_ASAP7_75t_R g209 ( .A(n_55), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_56), .A2(n_211), .B(n_256), .C(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_57), .Y(n_569) );
INVx1_ASAP7_75t_L g483 ( .A(n_58), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_59), .A2(n_88), .B1(n_452), .B2(n_453), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_59), .Y(n_453) );
INVx1_ASAP7_75t_L g139 ( .A(n_60), .Y(n_139) );
INVx1_ASAP7_75t_L g157 ( .A(n_61), .Y(n_157) );
INVx1_ASAP7_75t_SL g255 ( .A(n_62), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_63), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_64), .B(n_239), .Y(n_272) );
INVx1_ASAP7_75t_L g192 ( .A(n_65), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_SL g503 ( .A1(n_66), .A2(n_256), .B(n_504), .C(n_505), .Y(n_503) );
INVxp67_ASAP7_75t_L g506 ( .A(n_67), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_68), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_68), .Y(n_123) );
INVx1_ASAP7_75t_L g115 ( .A(n_69), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_70), .A2(n_172), .B(n_208), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_71), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_72), .A2(n_172), .B(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_73), .Y(n_498) );
INVx1_ASAP7_75t_L g563 ( .A(n_74), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_75), .A2(n_171), .B(n_173), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_76), .Y(n_140) );
INVx1_ASAP7_75t_L g233 ( .A(n_77), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_78), .A2(n_138), .B(n_142), .C(n_565), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_79), .A2(n_172), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g236 ( .A(n_80), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_81), .B(n_147), .Y(n_529) );
INVx2_ASAP7_75t_L g155 ( .A(n_82), .Y(n_155) );
INVx1_ASAP7_75t_L g224 ( .A(n_83), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_84), .B(n_504), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_85), .A2(n_138), .B(n_142), .C(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g112 ( .A(n_86), .Y(n_112) );
OR2x2_ASAP7_75t_L g456 ( .A(n_86), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g469 ( .A(n_86), .B(n_458), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_87), .A2(n_142), .B(n_191), .C(n_199), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_88), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_89), .B(n_154), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_90), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_91), .A2(n_138), .B(n_142), .C(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_92), .Y(n_545) );
INVx1_ASAP7_75t_L g502 ( .A(n_93), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_94), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_95), .B(n_147), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_96), .B(n_162), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_97), .B(n_162), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_98), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g269 ( .A(n_99), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_100), .A2(n_172), .B(n_501), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_101), .A2(n_466), .B1(n_747), .B2(n_748), .C1(n_754), .C2(n_757), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_102), .A2(n_104), .B1(n_116), .B2(n_762), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g762 ( .A(n_106), .Y(n_762) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g472 ( .A(n_112), .B(n_458), .Y(n_472) );
NOR2x2_ASAP7_75t_L g759 ( .A(n_112), .B(n_457), .Y(n_759) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_464), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g761 ( .A(n_119), .Y(n_761) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_454), .B(n_461), .Y(n_121) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
XOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_451), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_126), .A2(n_467), .B1(n_470), .B2(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g755 ( .A(n_126), .Y(n_755) );
OR4x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_341), .C(n_388), .D(n_428), .Y(n_126) );
NAND3xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_287), .C(n_316), .Y(n_127) );
AOI211xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_202), .B(n_240), .C(n_280), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_129), .A2(n_300), .B(n_317), .C(n_321), .Y(n_316) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_164), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_131), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_SL g283 ( .A(n_131), .Y(n_283) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_131), .Y(n_295) );
AND2x4_ASAP7_75t_L g299 ( .A(n_131), .B(n_247), .Y(n_299) );
AND2x2_ASAP7_75t_L g310 ( .A(n_131), .B(n_187), .Y(n_310) );
OR2x2_ASAP7_75t_L g334 ( .A(n_131), .B(n_243), .Y(n_334) );
AND2x2_ASAP7_75t_L g347 ( .A(n_131), .B(n_248), .Y(n_347) );
AND2x2_ASAP7_75t_L g387 ( .A(n_131), .B(n_373), .Y(n_387) );
AND2x2_ASAP7_75t_L g394 ( .A(n_131), .B(n_357), .Y(n_394) );
AND2x2_ASAP7_75t_L g424 ( .A(n_131), .B(n_165), .Y(n_424) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_159), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_141), .C(n_154), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_133), .A2(n_189), .B(n_190), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_133), .A2(n_221), .B(n_222), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_133), .A2(n_182), .B1(n_492), .B2(n_496), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_133), .A2(n_513), .B(n_514), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_133), .A2(n_563), .B(n_564), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
AND2x4_ASAP7_75t_L g172 ( .A(n_134), .B(n_138), .Y(n_172) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g152 ( .A(n_135), .Y(n_152) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
INVx1_ASAP7_75t_L g271 ( .A(n_136), .Y(n_271) );
INVx1_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
INVx3_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
INVx1_ASAP7_75t_L g504 ( .A(n_137), .Y(n_504) );
BUFx3_ASAP7_75t_L g153 ( .A(n_138), .Y(n_153) );
INVx4_ASAP7_75t_SL g182 ( .A(n_138), .Y(n_182) );
INVx5_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_143), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_149), .C(n_151), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_147), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_147), .A2(n_516), .B(n_517), .C(n_518), .Y(n_515) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_148), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_148), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_148), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
INVx4_ASAP7_75t_L g253 ( .A(n_150), .Y(n_253) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_152), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_154), .A2(n_207), .B(n_214), .Y(n_206) );
INVx1_ASAP7_75t_L g219 ( .A(n_154), .Y(n_219) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_154), .A2(n_548), .B(n_554), .Y(n_547) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_L g163 ( .A(n_155), .B(n_156), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_161), .A2(n_188), .B(n_200), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_161), .B(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
NOR2xp33_ASAP7_75t_SL g531 ( .A(n_161), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_162), .Y(n_230) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_162), .A2(n_500), .B(n_507), .Y(n_499) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_164), .B(n_351), .Y(n_363) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_186), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_165), .B(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g301 ( .A(n_165), .B(n_186), .Y(n_301) );
BUFx3_ASAP7_75t_L g309 ( .A(n_165), .Y(n_309) );
OR2x2_ASAP7_75t_L g330 ( .A(n_165), .B(n_205), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_165), .B(n_351), .Y(n_441) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_170), .B(n_183), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_167), .A2(n_244), .B(n_245), .Y(n_243) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_167), .A2(n_562), .B(n_568), .Y(n_561) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_168), .A2(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_169), .A2(n_491), .B(n_497), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_169), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_169), .A2(n_512), .B(n_519), .Y(n_511) );
INVx1_ASAP7_75t_L g244 ( .A(n_170), .Y(n_244) );
BUFx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_182), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g208 ( .A1(n_175), .A2(n_182), .B(n_209), .C(n_210), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_175), .A2(n_182), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_175), .A2(n_182), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_175), .A2(n_182), .B(n_266), .C(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_175), .A2(n_182), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_175), .A2(n_182), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_175), .A2(n_182), .B(n_550), .C(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_180), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_180), .B(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_180), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g194 ( .A(n_181), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_181), .A2(n_194), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g199 ( .A(n_182), .Y(n_199) );
INVx1_ASAP7_75t_L g245 ( .A(n_183), .Y(n_245) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_185), .B(n_201), .Y(n_200) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_185), .A2(n_537), .B(n_544), .Y(n_536) );
AND2x2_ASAP7_75t_L g246 ( .A(n_186), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g294 ( .A(n_186), .Y(n_294) );
AND2x2_ASAP7_75t_L g357 ( .A(n_186), .B(n_248), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_186), .A2(n_360), .B1(n_362), .B2(n_364), .C(n_365), .Y(n_359) );
AND2x2_ASAP7_75t_L g373 ( .A(n_186), .B(n_243), .Y(n_373) );
AND2x2_ASAP7_75t_L g399 ( .A(n_186), .B(n_283), .Y(n_399) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g279 ( .A(n_187), .B(n_248), .Y(n_279) );
BUFx2_ASAP7_75t_L g413 ( .A(n_187), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .C(n_196), .Y(n_191) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_193), .A2(n_196), .B(n_224), .C(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_196), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_196), .A2(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OAI32xp33_ASAP7_75t_L g379 ( .A1(n_203), .A2(n_340), .A3(n_354), .B1(n_380), .B2(n_381), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_215), .Y(n_203) );
AND2x2_ASAP7_75t_L g320 ( .A(n_204), .B(n_262), .Y(n_320) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g302 ( .A(n_205), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_205), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g374 ( .A(n_205), .B(n_262), .Y(n_374) );
AND2x2_ASAP7_75t_L g385 ( .A(n_205), .B(n_277), .Y(n_385) );
BUFx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g286 ( .A(n_206), .B(n_263), .Y(n_286) );
AND2x2_ASAP7_75t_L g290 ( .A(n_206), .B(n_263), .Y(n_290) );
AND2x2_ASAP7_75t_L g325 ( .A(n_206), .B(n_276), .Y(n_325) );
AND2x2_ASAP7_75t_L g332 ( .A(n_206), .B(n_228), .Y(n_332) );
OAI211xp5_ASAP7_75t_L g337 ( .A1(n_206), .A2(n_283), .B(n_294), .C(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g391 ( .A(n_206), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_206), .B(n_217), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_215), .B(n_274), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_215), .B(n_290), .Y(n_380) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g285 ( .A(n_216), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_228), .Y(n_216) );
AND2x2_ASAP7_75t_L g277 ( .A(n_217), .B(n_229), .Y(n_277) );
OR2x2_ASAP7_75t_L g292 ( .A(n_217), .B(n_229), .Y(n_292) );
AND2x2_ASAP7_75t_L g315 ( .A(n_217), .B(n_276), .Y(n_315) );
INVx1_ASAP7_75t_L g319 ( .A(n_217), .Y(n_319) );
AND2x2_ASAP7_75t_L g338 ( .A(n_217), .B(n_275), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_217), .A2(n_303), .B1(n_349), .B2(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_217), .B(n_391), .Y(n_415) );
AND2x2_ASAP7_75t_L g430 ( .A(n_217), .B(n_290), .Y(n_430) );
INVx4_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx3_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
AND2x2_ASAP7_75t_L g304 ( .A(n_218), .B(n_229), .Y(n_304) );
AND2x2_ASAP7_75t_L g306 ( .A(n_218), .B(n_262), .Y(n_306) );
AND3x2_ASAP7_75t_L g368 ( .A(n_218), .B(n_332), .C(n_369), .Y(n_368) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_219), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_219), .B(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_219), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g403 ( .A(n_228), .B(n_275), .Y(n_403) );
INVx1_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g262 ( .A(n_229), .B(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_229), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_229), .B(n_274), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_229), .B(n_315), .C(n_391), .Y(n_443) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_238), .Y(n_229) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_230), .A2(n_249), .B(n_258), .Y(n_248) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_230), .A2(n_264), .B(n_272), .Y(n_263) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_239), .A2(n_481), .B(n_487), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_259), .B1(n_273), .B2(n_278), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_246), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_243), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g355 ( .A(n_243), .Y(n_355) );
OAI31xp33_ASAP7_75t_L g371 ( .A1(n_246), .A2(n_372), .A3(n_373), .B(n_374), .Y(n_371) );
AND2x2_ASAP7_75t_L g396 ( .A(n_246), .B(n_283), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_246), .B(n_309), .Y(n_442) );
AND2x2_ASAP7_75t_L g351 ( .A(n_247), .B(n_283), .Y(n_351) );
AND2x2_ASAP7_75t_L g412 ( .A(n_247), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g282 ( .A(n_248), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g340 ( .A(n_248), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_253), .B(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_257), .Y(n_542) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_260), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_261), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AOI221x1_ASAP7_75t_SL g328 ( .A1(n_262), .A2(n_329), .B1(n_331), .B2(n_333), .C(n_335), .Y(n_328) );
INVx2_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_263), .Y(n_370) );
INVx2_ASAP7_75t_L g518 ( .A(n_270), .Y(n_518) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g358 ( .A(n_273), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_274), .B(n_291), .Y(n_383) );
INVx1_ASAP7_75t_SL g446 ( .A(n_274), .Y(n_446) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g364 ( .A(n_277), .B(n_290), .Y(n_364) );
INVx1_ASAP7_75t_L g432 ( .A(n_278), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_278), .B(n_361), .Y(n_445) );
INVx2_ASAP7_75t_SL g284 ( .A(n_279), .Y(n_284) );
AND2x2_ASAP7_75t_L g327 ( .A(n_279), .B(n_283), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_279), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_279), .B(n_354), .Y(n_381) );
AOI21xp33_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_284), .B(n_285), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_282), .B(n_354), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_282), .B(n_309), .Y(n_450) );
OR2x2_ASAP7_75t_L g322 ( .A(n_283), .B(n_301), .Y(n_322) );
AND2x2_ASAP7_75t_L g421 ( .A(n_283), .B(n_412), .Y(n_421) );
OAI22xp5_ASAP7_75t_SL g296 ( .A1(n_284), .A2(n_297), .B1(n_302), .B2(n_305), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_284), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g344 ( .A(n_286), .B(n_292), .Y(n_344) );
INVx1_ASAP7_75t_L g408 ( .A(n_286), .Y(n_408) );
AOI311xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_293), .A3(n_295), .B(n_296), .C(n_307), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_291), .A2(n_423), .B1(n_435), .B2(n_438), .C(n_440), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_291), .B(n_446), .Y(n_448) );
INVx2_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g345 ( .A(n_293), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_294), .A2(n_336), .B(n_337), .C(n_339), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_SL g404 ( .A1(n_298), .A2(n_300), .B(n_405), .C(n_406), .Y(n_404) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_299), .B(n_373), .Y(n_439) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_302), .A2(n_322), .B1(n_323), .B2(n_326), .C(n_328), .Y(n_321) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g324 ( .A(n_304), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g407 ( .A(n_304), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_308), .A2(n_366), .B(n_367), .C(n_371), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_309), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_309), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g331 ( .A(n_315), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_319), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g433 ( .A(n_322), .Y(n_433) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_325), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_325), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g437 ( .A(n_325), .Y(n_437) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g378 ( .A(n_327), .B(n_354), .Y(n_378) );
INVx1_ASAP7_75t_SL g372 ( .A(n_334), .Y(n_372) );
INVx1_ASAP7_75t_L g349 ( .A(n_340), .Y(n_349) );
NAND3xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_359), .C(n_375), .Y(n_341) );
AOI322xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .A3(n_346), .B1(n_348), .B2(n_352), .C1(n_356), .C2(n_358), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g395 ( .A1(n_343), .A2(n_396), .B(n_397), .C(n_404), .Y(n_395) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_346), .A2(n_367), .B1(n_398), .B2(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g356 ( .A(n_354), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g393 ( .A(n_354), .B(n_394), .Y(n_393) );
AOI32xp33_ASAP7_75t_L g444 ( .A1(n_354), .A2(n_445), .A3(n_446), .B1(n_447), .B2(n_449), .Y(n_444) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g366 ( .A(n_357), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_357), .A2(n_410), .B1(n_414), .B2(n_416), .C(n_419), .Y(n_409) );
AND2x2_ASAP7_75t_L g423 ( .A(n_357), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g426 ( .A(n_361), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g436 ( .A(n_361), .B(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g427 ( .A(n_370), .B(n_391), .Y(n_427) );
AOI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_379), .C(n_382), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_392), .B(n_395), .C(n_409), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_403), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g418 ( .A(n_415), .Y(n_418) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_425), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI211xp5_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_431), .B(n_434), .C(n_444), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_456), .Y(n_463) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_461), .A2(n_465), .B(n_760), .Y(n_464) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22x1_ASAP7_75t_L g754 ( .A1(n_467), .A2(n_470), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g756 ( .A(n_474), .Y(n_756) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND3x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_669), .C(n_714), .Y(n_475) );
NOR4xp25_ASAP7_75t_L g476 ( .A(n_477), .B(n_592), .C(n_633), .D(n_650), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_508), .B(n_522), .C(n_555), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_479), .B(n_509), .Y(n_508) );
NOR4xp25_ASAP7_75t_L g616 ( .A(n_479), .B(n_610), .C(n_617), .D(n_623), .Y(n_616) );
AND2x2_ASAP7_75t_L g689 ( .A(n_479), .B(n_578), .Y(n_689) );
AND2x2_ASAP7_75t_L g708 ( .A(n_479), .B(n_654), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_479), .B(n_703), .Y(n_717) );
AND2x2_ASAP7_75t_L g730 ( .A(n_479), .B(n_521), .Y(n_730) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g575 ( .A(n_480), .Y(n_575) );
AND2x2_ASAP7_75t_L g582 ( .A(n_480), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g632 ( .A(n_480), .B(n_489), .Y(n_632) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_480), .B(n_578), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_480), .B(n_489), .Y(n_647) );
AND2x2_ASAP7_75t_L g656 ( .A(n_480), .B(n_581), .Y(n_656) );
BUFx2_ASAP7_75t_L g679 ( .A(n_480), .Y(n_679) );
AND2x2_ASAP7_75t_L g683 ( .A(n_480), .B(n_499), .Y(n_683) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_499), .Y(n_488) );
AND2x2_ASAP7_75t_L g521 ( .A(n_489), .B(n_499), .Y(n_521) );
BUFx2_ASAP7_75t_L g585 ( .A(n_489), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_489), .A2(n_618), .B1(n_620), .B2(n_621), .Y(n_617) );
OR2x2_ASAP7_75t_L g639 ( .A(n_489), .B(n_511), .Y(n_639) );
AND2x2_ASAP7_75t_L g703 ( .A(n_489), .B(n_581), .Y(n_703) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g571 ( .A(n_490), .B(n_511), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_490), .B(n_499), .Y(n_578) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_490), .Y(n_620) );
OR2x2_ASAP7_75t_L g655 ( .A(n_490), .B(n_510), .Y(n_655) );
INVx1_ASAP7_75t_L g574 ( .A(n_499), .Y(n_574) );
INVx3_ASAP7_75t_L g583 ( .A(n_499), .Y(n_583) );
BUFx2_ASAP7_75t_L g607 ( .A(n_499), .Y(n_607) );
AND2x2_ASAP7_75t_L g640 ( .A(n_499), .B(n_575), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_508), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_510), .B(n_583), .Y(n_587) );
INVx1_ASAP7_75t_L g615 ( .A(n_510), .Y(n_615) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g581 ( .A(n_511), .Y(n_581) );
INVx1_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
NAND2x1_ASAP7_75t_SL g522 ( .A(n_523), .B(n_533), .Y(n_522) );
AND2x2_ASAP7_75t_L g591 ( .A(n_523), .B(n_546), .Y(n_591) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_523), .Y(n_665) );
AND2x2_ASAP7_75t_L g692 ( .A(n_523), .B(n_612), .Y(n_692) );
AND2x2_ASAP7_75t_L g700 ( .A(n_523), .B(n_662), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_523), .B(n_558), .Y(n_727) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g559 ( .A(n_524), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g576 ( .A(n_524), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g597 ( .A(n_524), .Y(n_597) );
INVx1_ASAP7_75t_L g603 ( .A(n_524), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_524), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g636 ( .A(n_524), .B(n_561), .Y(n_636) );
OR2x2_ASAP7_75t_L g674 ( .A(n_524), .B(n_629), .Y(n_674) );
AOI32xp33_ASAP7_75t_L g686 ( .A1(n_524), .A2(n_687), .A3(n_690), .B1(n_691), .B2(n_692), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_524), .B(n_662), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_524), .B(n_622), .Y(n_737) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g648 ( .A(n_534), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_546), .Y(n_534) );
INVx1_ASAP7_75t_L g610 ( .A(n_535), .Y(n_610) );
AND2x2_ASAP7_75t_L g612 ( .A(n_535), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_535), .B(n_560), .Y(n_629) );
AND2x2_ASAP7_75t_L g662 ( .A(n_535), .B(n_638), .Y(n_662) );
AND2x2_ASAP7_75t_L g699 ( .A(n_535), .B(n_561), .Y(n_699) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g558 ( .A(n_536), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_536), .B(n_560), .Y(n_589) );
AND2x2_ASAP7_75t_L g596 ( .A(n_536), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g637 ( .A(n_536), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_543), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_542), .Y(n_539) );
INVx2_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_546), .B(n_560), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_546), .B(n_604), .Y(n_685) );
INVx1_ASAP7_75t_L g707 ( .A(n_546), .Y(n_707) );
INVx1_ASAP7_75t_L g724 ( .A(n_546), .Y(n_724) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g577 ( .A(n_547), .B(n_560), .Y(n_577) );
AND2x2_ASAP7_75t_L g599 ( .A(n_547), .B(n_561), .Y(n_599) );
INVx1_ASAP7_75t_L g638 ( .A(n_547), .Y(n_638) );
AOI221x1_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_570), .B1(n_576), .B2(n_578), .C(n_579), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_556), .A2(n_643), .B1(n_710), .B2(n_711), .Y(n_709) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
AND2x2_ASAP7_75t_L g601 ( .A(n_557), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g696 ( .A(n_557), .B(n_576), .Y(n_696) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g652 ( .A(n_558), .B(n_577), .Y(n_652) );
INVx1_ASAP7_75t_L g664 ( .A(n_559), .Y(n_664) );
AND2x2_ASAP7_75t_L g675 ( .A(n_559), .B(n_662), .Y(n_675) );
AND2x2_ASAP7_75t_L g742 ( .A(n_559), .B(n_637), .Y(n_742) );
INVx2_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_571), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g694 ( .A(n_571), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_572), .B(n_655), .Y(n_658) );
INVx3_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_573), .A2(n_694), .B(n_739), .Y(n_738) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NOR2xp33_ASAP7_75t_SL g716 ( .A(n_576), .B(n_602), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_577), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g668 ( .A(n_577), .B(n_596), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_577), .B(n_603), .Y(n_745) );
AND2x2_ASAP7_75t_L g614 ( .A(n_578), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g681 ( .A(n_578), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B(n_588), .Y(n_579) );
NAND2x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_581), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g630 ( .A(n_581), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g642 ( .A(n_581), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_581), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g666 ( .A(n_582), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_582), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_582), .B(n_585), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_585), .A2(n_624), .B(n_654), .C(n_656), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_585), .A2(n_672), .B1(n_675), .B2(n_676), .C(n_680), .Y(n_671) );
AND2x2_ASAP7_75t_L g667 ( .A(n_586), .B(n_620), .Y(n_667) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g627 ( .A(n_591), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g698 ( .A(n_591), .B(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_600), .C(n_625), .Y(n_592) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_593), .B(n_712), .C(n_713), .Y(n_711) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
OR2x2_ASAP7_75t_L g684 ( .A(n_595), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_605), .B1(n_608), .B2(n_614), .C(n_616), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_602), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g624 ( .A(n_607), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_607), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
OR2x2_ASAP7_75t_L g744 ( .A(n_607), .B(n_655), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVxp67_ASAP7_75t_L g718 ( .A(n_610), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_612), .B(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_L g619 ( .A(n_613), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_615), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_615), .B(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_615), .B(n_682), .Y(n_721) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_619), .Y(n_645) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g735 ( .A(n_624), .B(n_655), .Y(n_735) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g713 ( .A(n_630), .Y(n_713) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI322xp33_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_639), .A3(n_640), .B1(n_641), .B2(n_644), .C1(n_646), .C2(n_648), .Y(n_633) );
OAI322xp33_ASAP7_75t_L g715 ( .A1(n_634), .A2(n_716), .A3(n_717), .B1(n_718), .B2(n_719), .C1(n_720), .C2(n_722), .Y(n_715) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx4_ASAP7_75t_L g649 ( .A(n_636), .Y(n_649) );
AND2x2_ASAP7_75t_L g710 ( .A(n_636), .B(n_662), .Y(n_710) );
AND2x2_ASAP7_75t_L g723 ( .A(n_636), .B(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_639), .Y(n_734) );
INVx1_ASAP7_75t_L g712 ( .A(n_640), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g646 ( .A(n_642), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g729 ( .A(n_642), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_642), .B(n_683), .Y(n_740) );
OR2x2_ASAP7_75t_L g673 ( .A(n_645), .B(n_674), .Y(n_673) );
INVxp33_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
OAI221xp5_ASAP7_75t_SL g650 ( .A1(n_649), .A2(n_651), .B1(n_653), .B2(n_657), .C(n_659), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g706 ( .A(n_649), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g733 ( .A(n_649), .Y(n_733) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx3_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_656), .A2(n_681), .A3(n_698), .B1(n_700), .B2(n_701), .C1(n_704), .C2(n_708), .Y(n_697) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B1(n_667), .B2(n_668), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_693), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_686), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_674), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
NAND2xp33_ASAP7_75t_SL g691 ( .A(n_677), .B(n_688), .Y(n_691) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
OAI322xp33_ASAP7_75t_L g731 ( .A1(n_679), .A2(n_732), .A3(n_734), .B1(n_735), .B2(n_736), .C1(n_738), .C2(n_741), .Y(n_731) );
AOI21xp33_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_689), .B(n_737), .Y(n_746) );
OAI211xp5_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_695), .B(n_697), .C(n_709), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NOR4xp25_ASAP7_75t_L g714 ( .A(n_715), .B(n_725), .C(n_731), .D(n_743), .Y(n_714) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
CKINVDCx14_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
OAI21xp5_ASAP7_75t_SL g743 ( .A1(n_744), .A2(n_745), .B(n_746), .Y(n_743) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
endmodule