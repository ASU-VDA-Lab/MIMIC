module fake_jpeg_22529_n_280 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_23),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_50),
.B1(n_61),
.B2(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_34),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_53),
.Y(n_72)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_52),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_34),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_65),
.Y(n_96)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_33),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_64),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_25),
.B1(n_32),
.B2(n_17),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_SL g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_68),
.B(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_73),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_26),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_17),
.B1(n_32),
.B2(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_87),
.B1(n_90),
.B2(n_60),
.Y(n_108)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_17),
.B1(n_32),
.B2(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_39),
.B1(n_31),
.B2(n_38),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_97),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_44),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_100),
.B1(n_31),
.B2(n_27),
.Y(n_120)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_33),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_52),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_31),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_0),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_105),
.C(n_128),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_57),
.C(n_58),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_27),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_115),
.B(n_48),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_108),
.A2(n_120),
.B1(n_121),
.B2(n_48),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_57),
.B1(n_56),
.B2(n_18),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_112),
.B1(n_74),
.B2(n_92),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_22),
.B1(n_20),
.B2(n_31),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_0),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

OAI22x1_ASAP7_75t_SL g121 ( 
.A1(n_72),
.A2(n_96),
.B1(n_87),
.B2(n_82),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_27),
.B(n_33),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_71),
.C(n_72),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_132),
.B(n_133),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_134),
.B(n_138),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_146),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_101),
.B1(n_79),
.B2(n_98),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_97),
.B1(n_94),
.B2(n_88),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_147),
.B1(n_156),
.B2(n_158),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_91),
.B1(n_27),
.B2(n_100),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_70),
.B1(n_73),
.B2(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_84),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_100),
.B1(n_27),
.B2(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_84),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_84),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_27),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_157),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_114),
.B(n_102),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_102),
.B(n_1),
.Y(n_157)
);

AO21x2_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_119),
.B(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_163),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_158),
.A2(n_127),
.B1(n_105),
.B2(n_111),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_173),
.B1(n_178),
.B2(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_132),
.B(n_157),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_114),
.B(n_111),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_171),
.B(n_136),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_170),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_112),
.A3(n_123),
.B1(n_104),
.B2(n_119),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_123),
.B(n_117),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_116),
.B1(n_2),
.B2(n_3),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_1),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_180),
.C(n_184),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_4),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_139),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_147),
.B(n_145),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_194),
.B1(n_9),
.B2(n_10),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_176),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_195),
.Y(n_220)
);

AO21x2_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_133),
.B(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_202),
.B(n_203),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_131),
.C(n_148),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_9),
.C(n_10),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_205),
.B(n_174),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_152),
.B(n_7),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_6),
.B(n_8),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_149),
.B(n_110),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_8),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_110),
.C(n_7),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_180),
.C(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_168),
.B1(n_184),
.B2(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_208),
.B(n_162),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_215),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_166),
.A3(n_164),
.B1(n_160),
.B2(n_163),
.C1(n_171),
.C2(n_186),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_213),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_173),
.C(n_176),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_217),
.C(n_224),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_179),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_218),
.B(n_223),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_181),
.C(n_8),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_192),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_188),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_16),
.C(n_10),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_202),
.C(n_201),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_227),
.C(n_207),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_194),
.B(n_204),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_233),
.Y(n_252)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_224),
.Y(n_246)
);

BUFx12_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_194),
.B1(n_188),
.B2(n_202),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_211),
.B1(n_217),
.B2(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_239),
.C(n_214),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_240),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_194),
.C(n_196),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_194),
.B(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_222),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_247),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_248),
.A2(n_230),
.B(n_235),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_213),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_251),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_227),
.B1(n_12),
.B2(n_13),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_259),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_232),
.C(n_229),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_261),
.C(n_228),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_229),
.CI(n_232),
.CON(n_259),
.SN(n_259)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_233),
.B(n_231),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_247),
.C(n_245),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_267),
.B(n_254),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_245),
.B1(n_233),
.B2(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_249),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_258),
.B(n_260),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_269),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_259),
.C(n_9),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_256),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_238),
.A3(n_263),
.B1(n_259),
.B2(n_255),
.C1(n_12),
.C2(n_15),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_275),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_270),
.C(n_14),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_277),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_14),
.Y(n_280)
);


endmodule