module real_jpeg_23825_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_348, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_348;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_1),
.A2(n_26),
.B1(n_57),
.B2(n_58),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_5),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_131),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_131),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_131),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_59),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_7),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_57),
.B1(n_73),
.B2(n_129),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_129),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_129),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_8),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_68),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_8),
.B(n_47),
.C(n_50),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_8),
.B(n_30),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_8),
.A2(n_106),
.B1(n_211),
.B2(n_214),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_58),
.B1(n_66),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_10),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_138),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_138),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_138),
.Y(n_211)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_70),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_42),
.B1(n_75),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_14),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_123)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_15),
.Y(n_117)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_15),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_97),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_84),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_84),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.C(n_80),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_20),
.A2(n_76),
.B1(n_331),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_20),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_44),
.C(n_54),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_24),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_25),
.A2(n_30),
.B(n_38),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_25),
.A2(n_38),
.B(n_83),
.Y(n_275)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_29),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_27),
.A2(n_62),
.B(n_135),
.C(n_155),
.Y(n_154)
);

HAxp5_ASAP7_75t_SL g226 ( 
.A(n_27),
.B(n_134),
.CON(n_226),
.SN(n_226)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_29),
.B(n_58),
.C(n_64),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_29),
.B(n_32),
.C(n_34),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_30),
.A2(n_38),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_30),
.A2(n_38),
.B1(n_171),
.B2(n_226),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_30),
.A2(n_38),
.B1(n_82),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_31),
.A2(n_148),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_31),
.A2(n_37),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_31)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_33),
.A2(n_36),
.B(n_225),
.C(n_227),
.Y(n_224)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_34),
.B(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_38),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_38),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_76),
.C(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_43),
.A2(n_44),
.B1(n_81),
.B2(n_334),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_45),
.A2(n_49),
.B1(n_186),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_45),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_45),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_49),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_123),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_49),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_49),
.B(n_134),
.Y(n_209)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_51),
.B(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_53),
.A2(n_121),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_53),
.B(n_184),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_61),
.B(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_58),
.B(n_134),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_69),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_60),
.A2(n_68),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_60),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_60),
.A2(n_68),
.B1(n_145),
.B2(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_61),
.A2(n_137),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_67),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_68),
.B(n_296),
.Y(n_295)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_76),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_76),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_80),
.B(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_81),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_93),
.B2(n_94),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_90),
.A2(n_143),
.B(n_320),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_328),
.A3(n_340),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_305),
.B(n_327),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_278),
.B(n_304),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_173),
.B(n_259),
.C(n_277),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_157),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_102),
.B(n_157),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_139),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_124),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_104),
.B(n_124),
.C(n_139),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_118),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_105),
.B(n_118),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_110),
.B(n_112),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_106),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_106),
.A2(n_115),
.B1(n_204),
.B2(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_106),
.A2(n_112),
.B(n_193),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_106),
.A2(n_193),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_111),
.B1(n_114),
.B2(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_107),
.B(n_113),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_107),
.A2(n_191),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_109),
.B(n_134),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_117),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_119),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_120),
.B(n_249),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_121),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_121),
.A2(n_184),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_121),
.A2(n_184),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_132),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_127),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_126),
.Y(n_288)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_159),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_149),
.B2(n_156),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_142),
.B(n_146),
.C(n_156),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_143),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_164),
.B(n_166),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_160),
.B(n_162),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.C(n_169),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_166),
.B(n_190),
.Y(n_265)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_169),
.B(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_258),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_253),
.B(n_257),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_237),
.B(n_252),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_220),
.B(n_236),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_200),
.B(n_219),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_187),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_187),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_182),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_195),
.C(n_198),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_207),
.B(n_218),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_206),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_217),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_235),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_235),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_231),
.C(n_232),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_234),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_245),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_247),
.C(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_261),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_276),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_270),
.C(n_276),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_269),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_269),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_268),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_273),
.C(n_275),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_274),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_279),
.B(n_280),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_303),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_290),
.B1(n_301),
.B2(n_302),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_302),
.C(n_303),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_286),
.B2(n_289),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_283),
.A2(n_284),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_283),
.A2(n_315),
.B(n_319),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_297),
.C(n_300),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_292)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_296),
.Y(n_320)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_306),
.B(n_307),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_307)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_312),
.B(n_313),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_313),
.A2(n_330),
.B1(n_335),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_322),
.C(n_326),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_324),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_337),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_337),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.C(n_336),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_341),
.B(n_342),
.Y(n_345)
);


endmodule