module fake_jpeg_28191_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_4),
.B(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_2),
.Y(n_11)
);

BUFx2_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx10_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_1),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_7),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_7),
.A2(n_2),
.B(n_3),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_21),
.B1(n_14),
.B2(n_19),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g21 ( 
.A(n_6),
.B(n_8),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_20),
.A2(n_9),
.B1(n_11),
.B2(n_6),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_21),
.B(n_13),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_11),
.B1(n_13),
.B2(n_4),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_32),
.B(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_33),
.B(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_13),
.B1(n_15),
.B2(n_26),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_35),
.B(n_33),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.C(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_29),
.Y(n_38)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_25),
.B(n_37),
.Y(n_40)
);


endmodule