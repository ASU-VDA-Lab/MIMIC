module fake_jpeg_28941_n_455 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_455);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_21),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_49),
.B(n_51),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_52),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_42),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_61),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_68),
.Y(n_108)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_64),
.Y(n_110)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_77),
.Y(n_111)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_28),
.B(n_8),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_37),
.B(n_8),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_87),
.Y(n_133)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_27),
.B(n_10),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_89),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_37),
.B(n_10),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_35),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_40),
.B1(n_18),
.B2(n_19),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_42),
.B1(n_44),
.B2(n_22),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_100),
.B1(n_113),
.B2(n_117),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_89),
.B1(n_88),
.B2(n_90),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_128),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_32),
.B1(n_44),
.B2(n_22),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_44),
.B1(n_34),
.B2(n_33),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_34),
.B1(n_47),
.B2(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_22),
.B1(n_46),
.B2(n_35),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_78),
.A2(n_32),
.B1(n_22),
.B2(n_16),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_58),
.A2(n_75),
.B1(n_84),
.B2(n_60),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_16),
.B1(n_18),
.B2(n_27),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_132),
.B1(n_138),
.B2(n_142),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_67),
.A2(n_46),
.B1(n_26),
.B2(n_20),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_63),
.B(n_30),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_41),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_56),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_69),
.A2(n_26),
.B1(n_30),
.B2(n_38),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_74),
.A2(n_19),
.B1(n_38),
.B2(n_41),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_41),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_72),
.A2(n_26),
.B1(n_38),
.B2(n_13),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_19),
.B1(n_55),
.B2(n_93),
.Y(n_187)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_147),
.Y(n_233)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_151),
.B(n_155),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_85),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_76),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_161),
.B(n_174),
.Y(n_227)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_116),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_168),
.Y(n_217)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_108),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_179),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_182),
.B(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_102),
.B(n_120),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_81),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_183),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_96),
.A2(n_66),
.B1(n_79),
.B2(n_18),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_178),
.A2(n_188),
.B1(n_110),
.B2(n_107),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_59),
.B1(n_19),
.B2(n_54),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_184),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_117),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_41),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_19),
.B(n_85),
.C(n_50),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_189),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_193),
.B1(n_152),
.B2(n_172),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_96),
.A2(n_18),
.B1(n_50),
.B2(n_11),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_110),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_97),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

OR2x4_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_7),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_141),
.B(n_127),
.C(n_110),
.Y(n_223)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_194),
.A2(n_144),
.B1(n_95),
.B2(n_124),
.Y(n_229)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_151),
.C(n_176),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_196),
.B(n_202),
.C(n_162),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_182),
.C(n_154),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_135),
.B1(n_118),
.B2(n_130),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_219),
.B1(n_171),
.B2(n_195),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_141),
.A3(n_127),
.B1(n_115),
.B2(n_98),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_226),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_154),
.B1(n_106),
.B2(n_153),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_223),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_182),
.B1(n_172),
.B2(n_173),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_130),
.B1(n_135),
.B2(n_140),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_232),
.B1(n_234),
.B2(n_194),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_153),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_173),
.A2(n_140),
.B1(n_114),
.B2(n_137),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_185),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_179),
.A2(n_183),
.B(n_192),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_190),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_154),
.C(n_184),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_239),
.B(n_269),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_250),
.B1(n_251),
.B2(n_259),
.Y(n_278)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_242),
.A2(n_256),
.B1(n_263),
.B2(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_168),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_243),
.B(n_264),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_163),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_245),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_150),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_246),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_219),
.B1(n_210),
.B2(n_214),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_248),
.A2(n_237),
.B(n_211),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_170),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_272),
.C(n_221),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_227),
.A2(n_160),
.B1(n_169),
.B2(n_167),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_254),
.A2(n_213),
.B(n_235),
.Y(n_291)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_225),
.B1(n_208),
.B2(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_212),
.A2(n_157),
.B1(n_149),
.B2(n_180),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_228),
.B1(n_226),
.B2(n_237),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_202),
.A2(n_148),
.B1(n_166),
.B2(n_164),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_271),
.Y(n_309)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_208),
.A2(n_137),
.B1(n_124),
.B2(n_181),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_98),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_208),
.A2(n_125),
.B1(n_112),
.B2(n_147),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_230),
.B(n_196),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_268),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_224),
.A2(n_144),
.B1(n_125),
.B2(n_95),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_270),
.B1(n_201),
.B2(n_204),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_5),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_215),
.B(n_0),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_232),
.A2(n_223),
.B1(n_215),
.B2(n_212),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_221),
.B(n_200),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_207),
.B(n_0),
.C(n_1),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_207),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_273),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_201),
.A2(n_11),
.B(n_14),
.C(n_4),
.D(n_5),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_233),
.B(n_228),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_216),
.A2(n_4),
.B1(n_12),
.B2(n_14),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_275),
.A2(n_231),
.B1(n_233),
.B2(n_198),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_281),
.A2(n_288),
.B(n_298),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_239),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_285),
.A2(n_302),
.B1(n_305),
.B2(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_204),
.C(n_235),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_294),
.C(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_270),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_271),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_293),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_213),
.C(n_218),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_299),
.B1(n_250),
.B2(n_267),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_254),
.A2(n_220),
.B(n_231),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_248),
.A2(n_198),
.B1(n_218),
.B2(n_206),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_240),
.A2(n_197),
.B1(n_206),
.B2(n_220),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_247),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_261),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_262),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_247),
.A2(n_197),
.B1(n_211),
.B2(n_1),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_247),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_1),
.C(n_2),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_311),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_280),
.B(n_293),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_312),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_313),
.A2(n_331),
.B1(n_333),
.B2(n_302),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_273),
.Y(n_314)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_276),
.A2(n_252),
.B1(n_253),
.B2(n_238),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_315),
.A2(n_316),
.B(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_284),
.Y(n_322)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_287),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_323),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_325),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_244),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_334),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_239),
.C(n_259),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_330),
.C(n_286),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_278),
.A2(n_256),
.B1(n_242),
.B2(n_243),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_329),
.A2(n_332),
.B1(n_339),
.B2(n_295),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_276),
.A2(n_268),
.B1(n_252),
.B2(n_251),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_278),
.A2(n_263),
.B1(n_265),
.B2(n_269),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_257),
.B1(n_241),
.B2(n_272),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_274),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_290),
.B(n_4),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_335),
.B(n_306),
.Y(n_365)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_338),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_304),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_289),
.Y(n_361)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_285),
.A2(n_1),
.B1(n_2),
.B2(n_12),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_309),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_341),
.B(n_352),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_300),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_348),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_317),
.B1(n_338),
.B2(n_336),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_300),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_351),
.C(n_356),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_294),
.C(n_283),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_311),
.B(n_296),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_353),
.A2(n_328),
.B(n_325),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_296),
.C(n_277),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_360),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_291),
.C(n_298),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_331),
.B(n_307),
.Y(n_360)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_362),
.A2(n_332),
.B1(n_317),
.B2(n_343),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_288),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_363),
.B(n_365),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_316),
.A2(n_277),
.B(n_279),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_364),
.A2(n_356),
.B(n_344),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_367),
.A2(n_385),
.B1(n_386),
.B2(n_347),
.Y(n_391)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_325),
.B(n_319),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_377),
.B(n_308),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_312),
.Y(n_371)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_319),
.Y(n_372)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_335),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_374),
.B(n_347),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_344),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_315),
.C(n_333),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_378),
.C(n_351),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_353),
.A2(n_328),
.B(n_313),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_337),
.C(n_279),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_326),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_384),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_381),
.A2(n_342),
.B1(n_354),
.B2(n_301),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_310),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_339),
.B1(n_310),
.B2(n_318),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_346),
.A2(n_321),
.B1(n_322),
.B2(n_301),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_387),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_391),
.Y(n_411)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_390),
.Y(n_408)
);

BUFx12_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_396),
.Y(n_413)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_373),
.B1(n_369),
.B2(n_381),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_345),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_397),
.Y(n_405)
);

AOI322xp5_ASAP7_75t_L g396 ( 
.A1(n_379),
.A2(n_354),
.A3(n_342),
.B1(n_364),
.B2(n_360),
.C1(n_355),
.C2(n_352),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_398),
.A2(n_385),
.B1(n_384),
.B2(n_380),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_370),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_341),
.C(n_292),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_401),
.A2(n_402),
.B(n_382),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_292),
.C(n_15),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_415),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_403),
.A2(n_369),
.B1(n_367),
.B2(n_386),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_407),
.A2(n_418),
.B1(n_389),
.B2(n_375),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_410),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_412),
.B(n_414),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_402),
.B(n_368),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_378),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_391),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_387),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_405),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_403),
.A2(n_371),
.B1(n_376),
.B2(n_377),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_408),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_418),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_421),
.A2(n_411),
.B1(n_416),
.B2(n_409),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_400),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_428),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_424),
.B(n_425),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_417),
.B(n_388),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_415),
.C(n_411),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_430),
.Y(n_437)
);

INVx11_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_433),
.B(n_434),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_423),
.B(n_393),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_435),
.B(n_439),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_427),
.B(n_404),
.Y(n_436)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_438),
.Y(n_440)
);

XOR2x1_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_400),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_392),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_437),
.A2(n_432),
.B(n_431),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_441),
.A2(n_445),
.B(n_429),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_420),
.C(n_422),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_443),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_420),
.C(n_429),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_447),
.B(n_448),
.C(n_449),
.Y(n_450)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_440),
.A2(n_404),
.B(n_395),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_442),
.C(n_440),
.Y(n_451)
);

OAI321xp33_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_436),
.A3(n_430),
.B1(n_395),
.B2(n_392),
.C(n_401),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_450),
.B(n_398),
.Y(n_453)
);

BUFx24_ASAP7_75t_SL g454 ( 
.A(n_453),
.Y(n_454)
);

AOI31xp33_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_382),
.A3(n_383),
.B(n_446),
.Y(n_455)
);


endmodule