module fake_netlist_1_12229_n_633 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_633);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_633;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_55), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_13), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_59), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_41), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_63), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_73), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_56), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_45), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_9), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_15), .Y(n_87) );
CKINVDCx14_ASAP7_75t_R g88 ( .A(n_43), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_30), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_5), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_19), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_34), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_42), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_51), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_49), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_6), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_36), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_52), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_50), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_1), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_19), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_64), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_28), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_60), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_23), .B(n_22), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_47), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_24), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_74), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_53), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_6), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_21), .Y(n_116) );
CKINVDCx14_ASAP7_75t_R g117 ( .A(n_58), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_1), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_2), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_86), .Y(n_121) );
AND3x2_ASAP7_75t_L g122 ( .A(n_119), .B(n_2), .C(n_3), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_86), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_76), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
AND2x6_ASAP7_75t_L g128 ( .A(n_80), .B(n_31), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_75), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_75), .Y(n_130) );
NAND2xp33_ASAP7_75t_R g131 ( .A(n_102), .B(n_29), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_78), .Y(n_136) );
INVx5_ASAP7_75t_L g137 ( .A(n_97), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_111), .B(n_4), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_97), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_99), .Y(n_147) );
CKINVDCx8_ASAP7_75t_R g148 ( .A(n_83), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_94), .B(n_4), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
INVxp33_ASAP7_75t_L g154 ( .A(n_76), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_109), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_109), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_117), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_100), .B(n_5), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_154), .B(n_95), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_149), .B(n_105), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_149), .B(n_81), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_139), .B(n_101), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_139), .B(n_101), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_160), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_160), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_129), .B(n_84), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_150), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_148), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_139), .B(n_106), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_148), .B(n_114), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
OAI22xp5_ASAP7_75t_SL g180 ( .A1(n_126), .A2(n_87), .B1(n_96), .B2(n_115), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_139), .B(n_106), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_128), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_124), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_126), .B(n_91), .Y(n_186) );
AND2x6_ASAP7_75t_L g187 ( .A(n_150), .B(n_103), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_127), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_129), .B(n_107), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_130), .B(n_107), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_127), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_140), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_130), .B(n_118), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_132), .B(n_110), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_132), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_140), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_128), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_133), .B(n_110), .Y(n_199) );
BUFx8_ASAP7_75t_SL g200 ( .A(n_141), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_133), .B(n_104), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_127), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_134), .B(n_104), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_128), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_134), .B(n_118), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_136), .B(n_90), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_128), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_136), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_152), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_128), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_138), .B(n_103), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_148), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_138), .B(n_113), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_159), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_159), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_142), .B(n_143), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_137), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_187), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_196), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_163), .B(n_142), .Y(n_223) );
CKINVDCx14_ASAP7_75t_R g224 ( .A(n_170), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_167), .B(n_141), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_213), .Y(n_227) );
BUFx4f_ASAP7_75t_SL g228 ( .A(n_214), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_196), .B(n_143), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_213), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_213), .Y(n_231) );
AND3x2_ASAP7_75t_SL g232 ( .A(n_187), .B(n_131), .C(n_122), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_209), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_209), .B(n_144), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_168), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_162), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_216), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_187), .A2(n_145), .B1(n_158), .B2(n_144), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_216), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
OR2x2_ASAP7_75t_SL g244 ( .A(n_184), .B(n_90), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_162), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_174), .B(n_145), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_187), .A2(n_93), .B1(n_158), .B2(n_151), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_187), .A2(n_146), .B1(n_155), .B2(n_151), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_175), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_206), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_186), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_174), .B(n_146), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_187), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_186), .B(n_155), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_164), .B(n_161), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_175), .Y(n_258) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_201), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_176), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_171), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_186), .B(n_135), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_183), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_173), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_165), .Y(n_265) );
AND2x6_ASAP7_75t_L g266 ( .A(n_175), .B(n_113), .Y(n_266) );
AND2x4_ASAP7_75t_SL g267 ( .A(n_186), .B(n_91), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_180), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_206), .B(n_135), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_206), .B(n_135), .Y(n_270) );
OR2x2_ASAP7_75t_SL g271 ( .A(n_180), .B(n_98), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_167), .B(n_114), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_165), .A2(n_120), .B1(n_112), .B2(n_98), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_169), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_179), .Y(n_275) );
INVx4_ASAP7_75t_L g276 ( .A(n_165), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_165), .A2(n_153), .B1(n_141), .B2(n_157), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_167), .B(n_137), .Y(n_278) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_219), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_206), .B(n_135), .Y(n_280) );
INVxp67_ASAP7_75t_SL g281 ( .A(n_220), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_166), .A2(n_157), .B1(n_153), .B2(n_141), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_265), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_261), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_235), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_279), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_261), .B(n_194), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_253), .B(n_172), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_259), .Y(n_289) );
AO21x1_ASAP7_75t_L g290 ( .A1(n_235), .A2(n_203), .B(n_191), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_221), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_247), .A2(n_195), .B1(n_190), .B2(n_199), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_256), .A2(n_211), .B(n_167), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_242), .Y(n_294) );
CKINVDCx8_ASAP7_75t_R g295 ( .A(n_260), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_224), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_227), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_236), .B(n_178), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_253), .A2(n_177), .B1(n_181), .B2(n_166), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_243), .B(n_166), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_249), .A2(n_177), .B1(n_166), .B2(n_181), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_227), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_226), .A2(n_212), .B(n_215), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_252), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_236), .B(n_200), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_221), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_242), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g309 ( .A1(n_273), .A2(n_194), .B1(n_207), .B2(n_217), .C(n_202), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_230), .Y(n_310) );
BUFx4_ASAP7_75t_R g311 ( .A(n_267), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_222), .A2(n_177), .B1(n_181), .B2(n_207), .Y(n_312) );
BUFx12f_ASAP7_75t_L g313 ( .A(n_260), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_244), .B(n_177), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_233), .B(n_181), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_267), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_265), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_250), .A2(n_211), .B1(n_179), .B2(n_198), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_223), .A2(n_192), .B(n_218), .C(n_217), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_278), .A2(n_211), .B(n_179), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_245), .B(n_211), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_265), .B(n_182), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_257), .A2(n_182), .B1(n_198), .B2(n_205), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_272), .A2(n_182), .B(n_198), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_229), .B(n_189), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_252), .B(n_189), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_240), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_301), .A2(n_238), .B1(n_225), .B2(n_255), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_284), .A2(n_268), .B1(n_228), .B2(n_225), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_285), .Y(n_332) );
INVx5_ASAP7_75t_L g333 ( .A(n_297), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_315), .A2(n_268), .B1(n_276), .B2(n_255), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_286), .B(n_252), .Y(n_335) );
O2A1O1Ixp5_ASAP7_75t_L g336 ( .A1(n_290), .A2(n_246), .B(n_254), .C(n_280), .Y(n_336) );
NAND2x1_ASAP7_75t_L g337 ( .A(n_285), .B(n_231), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_315), .A2(n_276), .B1(n_234), .B2(n_266), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_311), .Y(n_339) );
OAI22xp5_ASAP7_75t_SL g340 ( .A1(n_295), .A2(n_271), .B1(n_244), .B2(n_232), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_315), .A2(n_276), .B1(n_266), .B2(n_262), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_319), .A2(n_248), .B(n_274), .C(n_270), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_294), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_294), .Y(n_344) );
BUFx4f_ASAP7_75t_SL g345 ( .A(n_313), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_300), .B(n_269), .Y(n_346) );
OAI21xp33_ASAP7_75t_SL g347 ( .A1(n_307), .A2(n_274), .B(n_282), .Y(n_347) );
OR2x6_ASAP7_75t_L g348 ( .A(n_300), .B(n_226), .Y(n_348) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_316), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_300), .B(n_226), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_311), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_307), .Y(n_352) );
OAI22xp5_ASAP7_75t_SL g353 ( .A1(n_295), .A2(n_271), .B1(n_232), .B2(n_277), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_308), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_328), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_287), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_344), .A2(n_292), .B1(n_319), .B2(n_299), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_358), .A2(n_314), .B1(n_287), .B2(n_309), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_340), .A2(n_305), .B1(n_314), .B2(n_313), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_348), .B(n_303), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_332), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_353), .A2(n_290), .B1(n_312), .B2(n_298), .C(n_288), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_339), .A2(n_345), .B1(n_351), .B2(n_349), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_344), .A2(n_289), .B1(n_326), .B2(n_291), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_352), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_356), .B(n_303), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_346), .A2(n_296), .B1(n_322), .B2(n_291), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_348), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g372 ( .A1(n_336), .A2(n_293), .B(n_318), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_347), .A2(n_320), .B(n_325), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_348), .Y(n_374) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_331), .A2(n_122), .B(n_306), .Y(n_375) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_347), .A2(n_125), .B(n_121), .C(n_123), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_346), .A2(n_306), .B1(n_304), .B2(n_317), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_357), .A2(n_121), .B1(n_123), .B2(n_125), .C(n_157), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_346), .A2(n_317), .B1(n_266), .B2(n_283), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_356), .B(n_283), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_348), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_352), .B(n_283), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_346), .A2(n_317), .B1(n_266), .B2(n_310), .Y(n_383) );
BUFx6f_ASAP7_75t_SL g384 ( .A(n_348), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_360), .B(n_357), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_375), .B(n_334), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_362), .Y(n_387) );
NAND4xp25_ASAP7_75t_L g388 ( .A(n_364), .B(n_153), .C(n_157), .D(n_338), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_364), .A2(n_335), .B1(n_342), .B2(n_153), .C(n_330), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_361), .A2(n_341), .B1(n_346), .B2(n_350), .C(n_335), .Y(n_390) );
AOI33xp33_ASAP7_75t_L g391 ( .A1(n_365), .A2(n_202), .A3(n_185), .B1(n_192), .B2(n_204), .B3(n_218), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_362), .Y(n_392) );
OAI31xp33_ASAP7_75t_L g393 ( .A1(n_375), .A2(n_355), .A3(n_354), .B(n_343), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_367), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_367), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_369), .A2(n_350), .B1(n_337), .B2(n_355), .C(n_343), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
OAI33xp33_ASAP7_75t_L g399 ( .A1(n_359), .A2(n_185), .A3(n_204), .B1(n_210), .B2(n_173), .B3(n_193), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_368), .B(n_332), .Y(n_400) );
OAI31xp33_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_354), .A3(n_232), .B(n_116), .Y(n_401) );
OAI211xp5_ASAP7_75t_L g402 ( .A1(n_370), .A2(n_82), .B(n_210), .C(n_337), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_384), .A2(n_350), .B1(n_333), .B2(n_329), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_363), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_382), .B(n_350), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_382), .B(n_350), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_362), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_362), .B(n_333), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_366), .A2(n_333), .B(n_329), .Y(n_410) );
OAI33xp33_ASAP7_75t_L g411 ( .A1(n_359), .A2(n_173), .A3(n_188), .B1(n_193), .B2(n_197), .B3(n_11), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_378), .A2(n_147), .B1(n_156), .B2(n_140), .C(n_137), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_371), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_376), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_384), .A2(n_266), .B1(n_323), .B2(n_231), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_380), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_384), .A2(n_266), .B1(n_323), .B2(n_231), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
OAI33xp33_ASAP7_75t_L g419 ( .A1(n_381), .A2(n_188), .A3(n_193), .B1(n_197), .B2(n_10), .B3(n_11), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_394), .B(n_374), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_394), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_404), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_400), .B(n_371), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_388), .B(n_378), .C(n_374), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g426 ( .A1(n_386), .A2(n_390), .B(n_385), .C(n_419), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_400), .B(n_380), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_393), .B(n_147), .C(n_156), .Y(n_428) );
BUFx2_ASAP7_75t_SL g429 ( .A(n_409), .Y(n_429) );
INVx2_ASAP7_75t_SL g430 ( .A(n_409), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_395), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_404), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_405), .B(n_372), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_414), .A2(n_384), .B1(n_377), .B2(n_379), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_414), .A2(n_373), .B(n_372), .Y(n_438) );
OAI33xp33_ASAP7_75t_L g439 ( .A1(n_418), .A2(n_7), .A3(n_8), .B1(n_9), .B2(n_12), .B3(n_13), .Y(n_439) );
AND4x1_ASAP7_75t_L g440 ( .A(n_391), .B(n_383), .C(n_108), .D(n_12), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_416), .Y(n_441) );
AND2x4_ASAP7_75t_SL g442 ( .A(n_409), .B(n_302), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_389), .A2(n_418), .B1(n_411), .B2(n_407), .C1(n_406), .C2(n_399), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_416), .Y(n_444) );
OAI33xp33_ASAP7_75t_L g445 ( .A1(n_408), .A2(n_7), .A3(n_8), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_445) );
AOI32xp33_ASAP7_75t_L g446 ( .A1(n_406), .A2(n_14), .A3(n_16), .B1(n_17), .B2(n_18), .Y(n_446) );
OAI31xp33_ASAP7_75t_L g447 ( .A1(n_402), .A2(n_373), .A3(n_321), .B(n_310), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_401), .A2(n_147), .B1(n_156), .B2(n_321), .C(n_333), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_387), .B(n_333), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_408), .A2(n_17), .A3(n_20), .B1(n_197), .B2(n_188), .B3(n_156), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_387), .B(n_156), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_392), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_392), .B(n_333), .Y(n_456) );
OAI33xp33_ASAP7_75t_L g457 ( .A1(n_397), .A2(n_20), .A3(n_147), .B1(n_156), .B2(n_137), .B3(n_239), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_403), .B(n_237), .C(n_323), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_413), .A2(n_137), .B1(n_147), .B2(n_239), .C1(n_297), .C2(n_302), .Y(n_459) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_410), .A2(n_324), .B(n_264), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_412), .B(n_147), .C(n_137), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_392), .B(n_137), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_415), .B(n_329), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_417), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_394), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_394), .B(n_329), .Y(n_466) );
OAI322xp33_ASAP7_75t_L g467 ( .A1(n_386), .A2(n_237), .A3(n_264), .B1(n_263), .B2(n_241), .C1(n_327), .C2(n_297), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_394), .Y(n_468) );
AOI33xp33_ASAP7_75t_L g469 ( .A1(n_394), .A2(n_263), .A3(n_241), .B1(n_220), .B2(n_33), .B3(n_35), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_436), .B(n_25), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_446), .B(n_327), .C(n_302), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_441), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_422), .B(n_327), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_450), .B(n_26), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_425), .A2(n_327), .B1(n_302), .B2(n_297), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_427), .B(n_237), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_427), .B(n_27), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_436), .B(n_38), .Y(n_479) );
NAND3xp33_ASAP7_75t_SL g480 ( .A(n_440), .B(n_39), .C(n_40), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_465), .B(n_423), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_421), .B(n_424), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_465), .B(n_44), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_454), .B(n_46), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_468), .B(n_48), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_432), .B(n_54), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_449), .B(n_57), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_438), .B(n_61), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_423), .B(n_62), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_444), .B(n_66), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_433), .B(n_67), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_454), .B(n_438), .Y(n_492) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_469), .B(n_208), .C(n_205), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_438), .B(n_68), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_435), .B(n_69), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_426), .B(n_70), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_430), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_442), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_430), .A2(n_205), .B1(n_208), .B2(n_281), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_429), .B(n_72), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_443), .B(n_208), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_420), .B(n_251), .Y(n_503) );
NOR3xp33_ASAP7_75t_SL g504 ( .A(n_439), .B(n_445), .C(n_457), .Y(n_504) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_442), .B(n_469), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_429), .B(n_251), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_455), .B(n_251), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_453), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_456), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_460), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_451), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_451), .B(n_251), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_456), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_251), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_462), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_462), .Y(n_518) );
AOI31xp33_ASAP7_75t_SL g519 ( .A1(n_458), .A2(n_258), .A3(n_275), .B(n_437), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_464), .B(n_258), .Y(n_520) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_463), .B(n_467), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_481), .B(n_459), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_473), .B(n_428), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_497), .B(n_452), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_509), .B(n_447), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_492), .B(n_461), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_509), .B(n_448), .Y(n_528) );
AND2x2_ASAP7_75t_SL g529 ( .A(n_498), .B(n_258), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_512), .B(n_258), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_505), .A2(n_275), .B(n_521), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_510), .B(n_275), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_499), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g534 ( .A(n_480), .B(n_275), .C(n_471), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_472), .B(n_275), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_482), .Y(n_536) );
AND2x4_ASAP7_75t_SL g537 ( .A(n_514), .B(n_501), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_505), .A2(n_471), .B1(n_521), .B2(n_518), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_499), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_495), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_508), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_514), .B(n_516), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_514), .B(n_518), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_516), .B(n_474), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_504), .B(n_476), .C(n_522), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_522), .B(n_494), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_505), .B(n_478), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_521), .A2(n_493), .B(n_488), .Y(n_549) );
AOI21xp33_ASAP7_75t_L g550 ( .A1(n_488), .A2(n_475), .B(n_502), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_483), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_511), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_477), .B(n_489), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_489), .B(n_487), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_494), .B(n_470), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_511), .B(n_517), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_501), .A2(n_487), .B(n_493), .C(n_519), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_517), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_470), .B(n_479), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_479), .A2(n_486), .B1(n_485), .B2(n_491), .C(n_490), .Y(n_561) );
BUFx2_ASAP7_75t_L g562 ( .A(n_539), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_536), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_545), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_533), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_538), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_547), .Y(n_568) );
XNOR2xp5_ASAP7_75t_L g569 ( .A(n_543), .B(n_496), .Y(n_569) );
AOI21xp33_ASAP7_75t_SL g570 ( .A1(n_529), .A2(n_519), .B(n_486), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_542), .Y(n_571) );
NAND2x1_ASAP7_75t_L g572 ( .A(n_540), .B(n_531), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_544), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_537), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_554), .A2(n_484), .B1(n_513), .B2(n_496), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_541), .Y(n_576) );
NAND3x1_ASAP7_75t_L g577 ( .A(n_549), .B(n_506), .C(n_507), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_558), .A2(n_484), .B(n_506), .Y(n_578) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_558), .B(n_484), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_528), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_548), .A2(n_515), .B1(n_503), .B2(n_500), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_556), .Y(n_582) );
AND2x2_ASAP7_75t_SL g583 ( .A(n_537), .B(n_520), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_546), .B(n_527), .Y(n_584) );
O2A1O1Ixp5_ASAP7_75t_SL g585 ( .A1(n_550), .A2(n_526), .B(n_523), .C(n_535), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_546), .B(n_525), .Y(n_586) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_525), .A2(n_548), .B(n_524), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_524), .Y(n_588) );
OA22x2_ASAP7_75t_L g589 ( .A1(n_555), .A2(n_560), .B1(n_557), .B2(n_551), .Y(n_589) );
O2A1O1Ixp5_ASAP7_75t_SL g590 ( .A1(n_534), .A2(n_529), .B(n_561), .C(n_552), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_553), .B(n_559), .Y(n_591) );
NAND4xp75_ASAP7_75t_L g592 ( .A(n_532), .B(n_538), .C(n_531), .D(n_549), .Y(n_592) );
BUFx3_ASAP7_75t_L g593 ( .A(n_530), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_532), .B(n_559), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_537), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_536), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_548), .A2(n_538), .B1(n_525), .B2(n_545), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_531), .A2(n_549), .B(n_538), .C(n_558), .Y(n_598) );
XNOR2x1_ASAP7_75t_L g599 ( .A(n_538), .B(n_268), .Y(n_599) );
XNOR2x1_ASAP7_75t_L g600 ( .A(n_538), .B(n_268), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_565), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_566), .B(n_588), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_591), .Y(n_603) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_564), .A2(n_589), .B(n_566), .Y(n_604) );
OAI21xp33_ASAP7_75t_SL g605 ( .A1(n_579), .A2(n_583), .B(n_592), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_598), .B(n_578), .Y(n_606) );
AOI222xp33_ASAP7_75t_L g607 ( .A1(n_564), .A2(n_567), .B1(n_586), .B2(n_580), .C1(n_563), .C2(n_596), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_584), .Y(n_609) );
NOR4xp25_ASAP7_75t_L g610 ( .A(n_587), .B(n_577), .C(n_567), .D(n_568), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_597), .A2(n_578), .B(n_570), .Y(n_611) );
AOI211x1_ASAP7_75t_SL g612 ( .A1(n_585), .A2(n_575), .B(n_600), .C(n_599), .Y(n_612) );
XOR2xp5_ASAP7_75t_L g613 ( .A(n_569), .B(n_594), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_611), .A2(n_577), .B1(n_574), .B2(n_595), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_608), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_606), .B(n_590), .C(n_576), .Y(n_616) );
OAI221xp5_ASAP7_75t_R g617 ( .A1(n_613), .A2(n_581), .B1(n_595), .B2(n_573), .C(n_572), .Y(n_617) );
XNOR2x1_ASAP7_75t_L g618 ( .A(n_601), .B(n_602), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_606), .B(n_593), .Y(n_619) );
OAI31xp33_ASAP7_75t_L g620 ( .A1(n_610), .A2(n_575), .A3(n_571), .B(n_582), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_619), .A2(n_605), .B(n_604), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_615), .B(n_609), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_616), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_620), .B(n_612), .C(n_607), .D(n_603), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_622), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_623), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_624), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_625), .B(n_621), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_627), .B(n_614), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_628), .B(n_627), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_630), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_631), .A2(n_629), .B1(n_626), .B2(n_618), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_632), .A2(n_601), .B(n_617), .Y(n_633) );
endmodule