module fake_jpeg_28496_n_100 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_7),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_0),
.C(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_2),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_16),
.C(n_28),
.Y(n_48)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_42),
.CI(n_4),
.CON(n_55),
.SN(n_55)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_3),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_36),
.B1(n_40),
.B2(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_52),
.B1(n_8),
.B2(n_9),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_36),
.B1(n_40),
.B2(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_5),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_3),
.C(n_4),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_5),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_72),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_14),
.B(n_27),
.C(n_26),
.D(n_25),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_17),
.B(n_24),
.C(n_23),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_6),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_13),
.B1(n_22),
.B2(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_74),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_9),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_64),
.C(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.C(n_88),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_63),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_57),
.B1(n_58),
.B2(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_93),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_82),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_92),
.Y(n_97)
);

AOI321xp33_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_86),
.A3(n_79),
.B1(n_90),
.B2(n_76),
.C(n_75),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_98),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_57),
.Y(n_100)
);


endmodule