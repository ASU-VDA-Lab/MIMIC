module fake_jpeg_20159_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_31),
.B1(n_19),
.B2(n_23),
.Y(n_54)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_35),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_33),
.B1(n_28),
.B2(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_71),
.B(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_72),
.A2(n_86),
.B1(n_95),
.B2(n_97),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_57),
.B1(n_63),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_84),
.B1(n_100),
.B2(n_101),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_59),
.B(n_19),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_36),
.B(n_34),
.C(n_25),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_49),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_90),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_53),
.B1(n_36),
.B2(n_22),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_24),
.B1(n_28),
.B2(n_17),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_36),
.B(n_35),
.C(n_29),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_33),
.B1(n_21),
.B2(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2x1_ASAP7_75t_R g91 ( 
.A(n_56),
.B(n_36),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_94),
.Y(n_114)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_50),
.B1(n_44),
.B2(n_46),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

AO22x2_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_45),
.B1(n_43),
.B2(n_39),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_52),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_27),
.B1(n_39),
.B2(n_38),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_43),
.B1(n_35),
.B2(n_29),
.Y(n_101)
);

NAND2x1p5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_52),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_112),
.B(n_97),
.Y(n_145)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_111),
.Y(n_160)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_109),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_90),
.B1(n_94),
.B2(n_99),
.Y(n_136)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_123),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_34),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_25),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_92),
.B1(n_1),
.B2(n_2),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_68),
.A2(n_36),
.B1(n_22),
.B2(n_25),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_95),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_68),
.B1(n_85),
.B2(n_72),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_134),
.A2(n_10),
.B1(n_14),
.B2(n_6),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_99),
.B1(n_75),
.B2(n_87),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_77),
.B(n_89),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_116),
.B(n_118),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_97),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_88),
.B(n_93),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_76),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_151),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_89),
.C(n_98),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_129),
.C(n_104),
.Y(n_169)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_96),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_35),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_158),
.B(n_159),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_156),
.B1(n_113),
.B2(n_105),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_29),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_102),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_0),
.B(n_1),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_10),
.B1(n_15),
.B2(n_6),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_131),
.B1(n_113),
.B2(n_107),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

AO21x2_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_128),
.B(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_177),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_191),
.B1(n_154),
.B2(n_153),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_173),
.C(n_175),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_179),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_102),
.C(n_116),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_122),
.B(n_109),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_145),
.B(n_158),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_104),
.C(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_185),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_144),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_131),
.B1(n_127),
.B2(n_111),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_180),
.B1(n_153),
.B2(n_149),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_133),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_139),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_143),
.A2(n_127),
.B1(n_125),
.B2(n_106),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_190),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_16),
.C(n_9),
.Y(n_190)
);

AO21x2_ASAP7_75t_L g191 ( 
.A1(n_136),
.A2(n_3),
.B(n_4),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_176),
.B(n_182),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_199),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_161),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_202),
.B(n_211),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_146),
.B(n_152),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_216),
.B1(n_218),
.B2(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_139),
.B(n_160),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_213),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_190),
.B(n_135),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_169),
.B(n_10),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_250),
.B1(n_213),
.B2(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_179),
.C(n_178),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_229),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_172),
.C(n_139),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_167),
.B1(n_191),
.B2(n_6),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_210),
.B1(n_217),
.B2(n_232),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_241),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_167),
.C(n_191),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_247),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_210),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_205),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_193),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_195),
.A2(n_167),
.B1(n_191),
.B2(n_3),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_199),
.B(n_209),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_235),
.B(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_266),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_258),
.B1(n_240),
.B2(n_244),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_195),
.B1(n_220),
.B2(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_201),
.C(n_197),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_201),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_206),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_193),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_231),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_271),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_240),
.A2(n_214),
.B(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_246),
.B1(n_249),
.B2(n_242),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_229),
.C(n_243),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_281),
.C(n_285),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_237),
.B1(n_242),
.B2(n_246),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_234),
.C(n_233),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_234),
.C(n_231),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_288),
.B(n_226),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_198),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_263),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_214),
.B1(n_239),
.B2(n_232),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_265),
.B1(n_226),
.B2(n_251),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_259),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_260),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_300),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_252),
.Y(n_294)
);

XOR2x1_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_239),
.Y(n_296)
);

FAx1_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_290),
.CI(n_288),
.CON(n_310),
.SN(n_310)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_262),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_301),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_258),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_302),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_283),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_261),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_275),
.A2(n_269),
.B(n_266),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_287),
.B(n_296),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_306),
.C(n_273),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_268),
.B1(n_251),
.B2(n_265),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_274),
.B1(n_272),
.B2(n_282),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_309),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_291),
.A2(n_274),
.B1(n_272),
.B2(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_316),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_277),
.C(n_276),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_318),
.C(n_292),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_287),
.C(n_196),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_321),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_326),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_301),
.C(n_306),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_196),
.C(n_167),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_310),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_191),
.CI(n_7),
.CON(n_324),
.SN(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_8),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_310),
.B1(n_314),
.B2(n_16),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_312),
.B(n_311),
.Y(n_329)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_307),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_325),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_331),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_319),
.C(n_334),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_320),
.C(n_335),
.Y(n_341)
);

AOI221xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_336),
.B1(n_328),
.B2(n_321),
.C(n_326),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_16),
.C(n_13),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_13),
.B(n_4),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_13),
.Y(n_345)
);


endmodule