module real_jpeg_5187_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_0),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_0),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_0),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_0),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_0),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_0),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_0),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_0),
.B(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_1),
.Y(n_169)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_1),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_1),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_2),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_3),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_3),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_4),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_4),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_4),
.B(n_146),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_4),
.B(n_211),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_4),
.B(n_296),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_4),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_5),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_5),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_5),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_5),
.B(n_323),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_5),
.B(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_5),
.B(n_221),
.Y(n_423)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_6),
.Y(n_413)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_7),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_8),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_8),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_8),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_8),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_8),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_8),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_9),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_9),
.Y(n_362)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_11),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_11),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_13),
.B(n_100),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_13),
.B(n_87),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_13),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_13),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_13),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_13),
.B(n_395),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_13),
.B(n_407),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_14),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_14),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_14),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_15),
.B(n_59),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_15),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_15),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_15),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_15),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_15),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_15),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_15),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_16),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_16),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_16),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_16),
.B(n_59),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_16),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_16),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_16),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_17),
.B(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_17),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_17),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_17),
.B(n_323),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_17),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_17),
.B(n_421),
.Y(n_420)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_19),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_19),
.B(n_194),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_19),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_19),
.B(n_69),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_19),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_19),
.B(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_19),
.B(n_411),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_544),
.B(n_547),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_77),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_48),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.C(n_35),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_26),
.A2(n_31),
.B1(n_40),
.B2(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_29),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_52),
.C(n_58),
.Y(n_74)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_33),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_34),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_34),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_38),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_73),
.C(n_75),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_49),
.B(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_62),
.C(n_63),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_50),
.B(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_52),
.A2(n_57),
.B1(n_68),
.B2(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_53),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_55),
.Y(n_360)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_55),
.Y(n_397)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_55),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_64),
.C(n_68),
.Y(n_63)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_60),
.B(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_63),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_64),
.A2(n_65),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_68),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_68),
.A2(n_116),
.B1(n_117),
.B2(n_123),
.Y(n_513)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_71),
.Y(n_231)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_72),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_72),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_72),
.Y(n_356)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_72),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_134),
.B(n_543),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_131),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_80),
.B(n_131),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_128),
.C(n_129),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_81),
.A2(n_82),
.B1(n_539),
.B2(n_540),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_111),
.C(n_124),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_83),
.A2(n_84),
.B1(n_517),
.B2(n_519),
.Y(n_516)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_96),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_90),
.C(n_96),
.Y(n_128)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_108),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_97),
.B(n_507),
.Y(n_506)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_100),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_101),
.A2(n_102),
.B1(n_108),
.B2(n_109),
.Y(n_507)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_111),
.A2(n_124),
.B1(n_125),
.B2(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_111),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_123),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_112),
.B(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_116),
.A2(n_117),
.B1(n_210),
.B2(n_213),
.Y(n_209)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_117),
.B(n_206),
.C(n_210),
.Y(n_514)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g422 ( 
.A(n_122),
.Y(n_422)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_128),
.B(n_129),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_537),
.B(n_542),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_500),
.B(n_534),
.Y(n_135)
);

OAI21x1_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_302),
.B(n_499),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_253),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_138),
.B(n_253),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_203),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_139),
.B(n_204),
.C(n_234),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_171),
.C(n_182),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_140),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_149),
.C(n_158),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_141),
.B(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_149),
.A2(n_150),
.B1(n_158),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.C(n_154),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_151),
.B(n_154),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_152),
.B(n_475),
.Y(n_474)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_158),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_159),
.B(n_163),
.C(n_168),
.Y(n_250)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_167),
.B(n_210),
.C(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_167),
.A2(n_168),
.B1(n_210),
.B2(n_213),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_171),
.B(n_182),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_181),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_177),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_177),
.B(n_179),
.C(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_177),
.A2(n_180),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_178),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_180),
.B(n_239),
.C(n_246),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.C(n_198),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_183),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.C(n_190),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_184),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_186),
.B(n_190),
.Y(n_265)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_189),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_189),
.Y(n_380)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_192),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_192),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_193),
.B(n_198),
.Y(n_282)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_197),
.Y(n_290)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_202),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_202),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_234),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_214),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_205),
.B(n_215),
.C(n_233),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_210),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_212),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g332 ( 
.A(n_212),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_223),
.B1(n_232),
.B2(n_233),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_220),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_219),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_224),
.B(n_226),
.C(n_229),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_247),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_236),
.B(n_238),
.C(n_247),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.C(n_251),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_255),
.B(n_258),
.Y(n_495)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_260),
.B(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_280),
.C(n_283),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_262),
.B(n_488),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_272),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_263),
.A2(n_264),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_266),
.A2(n_267),
.B(n_269),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_266),
.B(n_272),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.C(n_277),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_443)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_277),
.B(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_279),
.B(n_373),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_283),
.Y(n_489)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_295),
.C(n_299),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_285),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.C(n_291),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_286),
.B(n_455),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_288),
.A2(n_291),
.B1(n_292),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_288),
.Y(n_456)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_295),
.B(n_299),
.Y(n_477)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_298),
.Y(n_338)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_493),
.B(n_498),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_480),
.B(n_492),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_462),
.B(n_479),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_436),
.B(n_461),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_401),
.B(n_435),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_365),
.B(n_400),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_342),
.B(n_364),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_326),
.B(n_341),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_321),
.B(n_325),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_320),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_320),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_316),
.Y(n_327)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_315),
.Y(n_429)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_328),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_334),
.B2(n_335),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_337),
.C(n_339),
.Y(n_363)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_333),
.Y(n_350)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_363),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_363),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_351),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_350),
.C(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_349),
.Y(n_370)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_351),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_357),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_384),
.C(n_385),
.Y(n_383)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_368),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_382),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_369),
.B(n_383),
.C(n_386),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_372),
.C(n_375),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_378),
.B1(n_379),
.B2(n_381),
.Y(n_375)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_376),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_377),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_381),
.Y(n_414)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_394),
.C(n_398),
.Y(n_433)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_391),
.A2(n_394),
.B1(n_398),
.B2(n_399),
.Y(n_390)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_391),
.Y(n_398)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_394),
.Y(n_399)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_434),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_434),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_416),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_415),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_404),
.B(n_415),
.C(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_414),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_410),
.Y(n_405)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_406),
.Y(n_450)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_450),
.C(n_451),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_424),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_426),
.C(n_432),
.Y(n_439)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_417),
.Y(n_550)
);

FAx1_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_420),
.CI(n_423),
.CON(n_417),
.SN(n_417)
);

MAJx2_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_420),
.C(n_423),
.Y(n_447)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_432),
.B2(n_433),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_430),
.Y(n_446)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_459),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_459),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_448),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_440),
.C(n_448),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_441),
.A2(n_442),
.B1(n_444),
.B2(n_445),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_471),
.C(n_472),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_453),
.C(n_458),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_454),
.B1(n_457),
.B2(n_458),
.Y(n_452)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_453),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_454),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_478),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_478),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_469),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_468),
.C(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_474),
.C(n_476),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_490),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_490),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_482),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_487),
.C(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_496),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_529),
.Y(n_500)
);

OAI21xp33_ASAP7_75t_L g534 ( 
.A1(n_501),
.A2(n_535),
.B(n_536),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_521),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_502),
.B(n_521),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_510),
.B2(n_520),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_511),
.C(n_516),
.Y(n_541)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.C(n_508),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_505),
.B(n_524),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_506),
.A2(n_508),
.B1(n_509),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_506),
.Y(n_525)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_516),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.C(n_515),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_512),
.B(n_527),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_515),
.Y(n_527)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_517),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_526),
.C(n_528),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_522),
.A2(n_523),
.B1(n_526),
.B2(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_526),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_531),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_530),
.B(n_533),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_533),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_538),
.B(n_541),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_541),
.Y(n_542)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx13_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_546),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_549),
.Y(n_547)
);


endmodule