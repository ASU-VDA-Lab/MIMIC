module fake_jpeg_26237_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_17),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_55),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_36),
.Y(n_91)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_61),
.B(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_64),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_39),
.C(n_34),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_87),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_27),
.B1(n_16),
.B2(n_35),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_17),
.B1(n_27),
.B2(n_16),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_17),
.B1(n_29),
.B2(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_68),
.A2(n_30),
.B1(n_19),
.B2(n_26),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_R g69 ( 
.A(n_50),
.B(n_19),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_84),
.C(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_75),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_42),
.B1(n_41),
.B2(n_36),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_20),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_47),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_18),
.B(n_24),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_71),
.B(n_23),
.Y(n_146)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_88),
.B1(n_73),
.B2(n_76),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_24),
.B1(n_18),
.B2(n_30),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_119),
.B(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_113),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_63),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_142),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_81),
.B1(n_78),
.B2(n_92),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_132),
.B1(n_145),
.B2(n_150),
.Y(n_167)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_75),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_139),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_85),
.B1(n_73),
.B2(n_76),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_78),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_112),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_79),
.B1(n_80),
.B2(n_61),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_121),
.B1(n_104),
.B2(n_86),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_117),
.B1(n_98),
.B2(n_109),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_82),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_22),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_71),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_66),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_146),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_107),
.B1(n_118),
.B2(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_99),
.B(n_107),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_82),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_151),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_80),
.B1(n_72),
.B2(n_34),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_150),
.B1(n_132),
.B2(n_127),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_124),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_154),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_157),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_126),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_100),
.B(n_105),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_176),
.B(n_184),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_123),
.C(n_105),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_161),
.B(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_169),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_100),
.B1(n_104),
.B2(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_21),
.B1(n_31),
.B2(n_9),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_129),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_172),
.A2(n_173),
.B1(n_188),
.B2(n_0),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_41),
.C(n_86),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_19),
.B(n_31),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_177),
.B(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_38),
.B1(n_26),
.B2(n_22),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_181),
.A2(n_183),
.B1(n_179),
.B2(n_176),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_38),
.C(n_33),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_0),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_26),
.B1(n_22),
.B2(n_115),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_33),
.B1(n_23),
.B2(n_21),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_204),
.B(n_179),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_198),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_130),
.B(n_1),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_33),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_210),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_31),
.B1(n_23),
.B2(n_21),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_211),
.B1(n_184),
.B2(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_15),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_12),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_156),
.B(n_14),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_13),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_220),
.A2(n_222),
.B1(n_190),
.B2(n_213),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_157),
.C(n_163),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_223),
.C(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_155),
.C(n_182),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_184),
.B1(n_171),
.B2(n_181),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_215),
.B1(n_209),
.B2(n_204),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_226),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_166),
.C(n_13),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_201),
.C(n_196),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_189),
.Y(n_246)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

HAxp5_ASAP7_75t_SL g239 ( 
.A(n_203),
.B(n_13),
.CON(n_239),
.SN(n_239)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_9),
.C(n_12),
.Y(n_256)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_212),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_241),
.B(n_216),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_250),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_190),
.B1(n_208),
.B2(n_198),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_255),
.B1(n_262),
.B2(n_235),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_248),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_189),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_258),
.B1(n_261),
.B2(n_236),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_253),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_259),
.B(n_228),
.Y(n_271)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_242),
.B(n_237),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_230),
.B(n_193),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_222),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_219),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_231),
.C(n_225),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_266),
.C(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_225),
.C(n_233),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_268),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_227),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_224),
.C(n_220),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_252),
.C(n_229),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_249),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

AO221x1_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_251),
.B1(n_245),
.B2(n_234),
.C(n_229),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_286),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_289),
.Y(n_294)
);

NOR4xp25_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_245),
.C(n_243),
.D(n_241),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_2),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_236),
.C(n_10),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.C(n_1),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_7),
.C(n_2),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_273),
.B1(n_279),
.B2(n_263),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_304),
.B1(n_290),
.B2(n_285),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_270),
.B1(n_269),
.B2(n_3),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_297),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_270),
.B1(n_2),
.B2(n_3),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_283),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_2),
.C(n_3),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_293),
.C(n_288),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_5),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_309),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_300),
.B1(n_298),
.B2(n_295),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_304),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_281),
.C(n_6),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_294),
.B(n_299),
.Y(n_313)
);

AOI221xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_306),
.B1(n_308),
.B2(n_305),
.C(n_302),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_315),
.B1(n_314),
.B2(n_317),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_312),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

NAND2x1_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_310),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_6),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_7),
.Y(n_325)
);


endmodule