module real_jpeg_5091_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_366;
wire n_149;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_2),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_2),
.A2(n_88),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_2),
.A2(n_88),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_2),
.A2(n_88),
.B1(n_250),
.B2(n_328),
.Y(n_327)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_3),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_45),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_4),
.A2(n_45),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_5),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_5),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_6),
.A2(n_105),
.B1(n_186),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_6),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_6),
.A2(n_178),
.B1(n_258),
.B2(n_298),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_6),
.A2(n_258),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_6),
.A2(n_258),
.B1(n_405),
.B2(n_408),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_9),
.A2(n_140),
.B1(n_142),
.B2(n_145),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_9),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_145),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_9),
.A2(n_145),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_9),
.A2(n_29),
.B1(n_145),
.B2(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_11),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_11),
.A2(n_29),
.B1(n_75),
.B2(n_163),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_75),
.B1(n_179),
.B2(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_12),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_12),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_12),
.A2(n_187),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_12),
.A2(n_37),
.B1(n_187),
.B2(n_371),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_12),
.A2(n_187),
.B1(n_432),
.B2(n_434),
.Y(n_431)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_13),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_13),
.A2(n_238),
.B1(n_276),
.B2(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_13),
.B(n_365),
.C(n_366),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_13),
.B(n_133),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_13),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_13),
.B(n_82),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_13),
.B(n_270),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_14),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_15),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_15),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_15),
.A2(n_103),
.B1(n_140),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_15),
.A2(n_77),
.B1(n_103),
.B2(n_287),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_15),
.A2(n_103),
.B1(n_329),
.B2(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_16),
.A2(n_36),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_218),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_216),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_192),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_20),
.B(n_192),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_116),
.C(n_159),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_21),
.A2(n_22),
.B1(n_116),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_23),
.A2(n_24),
.B(n_85),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_84),
.B1(n_85),
.B2(n_115),
.Y(n_83)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_24),
.A2(n_43),
.B1(n_115),
.B2(n_343),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_25),
.A2(n_35),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_25),
.A2(n_241),
.B1(n_244),
.B2(n_247),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_25),
.A2(n_370),
.B(n_374),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_25),
.A2(n_238),
.B(n_374),
.Y(n_401)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_26),
.A2(n_248),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_26),
.A2(n_242),
.B1(n_327),
.B2(n_332),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_26),
.B(n_377),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_26),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_28),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_28),
.Y(n_400)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_28),
.Y(n_412)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_30),
.Y(n_243)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_31),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_31),
.Y(n_407)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_39),
.Y(n_409)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_43),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_53),
.B1(n_74),
.B2(n_82),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_44),
.A2(n_53),
.B1(n_82),
.B2(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_46),
.Y(n_275)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AO22x2_ASAP7_75t_L g133 ( 
.A1(n_47),
.A2(n_65),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_48),
.Y(n_288)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_48),
.Y(n_385)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_48),
.Y(n_448)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_49),
.Y(n_170)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_52),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_53),
.A2(n_74),
.B1(n_82),
.B2(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_53),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_53),
.B(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_66),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_65),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_58),
.Y(n_174)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx11_ASAP7_75t_L g383 ( 
.A(n_65),
.Y(n_383)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_66),
.A2(n_285),
.B(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_69),
.Y(n_250)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_70),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_71),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_71),
.Y(n_253)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_78),
.Y(n_277)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_81),
.Y(n_433)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_82),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_82),
.B(n_286),
.Y(n_360)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_101),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_91),
.B(n_102),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_91),
.Y(n_198)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_92),
.A2(n_183),
.B1(n_184),
.B2(n_257),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_92),
.B(n_238),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_97),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_99),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_99),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_105),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_101),
.A2(n_198),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_109),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_109),
.A2(n_291),
.B(n_295),
.Y(n_290)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_113),
.Y(n_232)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_114),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_114),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_116),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_152),
.B(n_158),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_153),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_133),
.B1(n_138),
.B2(n_146),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_119),
.A2(n_261),
.B(n_267),
.Y(n_260)
);

AOI22x1_ASAP7_75t_L g306 ( 
.A1(n_119),
.A2(n_133),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_119),
.B(n_307),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_119),
.A2(n_267),
.B(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_120),
.A2(n_139),
.B1(n_176),
.B2(n_181),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_120),
.A2(n_181),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_120),
.A2(n_181),
.B1(n_262),
.B2(n_297),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_133),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_125),
.Y(n_445)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_127),
.Y(n_270)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_132),
.Y(n_299)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_136),
.Y(n_449)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g437 ( 
.A1(n_142),
.A2(n_238),
.B(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_155),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_193),
.CI(n_194),
.CON(n_192),
.SN(n_192)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_159),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_175),
.C(n_182),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_160),
.B(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_161),
.B(n_168),
.Y(n_312)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_162),
.Y(n_280)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_163),
.Y(n_378)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_164),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_169),
.Y(n_278)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_174),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_175),
.B(n_182),
.Y(n_341)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_176),
.Y(n_308)
);

AOI32xp33_ASAP7_75t_L g443 ( 
.A1(n_178),
.A2(n_288),
.A3(n_439),
.B1(n_444),
.B2(n_446),
.Y(n_443)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_181),
.B(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_181),
.A2(n_297),
.B(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B(n_191),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_196)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_190),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_191),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_192),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_204),
.B2(n_215),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_208),
.B1(n_209),
.B2(n_214),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_206),
.A2(n_207),
.B1(n_274),
.B2(n_278),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_206),
.A2(n_358),
.B(n_360),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_206),
.A2(n_207),
.B1(n_382),
.B2(n_431),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_206),
.A2(n_360),
.B(n_431),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_207),
.A2(n_274),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI311xp33_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_337),
.A3(n_351),
.B1(n_468),
.C1(n_473),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_315),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_222),
.A2(n_470),
.B(n_471),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_300),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_223),
.B(n_300),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_271),
.C(n_283),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_224),
.B(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_254),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_225),
.B(n_255),
.C(n_260),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_239),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_226),
.A2(n_239),
.B1(n_240),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_229),
.A3(n_230),
.B1(n_233),
.B2(n_237),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_234),
.Y(n_233)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g291 ( 
.A1(n_237),
.A2(n_238),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_253),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_271),
.A2(n_272),
.B1(n_283),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_279),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_273),
.B(n_279),
.Y(n_304)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.C(n_296),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_284),
.B(n_296),
.Y(n_318)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_290),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_312),
.C(n_313),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_306),
.C(n_311),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_306),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_334),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_316),
.B(n_334),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.C(n_323),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_317),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_320),
.A2(n_321),
.B1(n_323),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_323),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.C(n_333),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_324),
.B(n_459),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_326),
.B(n_333),
.Y(n_459)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_327),
.Y(n_442)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_348),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g468 ( 
.A1(n_338),
.A2(n_348),
.B(n_469),
.C(n_472),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_345),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_339),
.B(n_345),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.C(n_344),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_340),
.B(n_342),
.CI(n_344),
.CON(n_350),
.SN(n_350)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_349),
.B(n_350),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_350),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_462),
.B(n_467),
.Y(n_351)
);

AO21x1_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_451),
.B(n_461),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_425),
.B(n_450),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_388),
.B(n_424),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_368),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_368),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_361),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_357),
.A2(n_361),
.B1(n_362),
.B2(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_379),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_369),
.B(n_380),
.C(n_387),
.Y(n_426)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_381),
.B1(n_386),
.B2(n_387),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_416),
.B(n_423),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_402),
.B(n_415),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_401),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_398),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_399),
.Y(n_420)
);

INVx8_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_414),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_414),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_410),
.B(n_413),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_404),
.Y(n_418)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_412),
.A2(n_413),
.B(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_421),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_421),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_427),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_440),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_435),
.B2(n_436),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_435),
.C(n_440),
.Y(n_452)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_443),
.Y(n_457)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_452),
.B(n_453),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_458),
.B2(n_460),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_457),
.C(n_460),
.Y(n_463)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_458),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_463),
.B(n_464),
.Y(n_467)
);


endmodule