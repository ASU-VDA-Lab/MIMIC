module fake_jpeg_3023_n_198 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_10),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_0),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_28),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_51),
.B1(n_65),
.B2(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_84),
.B1(n_75),
.B2(n_60),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_51),
.B1(n_65),
.B2(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_50),
.B1(n_57),
.B2(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_61),
.B1(n_67),
.B2(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_50),
.B1(n_67),
.B2(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_62),
.B1(n_54),
.B2(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_98),
.B(n_1),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_97),
.B1(n_104),
.B2(n_7),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_77),
.B(n_60),
.C(n_58),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_112),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_80),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_52),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_59),
.B1(n_58),
.B2(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_66),
.Y(n_105)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_53),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_69),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_29),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_34),
.B(n_47),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_12),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_130),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_4),
.B(n_6),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_15),
.B(n_21),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_98),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_31),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_9),
.C(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_131),
.Y(n_139)
);

AO21x2_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_30),
.B(n_48),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_126),
.B1(n_122),
.B2(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_7),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_12),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_150),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_146),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_156),
.B(n_24),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_142),
.B1(n_138),
.B2(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_32),
.C(n_43),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_153),
.C(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_14),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_14),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_129),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_35),
.C(n_16),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_36),
.C(n_18),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_49),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_162),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_164),
.B1(n_160),
.B2(n_167),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_42),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_168),
.C(n_134),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_135),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_137),
.B1(n_156),
.B2(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_176),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_154),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_166),
.B1(n_163),
.B2(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_165),
.C(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_25),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_162),
.Y(n_185)
);

AOI31xp67_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_178),
.A3(n_176),
.B(n_37),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_178),
.B1(n_174),
.B2(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_191),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_186),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_185),
.B(n_189),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_192),
.B(n_187),
.Y(n_195)
);

AOI21x1_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_182),
.B(n_41),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_40),
.Y(n_198)
);


endmodule