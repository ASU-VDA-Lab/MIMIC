module fake_netlist_1_12385_n_728 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_728);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_728;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g99 ( .A(n_93), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_36), .Y(n_100) );
BUFx5_ASAP7_75t_L g101 ( .A(n_31), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_13), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_95), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_22), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_45), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_59), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_60), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_30), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_82), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_65), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_69), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_78), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_23), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_47), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_29), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_54), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_49), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_55), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_26), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_7), .B(n_5), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_53), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_32), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_25), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_44), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_14), .Y(n_129) );
INVxp33_ASAP7_75t_SL g130 ( .A(n_12), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_12), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_11), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_43), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_71), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_61), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_38), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_99), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_116), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_101), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
NOR2x1_ASAP7_75t_L g144 ( .A(n_117), .B(n_0), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_100), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_103), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_101), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_118), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_103), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_104), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_134), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_129), .B(n_0), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_101), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_108), .B(n_1), .Y(n_155) );
BUFx12f_ASAP7_75t_L g156 ( .A(n_106), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_104), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_154), .B(n_105), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_138), .B(n_115), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_154), .B(n_121), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_156), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_142), .Y(n_163) );
BUFx10_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_153), .A2(n_130), .B1(n_102), .B2(n_129), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_138), .B(n_145), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_145), .B(n_137), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_146), .B(n_134), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_146), .B(n_123), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_147), .B(n_109), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_147), .B(n_132), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_151), .B(n_136), .C(n_135), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_155), .B(n_132), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_151), .B(n_123), .Y(n_184) );
CKINVDCx11_ASAP7_75t_R g185 ( .A(n_156), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_161), .B(n_153), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_167), .A2(n_153), .B1(n_155), .B2(n_157), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_181), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_179), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_161), .B(n_114), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_167), .A2(n_157), .B1(n_150), .B2(n_140), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_166), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_181), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_164), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_159), .B(n_140), .Y(n_196) );
INVx5_ASAP7_75t_L g197 ( .A(n_165), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_166), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_175), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_182), .B(n_140), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_182), .B(n_140), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_175), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_176), .B(n_140), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_178), .B(n_144), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_165), .B(n_119), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_169), .B(n_150), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_165), .B(n_133), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_178), .B(n_150), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_181), .B(n_150), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_181), .B(n_150), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_160), .B(n_157), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_177), .B(n_157), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_170), .B(n_157), .Y(n_217) );
OR2x2_ASAP7_75t_L g218 ( .A(n_162), .B(n_1), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
O2A1O1Ixp5_ASAP7_75t_L g220 ( .A1(n_158), .A2(n_112), .B(n_148), .C(n_107), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_180), .A2(n_144), .B1(n_148), .B2(n_149), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_177), .Y(n_222) );
NAND2xp33_ASAP7_75t_L g223 ( .A(n_163), .B(n_101), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_162), .A2(n_131), .B1(n_124), .B2(n_148), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_224), .A2(n_180), .B(n_184), .C(n_173), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_216), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_197), .B(n_164), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_187), .A2(n_163), .B(n_172), .Y(n_228) );
OAI22xp33_ASAP7_75t_SL g229 ( .A1(n_218), .A2(n_179), .B1(n_185), .B2(n_111), .Y(n_229) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_214), .A2(n_186), .B(n_168), .Y(n_230) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_193), .A2(n_172), .B(n_168), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_200), .A2(n_171), .B(n_125), .C(n_136), .Y(n_232) );
AO21x1_ASAP7_75t_L g233 ( .A1(n_223), .A2(n_120), .B(n_107), .Y(n_233) );
CKINVDCx8_ASAP7_75t_R g234 ( .A(n_204), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_190), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_192), .B(n_110), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_188), .A2(n_128), .B1(n_111), .B2(n_113), .Y(n_237) );
NOR3xp33_ASAP7_75t_SL g238 ( .A(n_191), .B(n_110), .C(n_113), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_188), .B(n_120), .Y(n_239) );
BUFx12f_ASAP7_75t_L g240 ( .A(n_218), .Y(n_240) );
NOR3xp33_ASAP7_75t_SL g241 ( .A(n_201), .B(n_122), .C(n_125), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_197), .B(n_122), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_192), .B(n_126), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_204), .B(n_126), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_204), .B(n_128), .Y(n_245) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_220), .A2(n_186), .B(n_127), .C(n_135), .Y(n_246) );
NAND2xp33_ASAP7_75t_L g247 ( .A(n_197), .B(n_101), .Y(n_247) );
INVxp67_ASAP7_75t_SL g248 ( .A(n_216), .Y(n_248) );
BUFx4f_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_211), .A2(n_212), .B(n_194), .C(n_189), .Y(n_250) );
OAI22x1_ASAP7_75t_L g251 ( .A1(n_213), .A2(n_127), .B1(n_3), .B2(n_4), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_197), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_208), .A2(n_149), .B1(n_152), .B2(n_143), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_210), .B(n_149), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_197), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_189), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_249), .B(n_216), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_234), .B(n_196), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_235), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_231), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_225), .A2(n_203), .B(n_217), .C(n_194), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_256), .Y(n_262) );
AO31x2_ASAP7_75t_L g263 ( .A1(n_250), .A2(n_198), .A3(n_215), .B(n_206), .Y(n_263) );
O2A1O1Ixp5_ASAP7_75t_SL g264 ( .A1(n_253), .A2(n_209), .B(n_205), .C(n_101), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_251), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_252), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_248), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_237), .A2(n_221), .B(n_219), .C(n_195), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_240), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_249), .B(n_219), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_232), .A2(n_195), .B(n_207), .C(n_213), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_244), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_229), .B(n_195), .Y(n_273) );
O2A1O1Ixp5_ASAP7_75t_L g274 ( .A1(n_233), .A2(n_202), .B(n_215), .C(n_198), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_248), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_255), .B(n_197), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_228), .A2(n_222), .B(n_195), .Y(n_277) );
CKINVDCx16_ASAP7_75t_R g278 ( .A(n_226), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_262), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_260), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_262), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_272), .B(n_239), .Y(n_282) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_260), .A2(n_246), .B(n_254), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_263), .Y(n_284) );
OR2x6_ASAP7_75t_L g285 ( .A(n_267), .B(n_226), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_264), .A2(n_230), .B(n_236), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_261), .A2(n_241), .B(n_243), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_277), .A2(n_247), .B(n_230), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_275), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_278), .B(n_244), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_275), .Y(n_292) );
BUFx12f_ASAP7_75t_L g293 ( .A(n_259), .Y(n_293) );
OAI221xp5_ASAP7_75t_L g294 ( .A1(n_265), .A2(n_245), .B1(n_241), .B2(n_238), .C(n_242), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_258), .A2(n_238), .B1(n_149), .B2(n_139), .C(n_143), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_274), .A2(n_198), .B(n_193), .Y(n_296) );
CKINVDCx6p67_ASAP7_75t_R g297 ( .A(n_257), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_257), .B(n_255), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_264), .B(n_149), .C(n_152), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_263), .Y(n_300) );
OA21x2_ASAP7_75t_L g301 ( .A1(n_299), .A2(n_271), .B(n_273), .Y(n_301) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_299), .A2(n_202), .B(n_206), .Y(n_302) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_288), .A2(n_202), .B(n_206), .Y(n_303) );
AOI21x1_ASAP7_75t_L g304 ( .A1(n_288), .A2(n_227), .B(n_215), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_285), .B(n_266), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_290), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_289), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
OAI21xp33_ASAP7_75t_L g309 ( .A1(n_282), .A2(n_270), .B(n_266), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_280), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_279), .B(n_263), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_300), .A2(n_268), .B(n_193), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_285), .B(n_276), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_295), .A2(n_276), .B(n_222), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_280), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_280), .A2(n_276), .B(n_252), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_285), .B(n_263), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_286), .A2(n_199), .B(n_207), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_286), .A2(n_199), .B(n_263), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_300), .A2(n_199), .B(n_139), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_279), .B(n_101), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_292), .Y(n_323) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_286), .A2(n_139), .B(n_141), .Y(n_324) );
OR2x6_ASAP7_75t_L g325 ( .A(n_285), .B(n_252), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_292), .B(n_252), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
AOI22xp33_ASAP7_75t_SL g328 ( .A1(n_287), .A2(n_259), .B1(n_269), .B2(n_101), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_281), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_285), .B(n_149), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_298), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_284), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_321), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_313), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_307), .B(n_308), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_306), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_310), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g340 ( .A(n_327), .B(n_284), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_316), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_318), .B(n_284), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_311), .B(n_298), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_313), .B(n_287), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_311), .B(n_287), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_318), .B(n_296), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_308), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_322), .B(n_287), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_323), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_322), .B(n_297), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_322), .B(n_297), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_313), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_313), .B(n_294), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_316), .B(n_291), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_313), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_329), .B(n_291), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
INVx4_ASAP7_75t_R g367 ( .A(n_330), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_309), .B(n_282), .Y(n_368) );
INVxp33_ASAP7_75t_L g369 ( .A(n_305), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_318), .Y(n_370) );
OAI321xp33_ASAP7_75t_L g371 ( .A1(n_309), .A2(n_294), .A3(n_295), .B1(n_296), .B2(n_149), .C(n_152), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_318), .B(n_283), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_331), .B(n_283), .Y(n_373) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_305), .B(n_283), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_313), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_331), .B(n_283), .Y(n_376) );
INVx5_ASAP7_75t_SL g377 ( .A(n_325), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_321), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_325), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
OR2x6_ASAP7_75t_L g381 ( .A(n_325), .B(n_305), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_325), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_321), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_324), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_357), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_321), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_347), .B(n_321), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_354), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_365), .B(n_305), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_365), .B(n_305), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_338), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_345), .B(n_328), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_354), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_357), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_338), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_345), .B(n_328), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_363), .B(n_326), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_367), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_338), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_332), .B(n_312), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_363), .B(n_326), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_332), .B(n_312), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_337), .B(n_312), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_336), .B(n_330), .Y(n_405) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_362), .B(n_325), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_358), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_351), .B(n_366), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_336), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_350), .B(n_330), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_351), .B(n_312), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_337), .B(n_312), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_341), .B(n_320), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_350), .B(n_325), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_341), .B(n_320), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_352), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_343), .B(n_320), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_339), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_366), .B(n_325), .Y(n_420) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_340), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_352), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_353), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_362), .B(n_333), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_353), .B(n_317), .Y(n_425) );
INVx5_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_339), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_339), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_370), .B(n_320), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_342), .Y(n_430) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_340), .Y(n_431) );
NAND2xp33_ASAP7_75t_R g432 ( .A(n_359), .B(n_269), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_342), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_342), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_370), .B(n_320), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_355), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_368), .B(n_317), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_373), .B(n_324), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_334), .B(n_324), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_373), .B(n_301), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_335), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_376), .B(n_301), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_343), .Y(n_443) );
OAI21x1_ASAP7_75t_SL g444 ( .A1(n_334), .A2(n_314), .B(n_301), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_348), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_355), .B(n_293), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_381), .B(n_303), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_368), .B(n_141), .C(n_143), .Y(n_448) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_334), .B(n_303), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_335), .B(n_301), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_376), .B(n_301), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g452 ( .A(n_333), .B(n_293), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_367), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_344), .B(n_301), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_348), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_348), .B(n_314), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_382), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_377), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_344), .B(n_303), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_360), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_344), .B(n_303), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_344), .B(n_303), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_359), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_360), .Y(n_464) );
NAND2x1_ASAP7_75t_L g465 ( .A(n_399), .B(n_381), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_389), .B(n_369), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_394), .B(n_381), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_443), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_408), .B(n_381), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_390), .B(n_381), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_441), .B(n_378), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_391), .B(n_375), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_412), .B(n_378), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_408), .B(n_375), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_387), .B(n_375), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_386), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_387), .B(n_360), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_464), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_464), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_412), .B(n_383), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_436), .B(n_356), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_395), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_445), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_457), .B(n_356), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_426), .B(n_356), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_401), .B(n_383), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_401), .B(n_333), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_392), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_407), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_409), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_463), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_388), .B(n_364), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_388), .B(n_364), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_446), .B(n_293), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_398), .B(n_361), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_420), .B(n_364), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_403), .B(n_333), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_403), .B(n_361), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_410), .B(n_361), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_426), .B(n_374), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_420), .B(n_346), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_417), .B(n_380), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_402), .B(n_379), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_426), .B(n_346), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_422), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_405), .B(n_377), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_392), .Y(n_507) );
NAND2xp33_ASAP7_75t_L g508 ( .A(n_399), .B(n_372), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_423), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_415), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_440), .B(n_380), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_411), .B(n_377), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_438), .B(n_377), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_393), .A2(n_346), .B1(n_349), .B2(n_377), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_438), .B(n_414), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_440), .B(n_380), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_442), .B(n_384), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_442), .B(n_384), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_451), .B(n_384), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_420), .B(n_346), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_396), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_425), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_414), .B(n_372), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_451), .B(n_346), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_416), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_416), .B(n_349), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_454), .B(n_374), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_450), .B(n_385), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_418), .B(n_349), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_454), .B(n_374), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_453), .B(n_349), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_429), .B(n_385), .Y(n_532) );
NOR2xp67_ASAP7_75t_L g533 ( .A(n_426), .B(n_371), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_453), .B(n_385), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_460), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_396), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_418), .Y(n_537) );
OAI211xp5_ASAP7_75t_L g538 ( .A1(n_452), .A2(n_152), .B(n_143), .C(n_141), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_429), .B(n_319), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_397), .B(n_2), .C(n_3), .D(n_4), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_459), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_426), .B(n_319), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_459), .B(n_319), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_400), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_461), .B(n_302), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_435), .B(n_302), .Y(n_546) );
NAND4xp75_ASAP7_75t_L g547 ( .A(n_406), .B(n_302), .C(n_371), .D(n_6), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_400), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_419), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_404), .B(n_2), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_458), .B(n_5), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_419), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_427), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_435), .B(n_302), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_461), .B(n_302), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_468), .Y(n_556) );
AND3x2_ASAP7_75t_L g557 ( .A(n_494), .B(n_421), .C(n_431), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_476), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_540), .A2(n_432), .B1(n_458), .B2(n_462), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_515), .B(n_404), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_491), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_491), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_482), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_489), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_551), .A2(n_447), .B1(n_424), .B2(n_437), .C(n_413), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_501), .B(n_439), .Y(n_567) );
OAI32xp33_ASAP7_75t_L g568 ( .A1(n_541), .A2(n_447), .A3(n_424), .B1(n_413), .B2(n_462), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_533), .A2(n_449), .B1(n_439), .B2(n_456), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_479), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_522), .B(n_427), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_490), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_510), .B(n_428), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_505), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_537), .Y(n_575) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_550), .A2(n_439), .B(n_449), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_525), .B(n_428), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_509), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_473), .B(n_430), .Y(n_579) );
AOI21xp33_ASAP7_75t_L g580 ( .A1(n_471), .A2(n_444), .B(n_448), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_471), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_473), .B(n_430), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_541), .Y(n_583) );
NOR2xp67_ASAP7_75t_L g584 ( .A(n_500), .B(n_433), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_503), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_480), .B(n_433), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_469), .B(n_434), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_495), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_535), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_523), .B(n_434), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_511), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_520), .B(n_455), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_524), .B(n_455), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_511), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_467), .B(n_302), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_474), .B(n_304), .Y(n_596) );
NOR3xp33_ASAP7_75t_L g597 ( .A(n_547), .B(n_304), .C(n_7), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_508), .A2(n_444), .B1(n_152), .B2(n_143), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_480), .B(n_141), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_465), .B(n_304), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_470), .B(n_6), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_479), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_486), .B(n_141), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_504), .B(n_8), .Y(n_604) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_514), .A2(n_141), .B(n_143), .C(n_152), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_492), .B(n_141), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_504), .B(n_141), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_538), .A2(n_8), .B(n_9), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_486), .B(n_143), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_516), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_466), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_493), .B(n_143), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_516), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_517), .B(n_518), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_517), .B(n_152), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_518), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_472), .B(n_9), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_519), .B(n_152), .Y(n_618) );
AOI31xp33_ASAP7_75t_L g619 ( .A1(n_485), .A2(n_10), .A3(n_11), .B(n_13), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_519), .B(n_487), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_499), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_485), .B(n_542), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_484), .Y(n_623) );
OR2x6_ASAP7_75t_L g624 ( .A(n_542), .B(n_10), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_487), .A2(n_174), .B(n_15), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_497), .B(n_14), .Y(n_626) );
AOI321xp33_ASAP7_75t_L g627 ( .A1(n_497), .A2(n_15), .A3(n_16), .B1(n_17), .B2(n_18), .C(n_19), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_532), .B(n_16), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_619), .A2(n_530), .B(n_527), .C(n_475), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_624), .A2(n_539), .B(n_528), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_560), .A2(n_478), .B(n_532), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_621), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_581), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_561), .B(n_498), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_589), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_624), .A2(n_528), .B(n_502), .C(n_529), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_560), .A2(n_526), .B(n_481), .C(n_496), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_611), .B(n_531), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_604), .A2(n_498), .B1(n_554), .B2(n_546), .C1(n_502), .C2(n_539), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_620), .B(n_477), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_556), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_591), .B(n_543), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_614), .B(n_546), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_558), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_567), .B(n_534), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_590), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_566), .B(n_544), .C(n_553), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_564), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_594), .B(n_549), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_565), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_610), .B(n_499), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_563), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_613), .B(n_616), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_572), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_601), .A2(n_555), .B1(n_545), .B2(n_554), .C1(n_548), .C2(n_552), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_570), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_588), .B(n_513), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_574), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_578), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_604), .A2(n_512), .B1(n_506), .B2(n_536), .Y(n_660) );
O2A1O1Ixp5_ASAP7_75t_L g661 ( .A1(n_568), .A2(n_521), .B(n_507), .C(n_488), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_608), .A2(n_17), .B(n_18), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_584), .B(n_569), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_617), .A2(n_174), .B1(n_19), .B2(n_20), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_585), .A2(n_174), .B1(n_20), .B2(n_207), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_606), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_625), .A2(n_207), .B(n_24), .Y(n_667) );
AOI32xp33_ASAP7_75t_L g668 ( .A1(n_597), .A2(n_21), .A3(n_27), .B1(n_28), .B2(n_33), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_562), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_612), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_599), .B(n_174), .C(n_35), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_584), .B(n_567), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g673 ( .A1(n_629), .A2(n_569), .B(n_625), .C(n_627), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_670), .A2(n_576), .B1(n_626), .B2(n_580), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_641), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_631), .A2(n_575), .B1(n_628), .B2(n_583), .C(n_586), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_663), .A2(n_607), .B(n_622), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_639), .A2(n_623), .B1(n_592), .B2(n_557), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_637), .A2(n_598), .B(n_603), .C(n_609), .Y(n_679) );
OAI221xp5_ASAP7_75t_SL g680 ( .A1(n_636), .A2(n_598), .B1(n_618), .B2(n_605), .C(n_602), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_632), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_672), .B(n_593), .Y(n_682) );
AOI332xp33_ASAP7_75t_L g683 ( .A1(n_633), .A2(n_559), .A3(n_582), .B1(n_579), .B2(n_573), .B3(n_571), .C1(n_577), .C2(n_592), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_639), .A2(n_615), .B(n_596), .C(n_595), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_647), .A2(n_587), .B1(n_600), .B2(n_174), .C(n_41), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_653), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g687 ( .A1(n_655), .A2(n_34), .B(n_37), .C(n_39), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_666), .A2(n_174), .B1(n_46), .B2(n_48), .Y(n_688) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_661), .A2(n_630), .B(n_672), .C(n_668), .Y(n_689) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_652), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_649), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_651), .Y(n_692) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_669), .A2(n_42), .B(n_50), .C(n_51), .Y(n_693) );
OAI21xp33_ASAP7_75t_SL g694 ( .A1(n_656), .A2(n_52), .B(n_56), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_656), .A2(n_662), .B(n_667), .C(n_666), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_683), .A2(n_660), .B(n_664), .C(n_638), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_673), .B(n_665), .C(n_671), .D(n_659), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_695), .B(n_658), .C(n_635), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_684), .A2(n_654), .B1(n_650), .B2(n_648), .C(n_644), .Y(n_699) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_690), .A2(n_642), .B1(n_646), .B2(n_645), .C1(n_657), .C2(n_643), .Y(n_700) );
NOR2xp33_ASAP7_75t_R g701 ( .A(n_675), .B(n_634), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_690), .A2(n_640), .B1(n_58), .B2(n_63), .C(n_64), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_689), .A2(n_57), .B(n_66), .Y(n_703) );
NOR4xp25_ASAP7_75t_L g704 ( .A(n_687), .B(n_67), .C(n_68), .D(n_70), .Y(n_704) );
NOR2xp67_ASAP7_75t_L g705 ( .A(n_694), .B(n_72), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_678), .A2(n_98), .B1(n_74), .B2(n_75), .C(n_76), .Y(n_706) );
AOI22xp5_ASAP7_75t_SL g707 ( .A1(n_677), .A2(n_73), .B1(n_77), .B2(n_79), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_699), .B(n_686), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_703), .B(n_693), .C(n_685), .Y(n_709) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_704), .B(n_674), .C(n_676), .Y(n_710) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_698), .B(n_674), .C(n_688), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_696), .A2(n_680), .B(n_679), .C(n_691), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_706), .B(n_692), .C(n_681), .Y(n_713) );
OA22x2_ASAP7_75t_L g714 ( .A1(n_708), .A2(n_701), .B1(n_682), .B2(n_700), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_712), .B(n_697), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_713), .Y(n_716) );
NOR5xp2_ASAP7_75t_L g717 ( .A(n_710), .B(n_707), .C(n_705), .D(n_702), .E(n_86), .Y(n_717) );
AND3x4_ASAP7_75t_L g718 ( .A(n_716), .B(n_709), .C(n_711), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_714), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_715), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_720), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_719), .Y(n_722) );
OA22x2_ASAP7_75t_L g723 ( .A1(n_722), .A2(n_718), .B1(n_717), .B2(n_85), .Y(n_723) );
NOR2xp67_ASAP7_75t_L g724 ( .A(n_721), .B(n_80), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_723), .A2(n_84), .B(n_87), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_724), .B(n_90), .Y(n_726) );
OA22x2_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_89), .B1(n_91), .B2(n_92), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_94), .B1(n_96), .B2(n_97), .Y(n_728) );
endmodule