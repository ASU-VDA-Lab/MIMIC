module fake_jpeg_20656_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_15),
.B1(n_14),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_14),
.B1(n_27),
.B2(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_15),
.B1(n_24),
.B2(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_38),
.B1(n_42),
.B2(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_22),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_16),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_70),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_32),
.C(n_38),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_85),
.C(n_58),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_75),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_28),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_84),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_59),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_88),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_26),
.C(n_30),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_64),
.B1(n_60),
.B2(n_44),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_1),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_46),
.B(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_60),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_82),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_7),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_10),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_88),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_76),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp67_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_74),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_60),
.B1(n_71),
.B2(n_65),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_77),
.B(n_84),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_119),
.Y(n_129)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_5),
.C(n_6),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_125),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_98),
.B1(n_105),
.B2(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_133),
.B1(n_117),
.B2(n_114),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_135),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_98),
.B1(n_105),
.B2(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_124),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_146),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_106),
.B1(n_123),
.B2(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_147),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_111),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_131),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_109),
.B(n_112),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_129),
.B(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_120),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_66),
.B(n_85),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_138),
.C(n_130),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_138),
.C(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_142),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_147),
.B(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_157),
.B(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_156),
.C(n_154),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_4),
.B1(n_102),
.B2(n_76),
.Y(n_167)
);

OAI321xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_161),
.A3(n_159),
.B1(n_153),
.B2(n_114),
.C(n_3),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_167),
.A2(n_4),
.B(n_69),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_168),
.B(n_59),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_170),
.B(n_59),
.Y(n_172)
);


endmodule